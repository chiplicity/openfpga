magic
tech EFS8A
magscale 1 2
timestamp 1602095330
<< locali >>
rect 8217 19873 8378 19907
rect 8217 19703 8251 19873
rect 14013 16031 14047 16201
rect 6279 13481 6285 13515
rect 11615 13481 11621 13515
rect 6279 13413 6313 13481
rect 11615 13413 11649 13481
rect 4537 12631 4571 12937
rect 7423 12257 7458 12291
rect 13380 11237 13448 11271
rect 8119 10455 8153 10523
rect 8119 10421 8125 10455
rect 5859 10081 5894 10115
rect 14473 9435 14507 9605
rect 11931 8993 11966 9027
rect 4905 7191 4939 7361
rect 6009 7259 6043 7429
rect 18791 6953 18797 6987
rect 18791 6885 18825 6953
rect 8027 5865 8033 5899
rect 8027 5797 8061 5865
rect 2415 5015 2449 5083
rect 2415 4981 2421 5015
rect 14013 4471 14047 4777
rect 15663 4777 15669 4811
rect 15663 4709 15697 4777
rect 8355 3689 8401 3723
rect 10051 3689 10057 3723
rect 10051 3621 10085 3689
rect 1547 2873 1685 2907
<< viali >>
rect 10952 20961 10986 20995
rect 11023 20757 11057 20791
rect 1593 20553 1627 20587
rect 3433 20553 3467 20587
rect 10701 20553 10735 20587
rect 11161 20553 11195 20587
rect 12633 20553 12667 20587
rect 17325 20553 17359 20587
rect 21097 20553 21131 20587
rect 22109 20553 22143 20587
rect 1409 20349 1443 20383
rect 3249 20349 3283 20383
rect 5432 20349 5466 20383
rect 5825 20349 5859 20383
rect 10517 20349 10551 20383
rect 12449 20349 12483 20383
rect 13001 20349 13035 20383
rect 16840 20349 16874 20383
rect 20612 20349 20646 20383
rect 21624 20349 21658 20383
rect 2053 20213 2087 20247
rect 3893 20213 3927 20247
rect 5503 20213 5537 20247
rect 10425 20213 10459 20247
rect 16911 20213 16945 20247
rect 20683 20213 20717 20247
rect 21695 20213 21729 20247
rect 8447 20009 8481 20043
rect 11483 20009 11517 20043
rect 1476 19873 1510 19907
rect 11412 19873 11446 19907
rect 1547 19669 1581 19703
rect 8217 19669 8251 19703
rect 1593 19465 1627 19499
rect 11713 19465 11747 19499
rect 14381 19465 14415 19499
rect 10609 19261 10643 19295
rect 10977 19261 11011 19295
rect 14197 19261 14231 19295
rect 8309 19125 8343 19159
rect 11161 19125 11195 19159
rect 14841 19125 14875 19159
rect 7113 18921 7147 18955
rect 11253 18853 11287 18887
rect 1444 18785 1478 18819
rect 6929 18785 6963 18819
rect 13645 18785 13679 18819
rect 20980 18785 21014 18819
rect 10057 18717 10091 18751
rect 11161 18717 11195 18751
rect 13369 18717 13403 18751
rect 11713 18649 11747 18683
rect 1547 18581 1581 18615
rect 8401 18581 8435 18615
rect 10885 18581 10919 18615
rect 21051 18581 21085 18615
rect 2237 18377 2271 18411
rect 6193 18377 6227 18411
rect 10609 18377 10643 18411
rect 11805 18377 11839 18411
rect 13369 18377 13403 18411
rect 15255 18377 15289 18411
rect 20913 18377 20947 18411
rect 6975 18309 7009 18343
rect 7665 18309 7699 18343
rect 8677 18241 8711 18275
rect 11529 18241 11563 18275
rect 14565 18241 14599 18275
rect 1444 18173 1478 18207
rect 1869 18173 1903 18207
rect 5800 18173 5834 18207
rect 6904 18173 6938 18207
rect 7297 18173 7331 18207
rect 15152 18173 15186 18207
rect 15577 18173 15611 18207
rect 8401 18105 8435 18139
rect 8493 18105 8527 18139
rect 10333 18105 10367 18139
rect 10885 18105 10919 18139
rect 10977 18105 11011 18139
rect 12541 18105 12575 18139
rect 13093 18105 13127 18139
rect 13645 18105 13679 18139
rect 13737 18105 13771 18139
rect 14289 18105 14323 18139
rect 1547 18037 1581 18071
rect 5871 18037 5905 18071
rect 8217 18037 8251 18071
rect 5733 17765 5767 17799
rect 8033 17765 8067 17799
rect 10241 17765 10275 17799
rect 10793 17765 10827 17799
rect 13645 17765 13679 17799
rect 14197 17765 14231 17799
rect 1444 17697 1478 17731
rect 2789 17697 2823 17731
rect 11713 17697 11747 17731
rect 15368 17697 15402 17731
rect 20980 17697 21014 17731
rect 5641 17629 5675 17663
rect 5917 17629 5951 17663
rect 7941 17629 7975 17663
rect 8585 17629 8619 17663
rect 10149 17629 10183 17663
rect 11621 17629 11655 17663
rect 13553 17629 13587 17663
rect 13277 17561 13311 17595
rect 1547 17493 1581 17527
rect 2697 17493 2731 17527
rect 5273 17493 5307 17527
rect 15439 17493 15473 17527
rect 21051 17493 21085 17527
rect 1869 17289 1903 17323
rect 8217 17289 8251 17323
rect 10057 17289 10091 17323
rect 11713 17289 11747 17323
rect 15393 17289 15427 17323
rect 21005 17289 21039 17323
rect 8953 17221 8987 17255
rect 2697 17153 2731 17187
rect 3157 17153 3191 17187
rect 4629 17153 4663 17187
rect 5273 17153 5307 17187
rect 5917 17153 5951 17187
rect 9597 17153 9631 17187
rect 10885 17153 10919 17187
rect 13277 17153 13311 17187
rect 13553 17153 13587 17187
rect 1476 17085 1510 17119
rect 2237 17085 2271 17119
rect 7481 17085 7515 17119
rect 7849 17085 7883 17119
rect 8401 17085 8435 17119
rect 2789 17017 2823 17051
rect 3617 17017 3651 17051
rect 3985 17017 4019 17051
rect 5365 17017 5399 17051
rect 6837 17017 6871 17051
rect 10609 17017 10643 17051
rect 10701 17017 10735 17051
rect 13369 17017 13403 17051
rect 1547 16949 1581 16983
rect 5089 16949 5123 16983
rect 6193 16949 6227 16983
rect 10425 16949 10459 16983
rect 13001 16949 13035 16983
rect 14197 16949 14231 16983
rect 3433 16745 3467 16779
rect 8401 16745 8435 16779
rect 13645 16745 13679 16779
rect 2605 16677 2639 16711
rect 3157 16677 3191 16711
rect 6009 16677 6043 16711
rect 7843 16677 7877 16711
rect 12817 16677 12851 16711
rect 13369 16677 13403 16711
rect 1476 16609 1510 16643
rect 5365 16609 5399 16643
rect 9965 16609 9999 16643
rect 10149 16609 10183 16643
rect 20980 16609 21014 16643
rect 2513 16541 2547 16575
rect 7481 16541 7515 16575
rect 10241 16541 10275 16575
rect 12725 16541 12759 16575
rect 1547 16405 1581 16439
rect 7113 16405 7147 16439
rect 10701 16405 10735 16439
rect 21051 16405 21085 16439
rect 1593 16201 1627 16235
rect 2421 16201 2455 16235
rect 3801 16201 3835 16235
rect 5641 16201 5675 16235
rect 5917 16201 5951 16235
rect 10517 16201 10551 16235
rect 11897 16201 11931 16235
rect 14013 16201 14047 16235
rect 21005 16201 21039 16235
rect 13461 16133 13495 16167
rect 7389 16065 7423 16099
rect 14289 16065 14323 16099
rect 1409 15997 1443 16031
rect 2881 15997 2915 16031
rect 4721 15997 4755 16031
rect 9597 15997 9631 16031
rect 10793 15997 10827 16031
rect 12541 15997 12575 16031
rect 13737 15997 13771 16031
rect 14013 15997 14047 16031
rect 14197 15997 14231 16031
rect 14381 15997 14415 16031
rect 2789 15929 2823 15963
rect 3202 15929 3236 15963
rect 4537 15929 4571 15963
rect 5042 15929 5076 15963
rect 7113 15929 7147 15963
rect 7205 15929 7239 15963
rect 9413 15929 9447 15963
rect 9918 15929 9952 15963
rect 12862 15929 12896 15963
rect 1961 15861 1995 15895
rect 4077 15861 4111 15895
rect 6561 15861 6595 15895
rect 8033 15861 8067 15895
rect 8401 15861 8435 15895
rect 9137 15861 9171 15895
rect 12265 15861 12299 15895
rect 1547 15657 1581 15691
rect 1869 15657 1903 15691
rect 2697 15657 2731 15691
rect 3433 15657 3467 15691
rect 8585 15657 8619 15691
rect 9965 15657 9999 15691
rect 10977 15657 11011 15691
rect 13093 15657 13127 15691
rect 6193 15589 6227 15623
rect 7205 15589 7239 15623
rect 10419 15589 10453 15623
rect 12494 15589 12528 15623
rect 1476 15521 1510 15555
rect 2697 15521 2731 15555
rect 2973 15521 3007 15555
rect 6101 15521 6135 15555
rect 10057 15521 10091 15555
rect 7113 15453 7147 15487
rect 7389 15453 7423 15487
rect 12173 15453 12207 15487
rect 4721 15317 4755 15351
rect 6837 15317 6871 15351
rect 13369 15317 13403 15351
rect 3157 15113 3191 15147
rect 3617 15113 3651 15147
rect 5549 15113 5583 15147
rect 6285 15113 6319 15147
rect 7757 15113 7791 15147
rect 15623 15113 15657 15147
rect 10609 15045 10643 15079
rect 14565 15045 14599 15079
rect 4721 14977 4755 15011
rect 9781 14977 9815 15011
rect 10333 14977 10367 15011
rect 12265 14977 12299 15011
rect 13185 14977 13219 15011
rect 1685 14909 1719 14943
rect 1869 14909 1903 14943
rect 4077 14909 4111 14943
rect 4445 14909 4479 14943
rect 4629 14909 4663 14943
rect 6837 14909 6871 14943
rect 9229 14909 9263 14943
rect 9689 14909 9723 14943
rect 11529 14909 11563 14943
rect 12449 14909 12483 14943
rect 12909 14909 12943 14943
rect 14381 14909 14415 14943
rect 14933 14909 14967 14943
rect 15552 14909 15586 14943
rect 15945 14909 15979 14943
rect 7158 14841 7192 14875
rect 11897 14841 11931 14875
rect 2053 14773 2087 14807
rect 2789 14773 2823 14807
rect 6561 14773 6595 14807
rect 9137 14773 9171 14807
rect 1593 14569 1627 14603
rect 9321 14569 9355 14603
rect 12449 14569 12483 14603
rect 13323 14569 13357 14603
rect 1869 14501 1903 14535
rect 1961 14501 1995 14535
rect 5641 14501 5675 14535
rect 6561 14501 6595 14535
rect 6653 14501 6687 14535
rect 12173 14501 12207 14535
rect 15485 14501 15519 14535
rect 5181 14433 5215 14467
rect 5457 14433 5491 14467
rect 10057 14433 10091 14467
rect 11437 14433 11471 14467
rect 11989 14433 12023 14467
rect 13252 14433 13286 14467
rect 2513 14365 2547 14399
rect 14197 14365 14231 14399
rect 15393 14365 15427 14399
rect 15669 14365 15703 14399
rect 7113 14297 7147 14331
rect 3801 14229 3835 14263
rect 7573 14229 7607 14263
rect 9965 14229 9999 14263
rect 14933 14229 14967 14263
rect 1777 14025 1811 14059
rect 2881 14025 2915 14059
rect 5089 14025 5123 14059
rect 5825 14025 5859 14059
rect 10057 14025 10091 14059
rect 11805 14025 11839 14059
rect 14749 14025 14783 14059
rect 15853 14025 15887 14059
rect 4721 13957 4755 13991
rect 1961 13889 1995 13923
rect 3249 13889 3283 13923
rect 3801 13889 3835 13923
rect 9137 13889 9171 13923
rect 14933 13889 14967 13923
rect 15577 13889 15611 13923
rect 16497 13889 16531 13923
rect 16773 13889 16807 13923
rect 6193 13821 6227 13855
rect 6561 13821 6595 13855
rect 6929 13821 6963 13855
rect 2053 13753 2087 13787
rect 2605 13753 2639 13787
rect 4123 13753 4157 13787
rect 7573 13753 7607 13787
rect 8953 13753 8987 13787
rect 9229 13753 9263 13787
rect 9781 13753 9815 13787
rect 12541 13753 12575 13787
rect 12633 13753 12667 13787
rect 13185 13753 13219 13787
rect 15025 13753 15059 13787
rect 16313 13753 16347 13787
rect 16589 13753 16623 13787
rect 3709 13685 3743 13719
rect 5457 13685 5491 13719
rect 11345 13685 11379 13719
rect 12173 13685 12207 13719
rect 13461 13685 13495 13719
rect 2605 13481 2639 13515
rect 4169 13481 4203 13515
rect 6285 13481 6319 13515
rect 6837 13481 6871 13515
rect 9045 13481 9079 13515
rect 11621 13481 11655 13515
rect 12817 13481 12851 13515
rect 15577 13481 15611 13515
rect 16497 13481 16531 13515
rect 7849 13413 7883 13447
rect 9873 13413 9907 13447
rect 13185 13413 13219 13447
rect 17049 13413 17083 13447
rect 1777 13345 1811 13379
rect 4077 13345 4111 13379
rect 4537 13345 4571 13379
rect 14933 13345 14967 13379
rect 15485 13345 15519 13379
rect 20980 13345 21014 13379
rect 5917 13277 5951 13311
rect 7757 13277 7791 13311
rect 8033 13277 8067 13311
rect 9781 13277 9815 13311
rect 10057 13277 10091 13311
rect 11253 13277 11287 13311
rect 13093 13277 13127 13311
rect 13461 13277 13495 13311
rect 16957 13277 16991 13311
rect 17325 13277 17359 13311
rect 1869 13141 1903 13175
rect 2973 13141 3007 13175
rect 3709 13141 3743 13175
rect 5273 13141 5307 13175
rect 7113 13141 7147 13175
rect 10793 13141 10827 13175
rect 12173 13141 12207 13175
rect 12449 13141 12483 13175
rect 14289 13141 14323 13175
rect 21051 13141 21085 13175
rect 3433 12937 3467 12971
rect 4537 12937 4571 12971
rect 7665 12937 7699 12971
rect 9965 12937 9999 12971
rect 10241 12937 10275 12971
rect 15209 12937 15243 12971
rect 15485 12937 15519 12971
rect 16681 12937 16715 12971
rect 21465 12937 21499 12971
rect 3065 12869 3099 12903
rect 1685 12801 1719 12835
rect 3617 12733 3651 12767
rect 4169 12733 4203 12767
rect 1777 12665 1811 12699
rect 2329 12665 2363 12699
rect 6193 12869 6227 12903
rect 6653 12869 6687 12903
rect 5917 12801 5951 12835
rect 7297 12801 7331 12835
rect 9045 12801 9079 12835
rect 11345 12801 11379 12835
rect 13185 12801 13219 12835
rect 13461 12801 13495 12835
rect 14289 12801 14323 12835
rect 20453 12801 20487 12835
rect 5457 12733 5491 12767
rect 5733 12733 5767 12767
rect 6872 12733 6906 12767
rect 10793 12733 10827 12767
rect 11253 12733 11287 12767
rect 12265 12733 12299 12767
rect 12541 12733 12575 12767
rect 16313 12733 16347 12767
rect 17049 12733 17083 12767
rect 17417 12733 17451 12767
rect 8861 12665 8895 12699
rect 9366 12665 9400 12699
rect 11805 12665 11839 12699
rect 14197 12665 14231 12699
rect 14651 12665 14685 12699
rect 20545 12665 20579 12699
rect 21097 12665 21131 12699
rect 2605 12597 2639 12631
rect 3893 12597 3927 12631
rect 4537 12597 4571 12631
rect 4721 12597 4755 12631
rect 5089 12597 5123 12631
rect 6975 12597 7009 12631
rect 8125 12597 8159 12631
rect 10609 12597 10643 12631
rect 20177 12597 20211 12631
rect 4997 12393 5031 12427
rect 6469 12393 6503 12427
rect 9137 12393 9171 12427
rect 9781 12393 9815 12427
rect 11161 12393 11195 12427
rect 13001 12393 13035 12427
rect 16589 12393 16623 12427
rect 20453 12393 20487 12427
rect 1777 12325 1811 12359
rect 3893 12325 3927 12359
rect 4439 12325 4473 12359
rect 11253 12325 11287 12359
rect 14381 12325 14415 12359
rect 16031 12325 16065 12359
rect 19993 12325 20027 12359
rect 21005 12325 21039 12359
rect 21097 12325 21131 12359
rect 4077 12257 4111 12291
rect 5825 12257 5859 12291
rect 7389 12257 7423 12291
rect 9689 12257 9723 12291
rect 10149 12257 10183 12291
rect 11400 12257 11434 12291
rect 13645 12257 13679 12291
rect 14197 12257 14231 12291
rect 19901 12257 19935 12291
rect 1685 12189 1719 12223
rect 2053 12189 2087 12223
rect 6193 12189 6227 12223
rect 11621 12189 11655 12223
rect 15669 12189 15703 12223
rect 21281 12189 21315 12223
rect 5990 12121 6024 12155
rect 6929 12121 6963 12155
rect 11529 12121 11563 12155
rect 2789 12053 2823 12087
rect 5365 12053 5399 12087
rect 5733 12053 5767 12087
rect 6101 12053 6135 12087
rect 7297 12053 7331 12087
rect 7527 12053 7561 12087
rect 9413 12053 9447 12087
rect 10701 12053 10735 12087
rect 11897 12053 11931 12087
rect 16957 12053 16991 12087
rect 18337 12053 18371 12087
rect 5641 11849 5675 11883
rect 8125 11849 8159 11883
rect 9045 11849 9079 11883
rect 10517 11849 10551 11883
rect 13001 11849 13035 11883
rect 19257 11849 19291 11883
rect 19625 11849 19659 11883
rect 20821 11849 20855 11883
rect 21741 11849 21775 11883
rect 5089 11781 5123 11815
rect 5457 11781 5491 11815
rect 10333 11781 10367 11815
rect 14657 11781 14691 11815
rect 21051 11781 21085 11815
rect 21465 11781 21499 11815
rect 1869 11713 1903 11747
rect 5549 11713 5583 11747
rect 10425 11713 10459 11747
rect 15853 11713 15887 11747
rect 16497 11713 16531 11747
rect 1476 11645 1510 11679
rect 2697 11645 2731 11679
rect 5328 11645 5362 11679
rect 7113 11645 7147 11679
rect 7481 11645 7515 11679
rect 7849 11645 7883 11679
rect 10204 11645 10238 11679
rect 11621 11645 11655 11679
rect 14013 11645 14047 11679
rect 15393 11645 15427 11679
rect 15577 11645 15611 11679
rect 18337 11645 18371 11679
rect 20980 11645 21014 11679
rect 2605 11577 2639 11611
rect 3059 11577 3093 11611
rect 5181 11577 5215 11611
rect 9321 11577 9355 11611
rect 10057 11577 10091 11611
rect 16221 11577 16255 11611
rect 18658 11577 18692 11611
rect 1547 11509 1581 11543
rect 3617 11509 3651 11543
rect 4169 11509 4203 11543
rect 4721 11509 4755 11543
rect 6285 11509 6319 11543
rect 6653 11509 6687 11543
rect 9689 11509 9723 11543
rect 11253 11509 11287 11543
rect 11989 11509 12023 11543
rect 12725 11509 12759 11543
rect 13369 11509 13403 11543
rect 13829 11509 13863 11543
rect 15025 11509 15059 11543
rect 2789 11305 2823 11339
rect 4169 11305 4203 11339
rect 5181 11305 5215 11339
rect 6561 11305 6595 11339
rect 7389 11305 7423 11339
rect 10241 11305 10275 11339
rect 13001 11305 13035 11339
rect 15393 11305 15427 11339
rect 18429 11305 18463 11339
rect 1961 11237 1995 11271
rect 3893 11237 3927 11271
rect 5917 11237 5951 11271
rect 8769 11237 8803 11271
rect 11713 11237 11747 11271
rect 13346 11237 13380 11271
rect 17877 11237 17911 11271
rect 4353 11169 4387 11203
rect 4537 11169 4571 11203
rect 6064 11169 6098 11203
rect 8033 11169 8067 11203
rect 9724 11169 9758 11203
rect 10977 11169 11011 11203
rect 12449 11169 12483 11203
rect 13093 11169 13127 11203
rect 14013 11169 14047 11203
rect 14289 11169 14323 11203
rect 15393 11169 15427 11203
rect 15853 11169 15887 11203
rect 17417 11169 17451 11203
rect 17601 11169 17635 11203
rect 1869 11101 1903 11135
rect 6285 11101 6319 11135
rect 8401 11101 8435 11135
rect 11345 11101 11379 11135
rect 1685 11033 1719 11067
rect 2421 11033 2455 11067
rect 9827 11033 9861 11067
rect 5733 10965 5767 10999
rect 6193 10965 6227 10999
rect 7113 10965 7147 10999
rect 7849 10965 7883 10999
rect 8198 10965 8232 10999
rect 8309 10965 8343 10999
rect 9413 10965 9447 10999
rect 10517 10965 10551 10999
rect 11115 10965 11149 10999
rect 11253 10965 11287 10999
rect 11989 10965 12023 10999
rect 3433 10761 3467 10795
rect 4997 10761 5031 10795
rect 5346 10761 5380 10795
rect 6561 10761 6595 10795
rect 7205 10761 7239 10795
rect 13461 10761 13495 10795
rect 13921 10761 13955 10795
rect 15301 10761 15335 10795
rect 2605 10693 2639 10727
rect 5457 10693 5491 10727
rect 7573 10693 7607 10727
rect 10977 10693 11011 10727
rect 12725 10693 12759 10727
rect 13093 10693 13127 10727
rect 16037 10693 16071 10727
rect 17509 10693 17543 10727
rect 1869 10625 1903 10659
rect 3525 10625 3559 10659
rect 4537 10625 4571 10659
rect 5549 10625 5583 10659
rect 5641 10625 5675 10659
rect 9873 10625 9907 10659
rect 12817 10625 12851 10659
rect 14381 10625 14415 10659
rect 3065 10557 3099 10591
rect 3617 10557 3651 10591
rect 7757 10557 7791 10591
rect 8677 10557 8711 10591
rect 9321 10557 9355 10591
rect 11412 10557 11446 10591
rect 12596 10557 12630 10591
rect 19901 10557 19935 10591
rect 20637 10557 20671 10591
rect 21624 10557 21658 10591
rect 2053 10489 2087 10523
rect 2145 10489 2179 10523
rect 5181 10489 5215 10523
rect 8953 10489 8987 10523
rect 9597 10489 9631 10523
rect 9689 10489 9723 10523
rect 11805 10489 11839 10523
rect 12449 10489 12483 10523
rect 14105 10489 14139 10523
rect 14197 10489 14231 10523
rect 6285 10421 6319 10455
rect 8125 10421 8159 10455
rect 10701 10421 10735 10455
rect 11483 10421 11517 10455
rect 12173 10421 12207 10455
rect 15577 10421 15611 10455
rect 17233 10421 17267 10455
rect 20269 10421 20303 10455
rect 21695 10421 21729 10455
rect 22109 10421 22143 10455
rect 3157 10217 3191 10251
rect 3617 10217 3651 10251
rect 4353 10217 4387 10251
rect 5365 10217 5399 10251
rect 5641 10217 5675 10251
rect 7941 10217 7975 10251
rect 8769 10217 8803 10251
rect 12817 10217 12851 10251
rect 14749 10217 14783 10251
rect 9413 10149 9447 10183
rect 13829 10149 13863 10183
rect 14381 10149 14415 10183
rect 21097 10149 21131 10183
rect 2237 10081 2271 10115
rect 4353 10081 4387 10115
rect 4721 10081 4755 10115
rect 5825 10081 5859 10115
rect 6745 10081 6779 10115
rect 7205 10081 7239 10115
rect 7481 10081 7515 10115
rect 7849 10081 7883 10115
rect 9781 10081 9815 10115
rect 11345 10081 11379 10115
rect 15945 10081 15979 10115
rect 17417 10081 17451 10115
rect 17601 10081 17635 10115
rect 2145 10013 2179 10047
rect 8401 10013 8435 10047
rect 9689 10013 9723 10047
rect 11253 10013 11287 10047
rect 13737 10013 13771 10047
rect 15393 10013 15427 10047
rect 17877 10013 17911 10047
rect 21005 10013 21039 10047
rect 1869 9945 1903 9979
rect 10793 9945 10827 9979
rect 13185 9945 13219 9979
rect 21557 9945 21591 9979
rect 5963 9877 5997 9911
rect 6377 9877 6411 9911
rect 12449 9877 12483 9911
rect 2145 9673 2179 9707
rect 3801 9673 3835 9707
rect 4169 9673 4203 9707
rect 5825 9673 5859 9707
rect 6653 9673 6687 9707
rect 9597 9673 9631 9707
rect 10609 9673 10643 9707
rect 11069 9673 11103 9707
rect 11437 9673 11471 9707
rect 11805 9673 11839 9707
rect 12173 9673 12207 9707
rect 14197 9673 14231 9707
rect 19165 9673 19199 9707
rect 20269 9673 20303 9707
rect 21465 9673 21499 9707
rect 21833 9673 21867 9707
rect 2973 9605 3007 9639
rect 7389 9605 7423 9639
rect 14473 9605 14507 9639
rect 14565 9605 14599 9639
rect 2421 9537 2455 9571
rect 6837 9537 6871 9571
rect 9137 9537 9171 9571
rect 10333 9537 10367 9571
rect 10940 9537 10974 9571
rect 11161 9537 11195 9571
rect 4629 9469 4663 9503
rect 13185 9469 13219 9503
rect 13645 9469 13679 9503
rect 13921 9469 13955 9503
rect 18245 9537 18279 9571
rect 20545 9537 20579 9571
rect 21189 9537 21223 9571
rect 14749 9469 14783 9503
rect 2513 9401 2547 9435
rect 4950 9401 4984 9435
rect 8493 9401 8527 9435
rect 8585 9401 8619 9435
rect 9965 9401 9999 9435
rect 10793 9401 10827 9435
rect 14473 9401 14507 9435
rect 15070 9401 15104 9435
rect 17785 9401 17819 9435
rect 18566 9401 18600 9435
rect 20637 9401 20671 9435
rect 1869 9333 1903 9367
rect 3433 9333 3467 9367
rect 4445 9333 4479 9367
rect 5549 9333 5583 9367
rect 7757 9333 7791 9367
rect 8309 9333 8343 9367
rect 13001 9333 13035 9367
rect 15669 9333 15703 9367
rect 15945 9333 15979 9367
rect 16497 9333 16531 9367
rect 17233 9333 17267 9367
rect 4261 9129 4295 9163
rect 4629 9129 4663 9163
rect 5273 9129 5307 9163
rect 8217 9129 8251 9163
rect 8677 9129 8711 9163
rect 12035 9129 12069 9163
rect 14289 9129 14323 9163
rect 14749 9129 14783 9163
rect 15669 9129 15703 9163
rect 17233 9129 17267 9163
rect 18245 9129 18279 9163
rect 20545 9129 20579 9163
rect 2053 9061 2087 9095
rect 5733 9061 5767 9095
rect 13369 9061 13403 9095
rect 15945 9061 15979 9095
rect 4065 8993 4099 9027
rect 10977 8993 11011 9027
rect 11897 8993 11931 9027
rect 20980 8993 21014 9027
rect 1961 8925 1995 8959
rect 5641 8925 5675 8959
rect 7113 8925 7147 8959
rect 10333 8925 10367 8959
rect 13277 8925 13311 8959
rect 15853 8925 15887 8959
rect 16221 8925 16255 8959
rect 2513 8857 2547 8891
rect 6193 8857 6227 8891
rect 13829 8857 13863 8891
rect 21051 8857 21085 8891
rect 1685 8789 1719 8823
rect 7849 8789 7883 8823
rect 2421 8585 2455 8619
rect 4169 8585 4203 8619
rect 5089 8585 5123 8619
rect 10609 8585 10643 8619
rect 14565 8585 14599 8619
rect 15393 8585 15427 8619
rect 16589 8585 16623 8619
rect 21465 8585 21499 8619
rect 21833 8585 21867 8619
rect 2053 8517 2087 8551
rect 4629 8517 4663 8551
rect 10149 8517 10183 8551
rect 11989 8517 12023 8551
rect 16221 8517 16255 8551
rect 3249 8449 3283 8483
rect 5273 8449 5307 8483
rect 9045 8449 9079 8483
rect 9597 8449 9631 8483
rect 11069 8449 11103 8483
rect 12541 8449 12575 8483
rect 13645 8449 13679 8483
rect 13921 8449 13955 8483
rect 15669 8449 15703 8483
rect 1409 8381 1443 8415
rect 7757 8381 7791 8415
rect 20980 8381 21014 8415
rect 3570 8313 3604 8347
rect 5365 8313 5399 8347
rect 5917 8313 5951 8347
rect 7573 8313 7607 8347
rect 8078 8313 8112 8347
rect 9689 8313 9723 8347
rect 13737 8313 13771 8347
rect 15761 8313 15795 8347
rect 1593 8245 1627 8279
rect 3065 8245 3099 8279
rect 6193 8245 6227 8279
rect 8677 8245 8711 8279
rect 9413 8245 9447 8279
rect 13277 8245 13311 8279
rect 15025 8245 15059 8279
rect 21051 8245 21085 8279
rect 3893 8041 3927 8075
rect 7849 8041 7883 8075
rect 15853 8041 15887 8075
rect 21051 8041 21085 8075
rect 2329 7973 2363 8007
rect 5917 7973 5951 8007
rect 9689 7973 9723 8007
rect 12862 7973 12896 8007
rect 4123 7905 4157 7939
rect 5089 7905 5123 7939
rect 5365 7905 5399 7939
rect 7205 7905 7239 7939
rect 7389 7905 7423 7939
rect 7757 7905 7791 7939
rect 9781 7905 9815 7939
rect 15368 7905 15402 7939
rect 20980 7905 21014 7939
rect 2237 7837 2271 7871
rect 2513 7837 2547 7871
rect 4537 7837 4571 7871
rect 12541 7837 12575 7871
rect 14381 7769 14415 7803
rect 1685 7701 1719 7735
rect 1961 7701 1995 7735
rect 3341 7701 3375 7735
rect 4215 7701 4249 7735
rect 8861 7701 8895 7735
rect 10793 7701 10827 7735
rect 13461 7701 13495 7735
rect 14105 7701 14139 7735
rect 15439 7701 15473 7735
rect 2697 7497 2731 7531
rect 4077 7497 4111 7531
rect 5346 7497 5380 7531
rect 8033 7497 8067 7531
rect 8677 7497 8711 7531
rect 9781 7497 9815 7531
rect 15393 7497 15427 7531
rect 21189 7497 21223 7531
rect 5457 7429 5491 7463
rect 6009 7429 6043 7463
rect 9413 7429 9447 7463
rect 11069 7429 11103 7463
rect 2329 7361 2363 7395
rect 4905 7361 4939 7395
rect 5549 7361 5583 7395
rect 3157 7293 3191 7327
rect 1685 7225 1719 7259
rect 1777 7225 1811 7259
rect 3478 7225 3512 7259
rect 4629 7225 4663 7259
rect 7389 7361 7423 7395
rect 10940 7361 10974 7395
rect 11161 7361 11195 7395
rect 11529 7361 11563 7395
rect 11897 7361 11931 7395
rect 6837 7293 6871 7327
rect 12449 7293 12483 7327
rect 13001 7293 13035 7327
rect 14013 7293 14047 7327
rect 14473 7293 14507 7327
rect 18061 7293 18095 7327
rect 18521 7293 18555 7327
rect 19993 7293 20027 7327
rect 20729 7293 20763 7327
rect 5181 7225 5215 7259
rect 6009 7225 6043 7259
rect 6285 7225 6319 7259
rect 8861 7225 8895 7259
rect 8953 7225 8987 7259
rect 10333 7225 10367 7259
rect 10793 7225 10827 7259
rect 14749 7225 14783 7259
rect 3065 7157 3099 7191
rect 4905 7157 4939 7191
rect 4997 7157 5031 7191
rect 5825 7157 5859 7191
rect 6653 7157 6687 7191
rect 7757 7157 7791 7191
rect 10609 7157 10643 7191
rect 12265 7157 12299 7191
rect 12725 7157 12759 7191
rect 13921 7157 13955 7191
rect 17785 7157 17819 7191
rect 18337 7157 18371 7191
rect 20361 7157 20395 7191
rect 2789 6953 2823 6987
rect 3249 6953 3283 6987
rect 4169 6953 4203 6987
rect 5273 6953 5307 6987
rect 7297 6953 7331 6987
rect 7849 6953 7883 6987
rect 10885 6953 10919 6987
rect 12817 6953 12851 6987
rect 13369 6953 13403 6987
rect 18061 6953 18095 6987
rect 18797 6953 18831 6987
rect 19349 6953 19383 6987
rect 5641 6885 5675 6919
rect 7021 6885 7055 6919
rect 8217 6885 8251 6919
rect 11989 6885 12023 6919
rect 16405 6885 16439 6919
rect 21097 6885 21131 6919
rect 1685 6817 1719 6851
rect 1777 6817 1811 6851
rect 2421 6817 2455 6851
rect 4353 6817 4387 6851
rect 4629 6817 4663 6851
rect 5788 6817 5822 6851
rect 9965 6817 9999 6851
rect 11253 6817 11287 6851
rect 13645 6817 13679 6851
rect 18429 6817 18463 6851
rect 3801 6749 3835 6783
rect 6009 6749 6043 6783
rect 8125 6749 8159 6783
rect 8769 6749 8803 6783
rect 9689 6749 9723 6783
rect 11400 6749 11434 6783
rect 11621 6749 11655 6783
rect 16313 6749 16347 6783
rect 21005 6749 21039 6783
rect 6101 6681 6135 6715
rect 11529 6681 11563 6715
rect 16865 6681 16899 6715
rect 21557 6681 21591 6715
rect 5917 6613 5951 6647
rect 9045 6613 9079 6647
rect 12449 6613 12483 6647
rect 2421 6409 2455 6443
rect 4813 6409 4847 6443
rect 6193 6409 6227 6443
rect 8401 6409 8435 6443
rect 9965 6409 9999 6443
rect 10425 6409 10459 6443
rect 11529 6409 11563 6443
rect 11897 6409 11931 6443
rect 12725 6409 12759 6443
rect 14841 6409 14875 6443
rect 15853 6409 15887 6443
rect 16313 6409 16347 6443
rect 18797 6409 18831 6443
rect 20361 6409 20395 6443
rect 21557 6409 21591 6443
rect 3249 6341 3283 6375
rect 21189 6341 21223 6375
rect 2053 6273 2087 6307
rect 9321 6273 9355 6307
rect 14933 6273 14967 6307
rect 16589 6273 16623 6307
rect 18521 6273 18555 6307
rect 20085 6273 20119 6307
rect 1409 6205 1443 6239
rect 2513 6205 2547 6239
rect 3617 6205 3651 6239
rect 3985 6205 4019 6239
rect 4261 6205 4295 6239
rect 5181 6205 5215 6239
rect 5549 6205 5583 6239
rect 7205 6205 7239 6239
rect 7389 6205 7423 6239
rect 7757 6205 7791 6239
rect 10977 6205 11011 6239
rect 13645 6205 13679 6239
rect 14013 6205 14047 6239
rect 16840 6205 16874 6239
rect 5365 6137 5399 6171
rect 5917 6137 5951 6171
rect 9045 6137 9079 6171
rect 9137 6137 9171 6171
rect 10517 6137 10551 6171
rect 15254 6137 15288 6171
rect 20637 6137 20671 6171
rect 20729 6137 20763 6171
rect 1593 6069 1627 6103
rect 2697 6069 2731 6103
rect 3801 6069 3835 6103
rect 6653 6069 6687 6103
rect 7849 6069 7883 6103
rect 8861 6069 8895 6103
rect 13277 6069 13311 6103
rect 16911 6069 16945 6103
rect 17325 6069 17359 6103
rect 2881 5865 2915 5899
rect 4169 5865 4203 5899
rect 8033 5865 8067 5899
rect 8585 5865 8619 5899
rect 9045 5865 9079 5899
rect 11897 5865 11931 5899
rect 13369 5865 13403 5899
rect 13645 5865 13679 5899
rect 14933 5865 14967 5899
rect 18429 5865 18463 5899
rect 20177 5865 20211 5899
rect 20637 5865 20671 5899
rect 21051 5865 21085 5899
rect 3525 5797 3559 5831
rect 12770 5797 12804 5831
rect 16589 5797 16623 5831
rect 1685 5729 1719 5763
rect 1869 5729 1903 5763
rect 4353 5729 4387 5763
rect 4629 5729 4663 5763
rect 6009 5729 6043 5763
rect 6285 5729 6319 5763
rect 6837 5729 6871 5763
rect 7665 5729 7699 5763
rect 10885 5729 10919 5763
rect 11437 5729 11471 5763
rect 20980 5729 21014 5763
rect 1777 5661 1811 5695
rect 3893 5661 3927 5695
rect 5457 5661 5491 5695
rect 11621 5661 11655 5695
rect 12449 5661 12483 5695
rect 16497 5661 16531 5695
rect 16865 5661 16899 5695
rect 5825 5525 5859 5559
rect 7297 5525 7331 5559
rect 2973 5321 3007 5355
rect 3801 5321 3835 5355
rect 6561 5321 6595 5355
rect 7113 5321 7147 5355
rect 7297 5321 7331 5355
rect 7941 5321 7975 5355
rect 9183 5321 9217 5355
rect 10958 5321 10992 5355
rect 12173 5321 12207 5355
rect 13277 5321 13311 5355
rect 15853 5321 15887 5355
rect 21189 5321 21223 5355
rect 5273 5253 5307 5287
rect 8861 5253 8895 5287
rect 9321 5253 9355 5287
rect 10609 5253 10643 5287
rect 11069 5253 11103 5287
rect 14473 5253 14507 5287
rect 2053 5185 2087 5219
rect 3433 5185 3467 5219
rect 7205 5185 7239 5219
rect 9413 5185 9447 5219
rect 11161 5185 11195 5219
rect 13461 5185 13495 5219
rect 13829 5185 13863 5219
rect 16681 5185 16715 5219
rect 16957 5185 16991 5219
rect 20177 5185 20211 5219
rect 20453 5185 20487 5219
rect 3893 5117 3927 5151
rect 4445 5117 4479 5151
rect 5492 5117 5526 5151
rect 6984 5117 7018 5151
rect 8585 5117 8619 5151
rect 9045 5117 9079 5151
rect 10793 5117 10827 5151
rect 11805 5117 11839 5151
rect 16037 5117 16071 5151
rect 17877 5117 17911 5151
rect 18337 5117 18371 5151
rect 5917 5049 5951 5083
rect 6837 5049 6871 5083
rect 11529 5049 11563 5083
rect 13553 5049 13587 5083
rect 18699 5049 18733 5083
rect 20269 5049 20303 5083
rect 1961 4981 1995 5015
rect 2421 4981 2455 5015
rect 3985 4981 4019 5015
rect 4997 4981 5031 5015
rect 5595 4981 5629 5015
rect 9689 4981 9723 5015
rect 10241 4981 10275 5015
rect 12633 4981 12667 5015
rect 19257 4981 19291 5015
rect 19901 4981 19935 5015
rect 3893 4777 3927 4811
rect 6101 4777 6135 4811
rect 7205 4777 7239 4811
rect 7757 4777 7791 4811
rect 9045 4777 9079 4811
rect 10885 4777 10919 4811
rect 14013 4777 14047 4811
rect 2421 4709 2455 4743
rect 4398 4709 4432 4743
rect 6837 4709 6871 4743
rect 11713 4709 11747 4743
rect 12449 4709 12483 4743
rect 13277 4709 13311 4743
rect 13829 4709 13863 4743
rect 5917 4641 5951 4675
rect 9689 4641 9723 4675
rect 10149 4641 10183 4675
rect 2329 4573 2363 4607
rect 2605 4573 2639 4607
rect 4077 4573 4111 4607
rect 8677 4573 8711 4607
rect 10241 4573 10275 4607
rect 11253 4573 11287 4607
rect 13185 4573 13219 4607
rect 15669 4777 15703 4811
rect 16589 4777 16623 4811
rect 18153 4709 18187 4743
rect 21097 4709 21131 4743
rect 17509 4641 17543 4675
rect 17877 4641 17911 4675
rect 19860 4641 19894 4675
rect 15301 4573 15335 4607
rect 19947 4573 19981 4607
rect 21005 4573 21039 4607
rect 21557 4505 21591 4539
rect 1869 4437 1903 4471
rect 4997 4437 5031 4471
rect 14013 4437 14047 4471
rect 14197 4437 14231 4471
rect 16221 4437 16255 4471
rect 1685 4233 1719 4267
rect 4997 4233 5031 4267
rect 9689 4233 9723 4267
rect 11345 4233 11379 4267
rect 12817 4233 12851 4267
rect 17049 4233 17083 4267
rect 19717 4233 19751 4267
rect 21281 4233 21315 4267
rect 2881 4165 2915 4199
rect 4537 4165 4571 4199
rect 8401 4165 8435 4199
rect 13369 4165 13403 4199
rect 17785 4165 17819 4199
rect 2513 4097 2547 4131
rect 3433 4097 3467 4131
rect 3985 4097 4019 4131
rect 12909 4097 12943 4131
rect 14749 4097 14783 4131
rect 16497 4097 16531 4131
rect 6872 4029 6906 4063
rect 7297 4029 7331 4063
rect 8585 4029 8619 4063
rect 9137 4029 9171 4063
rect 10149 4029 10183 4063
rect 13921 4029 13955 4063
rect 14013 4029 14047 4063
rect 14473 4029 14507 4063
rect 19901 4029 19935 4063
rect 1869 3961 1903 3995
rect 1961 3961 1995 3995
rect 3801 3961 3835 3995
rect 4086 3961 4120 3995
rect 9321 3961 9355 3995
rect 10057 3961 10091 3995
rect 10511 3961 10545 3995
rect 15301 3961 15335 3995
rect 16129 3961 16163 3995
rect 16221 3961 16255 3995
rect 20545 3961 20579 3995
rect 20913 3961 20947 3995
rect 5825 3893 5859 3927
rect 6975 3893 7009 3927
rect 11069 3893 11103 3927
rect 15945 3893 15979 3927
rect 17509 3893 17543 3927
rect 1593 3689 1627 3723
rect 2329 3689 2363 3723
rect 4261 3689 4295 3723
rect 8401 3689 8435 3723
rect 9413 3689 9447 3723
rect 10057 3689 10091 3723
rect 10885 3689 10919 3723
rect 12449 3689 12483 3723
rect 15669 3689 15703 3723
rect 19901 3689 19935 3723
rect 2513 3621 2547 3655
rect 4629 3621 4663 3655
rect 11621 3621 11655 3655
rect 15945 3621 15979 3655
rect 16865 3621 16899 3655
rect 1409 3553 1443 3587
rect 7056 3553 7090 3587
rect 8284 3553 8318 3587
rect 9689 3553 9723 3587
rect 13001 3553 13035 3587
rect 14140 3553 14174 3587
rect 16497 3553 16531 3587
rect 4537 3485 4571 3519
rect 4813 3485 4847 3519
rect 11529 3485 11563 3519
rect 12173 3485 12207 3519
rect 15853 3485 15887 3519
rect 17325 3485 17359 3519
rect 6837 3349 6871 3383
rect 7159 3349 7193 3383
rect 10609 3349 10643 3383
rect 13185 3349 13219 3383
rect 14243 3349 14277 3383
rect 2559 3145 2593 3179
rect 4077 3145 4111 3179
rect 10057 3145 10091 3179
rect 10425 3145 10459 3179
rect 13461 3145 13495 3179
rect 14105 3145 14139 3179
rect 15485 3145 15519 3179
rect 15117 3077 15151 3111
rect 2329 3009 2363 3043
rect 4997 3009 5031 3043
rect 5273 3009 5307 3043
rect 7389 3009 7423 3043
rect 10609 3009 10643 3043
rect 10977 3009 11011 3043
rect 12541 3009 12575 3043
rect 12817 3009 12851 3043
rect 16313 3009 16347 3043
rect 16589 3009 16623 3043
rect 1476 2941 1510 2975
rect 1869 2941 1903 2975
rect 2488 2941 2522 2975
rect 2881 2941 2915 2975
rect 4353 2941 4387 2975
rect 7021 2941 7055 2975
rect 8861 2941 8895 2975
rect 9597 2941 9631 2975
rect 14616 2941 14650 2975
rect 16221 2941 16255 2975
rect 18404 2941 18438 2975
rect 1685 2873 1719 2907
rect 6837 2873 6871 2907
rect 10701 2873 10735 2907
rect 12633 2873 12667 2907
rect 14703 2873 14737 2907
rect 6653 2805 6687 2839
rect 7757 2805 7791 2839
rect 8309 2805 8343 2839
rect 9413 2805 9447 2839
rect 11621 2805 11655 2839
rect 12265 2805 12299 2839
rect 18475 2805 18509 2839
rect 18889 2805 18923 2839
rect 1547 2601 1581 2635
rect 9505 2601 9539 2635
rect 10793 2601 10827 2635
rect 21327 2601 21361 2635
rect 6009 2533 6043 2567
rect 9873 2533 9907 2567
rect 9965 2533 9999 2567
rect 10517 2533 10551 2567
rect 11989 2533 12023 2567
rect 12633 2533 12667 2567
rect 1476 2465 1510 2499
rect 1869 2465 1903 2499
rect 4537 2465 4571 2499
rect 5181 2465 5215 2499
rect 5917 2465 5951 2499
rect 6377 2465 6411 2499
rect 6929 2465 6963 2499
rect 7297 2465 7331 2499
rect 7665 2465 7699 2499
rect 8493 2465 8527 2499
rect 9045 2465 9079 2499
rect 11437 2465 11471 2499
rect 12449 2465 12483 2499
rect 12725 2465 12759 2499
rect 14248 2465 14282 2499
rect 14657 2465 14691 2499
rect 15485 2465 15519 2499
rect 16037 2465 16071 2499
rect 16589 2465 16623 2499
rect 17141 2465 17175 2499
rect 20060 2465 20094 2499
rect 21256 2465 21290 2499
rect 6745 2397 6779 2431
rect 11161 2397 11195 2431
rect 13645 2397 13679 2431
rect 14335 2397 14369 2431
rect 8677 2329 8711 2363
rect 11621 2329 11655 2363
rect 15669 2261 15703 2295
rect 16773 2261 16807 2295
rect 20131 2261 20165 2295
rect 20545 2261 20579 2295
rect 21741 2261 21775 2295
<< metal1 >>
rect 1104 21786 22816 21808
rect 1104 21734 4982 21786
rect 5034 21734 5046 21786
rect 5098 21734 5110 21786
rect 5162 21734 5174 21786
rect 5226 21734 12982 21786
rect 13034 21734 13046 21786
rect 13098 21734 13110 21786
rect 13162 21734 13174 21786
rect 13226 21734 20982 21786
rect 21034 21734 21046 21786
rect 21098 21734 21110 21786
rect 21162 21734 21174 21786
rect 21226 21734 22816 21786
rect 1104 21712 22816 21734
rect 11146 21360 11152 21412
rect 11204 21400 11210 21412
rect 23566 21400 23572 21412
rect 11204 21372 23572 21400
rect 11204 21360 11210 21372
rect 23566 21360 23572 21372
rect 23624 21360 23630 21412
rect 1104 21242 22816 21264
rect 1104 21190 8982 21242
rect 9034 21190 9046 21242
rect 9098 21190 9110 21242
rect 9162 21190 9174 21242
rect 9226 21190 16982 21242
rect 17034 21190 17046 21242
rect 17098 21190 17110 21242
rect 17162 21190 17174 21242
rect 17226 21190 22816 21242
rect 1104 21168 22816 21190
rect 10940 20995 10998 21001
rect 10940 20961 10952 20995
rect 10986 20992 10998 20995
rect 11146 20992 11152 21004
rect 10986 20964 11152 20992
rect 10986 20961 10998 20964
rect 10940 20955 10998 20961
rect 11146 20952 11152 20964
rect 11204 20952 11210 21004
rect 9950 20748 9956 20800
rect 10008 20788 10014 20800
rect 11011 20791 11069 20797
rect 11011 20788 11023 20791
rect 10008 20760 11023 20788
rect 10008 20748 10014 20760
rect 11011 20757 11023 20760
rect 11057 20757 11069 20791
rect 11011 20751 11069 20757
rect 1104 20698 22816 20720
rect 1104 20646 4982 20698
rect 5034 20646 5046 20698
rect 5098 20646 5110 20698
rect 5162 20646 5174 20698
rect 5226 20646 12982 20698
rect 13034 20646 13046 20698
rect 13098 20646 13110 20698
rect 13162 20646 13174 20698
rect 13226 20646 20982 20698
rect 21034 20646 21046 20698
rect 21098 20646 21110 20698
rect 21162 20646 21174 20698
rect 21226 20646 22816 20698
rect 1104 20624 22816 20646
rect 1578 20584 1584 20596
rect 1539 20556 1584 20584
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 3418 20584 3424 20596
rect 3379 20556 3424 20584
rect 3418 20544 3424 20556
rect 3476 20544 3482 20596
rect 10686 20584 10692 20596
rect 10647 20556 10692 20584
rect 10686 20544 10692 20556
rect 10744 20544 10750 20596
rect 11146 20584 11152 20596
rect 11107 20556 11152 20584
rect 11146 20544 11152 20556
rect 11204 20544 11210 20596
rect 12621 20587 12679 20593
rect 12621 20553 12633 20587
rect 12667 20584 12679 20587
rect 12802 20584 12808 20596
rect 12667 20556 12808 20584
rect 12667 20553 12679 20556
rect 12621 20547 12679 20553
rect 12802 20544 12808 20556
rect 12860 20544 12866 20596
rect 17313 20587 17371 20593
rect 17313 20553 17325 20587
rect 17359 20584 17371 20587
rect 17678 20584 17684 20596
rect 17359 20556 17684 20584
rect 17359 20553 17371 20556
rect 17313 20547 17371 20553
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 3237 20383 3295 20389
rect 1443 20352 2084 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 2056 20256 2084 20352
rect 3237 20349 3249 20383
rect 3283 20380 3295 20383
rect 5420 20383 5478 20389
rect 3283 20352 3924 20380
rect 3283 20349 3295 20352
rect 3237 20343 3295 20349
rect 3896 20256 3924 20352
rect 5420 20349 5432 20383
rect 5466 20380 5478 20383
rect 5810 20380 5816 20392
rect 5466 20352 5816 20380
rect 5466 20349 5478 20352
rect 5420 20343 5478 20349
rect 5810 20340 5816 20352
rect 5868 20340 5874 20392
rect 10505 20383 10563 20389
rect 10505 20349 10517 20383
rect 10551 20349 10563 20383
rect 12434 20380 12440 20392
rect 12347 20352 12440 20380
rect 10505 20343 10563 20349
rect 2038 20244 2044 20256
rect 1999 20216 2044 20244
rect 2038 20204 2044 20216
rect 2096 20204 2102 20256
rect 3878 20244 3884 20256
rect 3839 20216 3884 20244
rect 3878 20204 3884 20216
rect 3936 20204 3942 20256
rect 5491 20247 5549 20253
rect 5491 20213 5503 20247
rect 5537 20244 5549 20247
rect 5810 20244 5816 20256
rect 5537 20216 5816 20244
rect 5537 20213 5549 20216
rect 5491 20207 5549 20213
rect 5810 20204 5816 20216
rect 5868 20204 5874 20256
rect 10413 20247 10471 20253
rect 10413 20213 10425 20247
rect 10459 20244 10471 20247
rect 10520 20244 10548 20343
rect 12434 20340 12440 20352
rect 12492 20380 12498 20392
rect 12989 20383 13047 20389
rect 12989 20380 13001 20383
rect 12492 20352 13001 20380
rect 12492 20340 12498 20352
rect 12989 20349 13001 20352
rect 13035 20349 13047 20383
rect 12989 20343 13047 20349
rect 16828 20383 16886 20389
rect 16828 20349 16840 20383
rect 16874 20380 16886 20383
rect 17328 20380 17356 20547
rect 17678 20544 17684 20556
rect 17736 20544 17742 20596
rect 21085 20587 21143 20593
rect 21085 20553 21097 20587
rect 21131 20584 21143 20587
rect 21634 20584 21640 20596
rect 21131 20556 21640 20584
rect 21131 20553 21143 20556
rect 21085 20547 21143 20553
rect 16874 20352 17356 20380
rect 20600 20383 20658 20389
rect 16874 20349 16886 20352
rect 16828 20343 16886 20349
rect 20600 20349 20612 20383
rect 20646 20380 20658 20383
rect 21100 20380 21128 20547
rect 21634 20544 21640 20556
rect 21692 20544 21698 20596
rect 22097 20587 22155 20593
rect 22097 20553 22109 20587
rect 22143 20584 22155 20587
rect 22462 20584 22468 20596
rect 22143 20556 22468 20584
rect 22143 20553 22155 20556
rect 22097 20547 22155 20553
rect 20646 20352 21128 20380
rect 21612 20383 21670 20389
rect 20646 20349 20658 20352
rect 20600 20343 20658 20349
rect 21612 20349 21624 20383
rect 21658 20380 21670 20383
rect 22112 20380 22140 20547
rect 22462 20544 22468 20556
rect 22520 20544 22526 20596
rect 21658 20352 22140 20380
rect 21658 20349 21670 20352
rect 21612 20343 21670 20349
rect 10686 20244 10692 20256
rect 10459 20216 10692 20244
rect 10459 20213 10471 20216
rect 10413 20207 10471 20213
rect 10686 20204 10692 20216
rect 10744 20204 10750 20256
rect 16482 20204 16488 20256
rect 16540 20244 16546 20256
rect 16899 20247 16957 20253
rect 16899 20244 16911 20247
rect 16540 20216 16911 20244
rect 16540 20204 16546 20216
rect 16899 20213 16911 20216
rect 16945 20213 16957 20247
rect 16899 20207 16957 20213
rect 20530 20204 20536 20256
rect 20588 20244 20594 20256
rect 20671 20247 20729 20253
rect 20671 20244 20683 20247
rect 20588 20216 20683 20244
rect 20588 20204 20594 20216
rect 20671 20213 20683 20216
rect 20717 20213 20729 20247
rect 20671 20207 20729 20213
rect 21683 20247 21741 20253
rect 21683 20213 21695 20247
rect 21729 20244 21741 20247
rect 21818 20244 21824 20256
rect 21729 20216 21824 20244
rect 21729 20213 21741 20216
rect 21683 20207 21741 20213
rect 21818 20204 21824 20216
rect 21876 20204 21882 20256
rect 1104 20154 22816 20176
rect 1104 20102 8982 20154
rect 9034 20102 9046 20154
rect 9098 20102 9110 20154
rect 9162 20102 9174 20154
rect 9226 20102 16982 20154
rect 17034 20102 17046 20154
rect 17098 20102 17110 20154
rect 17162 20102 17174 20154
rect 17226 20102 22816 20154
rect 1104 20080 22816 20102
rect 3878 20000 3884 20052
rect 3936 20040 3942 20052
rect 8435 20043 8493 20049
rect 8435 20040 8447 20043
rect 3936 20012 8447 20040
rect 3936 20000 3942 20012
rect 8435 20009 8447 20012
rect 8481 20009 8493 20043
rect 8435 20003 8493 20009
rect 11471 20043 11529 20049
rect 11471 20009 11483 20043
rect 11517 20040 11529 20043
rect 12434 20040 12440 20052
rect 11517 20012 12440 20040
rect 11517 20009 11529 20012
rect 11471 20003 11529 20009
rect 12434 20000 12440 20012
rect 12492 20000 12498 20052
rect 1210 19932 1216 19984
rect 1268 19972 1274 19984
rect 1268 19944 1507 19972
rect 1268 19932 1274 19944
rect 1479 19913 1507 19944
rect 1464 19907 1522 19913
rect 1464 19873 1476 19907
rect 1510 19873 1522 19907
rect 1464 19867 1522 19873
rect 11400 19907 11458 19913
rect 11400 19873 11412 19907
rect 11446 19904 11458 19907
rect 11698 19904 11704 19916
rect 11446 19876 11704 19904
rect 11446 19873 11458 19876
rect 11400 19867 11458 19873
rect 11698 19864 11704 19876
rect 11756 19864 11762 19916
rect 1535 19703 1593 19709
rect 1535 19669 1547 19703
rect 1581 19700 1593 19703
rect 2866 19700 2872 19712
rect 1581 19672 2872 19700
rect 1581 19669 1593 19672
rect 1535 19663 1593 19669
rect 2866 19660 2872 19672
rect 2924 19660 2930 19712
rect 8205 19703 8263 19709
rect 8205 19669 8217 19703
rect 8251 19700 8263 19703
rect 8294 19700 8300 19712
rect 8251 19672 8300 19700
rect 8251 19669 8263 19672
rect 8205 19663 8263 19669
rect 8294 19660 8300 19672
rect 8352 19660 8358 19712
rect 1104 19610 22816 19632
rect 1104 19558 4982 19610
rect 5034 19558 5046 19610
rect 5098 19558 5110 19610
rect 5162 19558 5174 19610
rect 5226 19558 12982 19610
rect 13034 19558 13046 19610
rect 13098 19558 13110 19610
rect 13162 19558 13174 19610
rect 13226 19558 20982 19610
rect 21034 19558 21046 19610
rect 21098 19558 21110 19610
rect 21162 19558 21174 19610
rect 21226 19558 22816 19610
rect 1104 19536 22816 19558
rect 1210 19456 1216 19508
rect 1268 19496 1274 19508
rect 1581 19499 1639 19505
rect 1581 19496 1593 19499
rect 1268 19468 1593 19496
rect 1268 19456 1274 19468
rect 1581 19465 1593 19468
rect 1627 19465 1639 19499
rect 11698 19496 11704 19508
rect 11659 19468 11704 19496
rect 1581 19459 1639 19465
rect 11698 19456 11704 19468
rect 11756 19456 11762 19508
rect 14369 19499 14427 19505
rect 14369 19465 14381 19499
rect 14415 19496 14427 19499
rect 15654 19496 15660 19508
rect 14415 19468 15660 19496
rect 14415 19465 14427 19468
rect 14369 19459 14427 19465
rect 15654 19456 15660 19468
rect 15712 19456 15718 19508
rect 10597 19295 10655 19301
rect 10597 19261 10609 19295
rect 10643 19292 10655 19295
rect 10962 19292 10968 19304
rect 10643 19264 10968 19292
rect 10643 19261 10655 19264
rect 10597 19255 10655 19261
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 14185 19295 14243 19301
rect 14185 19261 14197 19295
rect 14231 19292 14243 19295
rect 14231 19264 14872 19292
rect 14231 19261 14243 19264
rect 14185 19255 14243 19261
rect 14844 19168 14872 19264
rect 8294 19156 8300 19168
rect 8255 19128 8300 19156
rect 8294 19116 8300 19128
rect 8352 19116 8358 19168
rect 11146 19156 11152 19168
rect 11107 19128 11152 19156
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 14826 19156 14832 19168
rect 14787 19128 14832 19156
rect 14826 19116 14832 19128
rect 14884 19116 14890 19168
rect 1104 19066 22816 19088
rect 1104 19014 8982 19066
rect 9034 19014 9046 19066
rect 9098 19014 9110 19066
rect 9162 19014 9174 19066
rect 9226 19014 16982 19066
rect 17034 19014 17046 19066
rect 17098 19014 17110 19066
rect 17162 19014 17174 19066
rect 17226 19014 22816 19066
rect 1104 18992 22816 19014
rect 7101 18955 7159 18961
rect 7101 18921 7113 18955
rect 7147 18952 7159 18955
rect 8478 18952 8484 18964
rect 7147 18924 8484 18952
rect 7147 18921 7159 18924
rect 7101 18915 7159 18921
rect 8478 18912 8484 18924
rect 8536 18912 8542 18964
rect 11146 18844 11152 18896
rect 11204 18884 11210 18896
rect 11241 18887 11299 18893
rect 11241 18884 11253 18887
rect 11204 18856 11253 18884
rect 11204 18844 11210 18856
rect 11241 18853 11253 18856
rect 11287 18853 11299 18887
rect 11241 18847 11299 18853
rect 1302 18776 1308 18828
rect 1360 18816 1366 18828
rect 1432 18819 1490 18825
rect 1432 18816 1444 18819
rect 1360 18788 1444 18816
rect 1360 18776 1366 18788
rect 1432 18785 1444 18788
rect 1478 18785 1490 18819
rect 6914 18816 6920 18828
rect 6875 18788 6920 18816
rect 1432 18779 1490 18785
rect 6914 18776 6920 18788
rect 6972 18776 6978 18828
rect 13630 18816 13636 18828
rect 13591 18788 13636 18816
rect 13630 18776 13636 18788
rect 13688 18776 13694 18828
rect 20806 18776 20812 18828
rect 20864 18816 20870 18828
rect 20968 18819 21026 18825
rect 20968 18816 20980 18819
rect 20864 18788 20980 18816
rect 20864 18776 20870 18788
rect 20968 18785 20980 18788
rect 21014 18816 21026 18819
rect 21266 18816 21272 18828
rect 21014 18788 21272 18816
rect 21014 18785 21026 18788
rect 20968 18779 21026 18785
rect 21266 18776 21272 18788
rect 21324 18776 21330 18828
rect 10045 18751 10103 18757
rect 10045 18717 10057 18751
rect 10091 18748 10103 18751
rect 10594 18748 10600 18760
rect 10091 18720 10600 18748
rect 10091 18717 10103 18720
rect 10045 18711 10103 18717
rect 10594 18708 10600 18720
rect 10652 18748 10658 18760
rect 11149 18751 11207 18757
rect 11149 18748 11161 18751
rect 10652 18720 11161 18748
rect 10652 18708 10658 18720
rect 11149 18717 11161 18720
rect 11195 18717 11207 18751
rect 13354 18748 13360 18760
rect 13315 18720 13360 18748
rect 11149 18711 11207 18717
rect 13354 18708 13360 18720
rect 13412 18708 13418 18760
rect 11698 18680 11704 18692
rect 11659 18652 11704 18680
rect 11698 18640 11704 18652
rect 11756 18640 11762 18692
rect 1535 18615 1593 18621
rect 1535 18581 1547 18615
rect 1581 18612 1593 18615
rect 8110 18612 8116 18624
rect 1581 18584 8116 18612
rect 1581 18581 1593 18584
rect 1535 18575 1593 18581
rect 8110 18572 8116 18584
rect 8168 18572 8174 18624
rect 8386 18612 8392 18624
rect 8347 18584 8392 18612
rect 8386 18572 8392 18584
rect 8444 18572 8450 18624
rect 10873 18615 10931 18621
rect 10873 18581 10885 18615
rect 10919 18612 10931 18615
rect 10962 18612 10968 18624
rect 10919 18584 10968 18612
rect 10919 18581 10931 18584
rect 10873 18575 10931 18581
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 16022 18572 16028 18624
rect 16080 18612 16086 18624
rect 21039 18615 21097 18621
rect 21039 18612 21051 18615
rect 16080 18584 21051 18612
rect 16080 18572 16086 18584
rect 21039 18581 21051 18584
rect 21085 18581 21097 18615
rect 21039 18575 21097 18581
rect 1104 18522 22816 18544
rect 1104 18470 4982 18522
rect 5034 18470 5046 18522
rect 5098 18470 5110 18522
rect 5162 18470 5174 18522
rect 5226 18470 12982 18522
rect 13034 18470 13046 18522
rect 13098 18470 13110 18522
rect 13162 18470 13174 18522
rect 13226 18470 20982 18522
rect 21034 18470 21046 18522
rect 21098 18470 21110 18522
rect 21162 18470 21174 18522
rect 21226 18470 22816 18522
rect 1104 18448 22816 18470
rect 1302 18368 1308 18420
rect 1360 18408 1366 18420
rect 2225 18411 2283 18417
rect 2225 18408 2237 18411
rect 1360 18380 2237 18408
rect 1360 18368 1366 18380
rect 2225 18377 2237 18380
rect 2271 18377 2283 18411
rect 6178 18408 6184 18420
rect 6139 18380 6184 18408
rect 2225 18371 2283 18377
rect 6178 18368 6184 18380
rect 6236 18368 6242 18420
rect 10594 18408 10600 18420
rect 10555 18380 10600 18408
rect 10594 18368 10600 18380
rect 10652 18368 10658 18420
rect 11146 18368 11152 18420
rect 11204 18408 11210 18420
rect 11793 18411 11851 18417
rect 11793 18408 11805 18411
rect 11204 18380 11805 18408
rect 11204 18368 11210 18380
rect 11793 18377 11805 18380
rect 11839 18377 11851 18411
rect 13354 18408 13360 18420
rect 13315 18380 13360 18408
rect 11793 18371 11851 18377
rect 13354 18368 13360 18380
rect 13412 18368 13418 18420
rect 14826 18368 14832 18420
rect 14884 18408 14890 18420
rect 15243 18411 15301 18417
rect 15243 18408 15255 18411
rect 14884 18380 15255 18408
rect 14884 18368 14890 18380
rect 15243 18377 15255 18380
rect 15289 18377 15301 18411
rect 15243 18371 15301 18377
rect 20806 18368 20812 18420
rect 20864 18408 20870 18420
rect 20901 18411 20959 18417
rect 20901 18408 20913 18411
rect 20864 18380 20913 18408
rect 20864 18368 20870 18380
rect 20901 18377 20913 18380
rect 20947 18377 20959 18411
rect 20901 18371 20959 18377
rect 6914 18340 6920 18352
rect 6873 18312 6920 18340
rect 6914 18300 6920 18312
rect 6972 18349 6978 18352
rect 6972 18343 7021 18349
rect 6972 18309 6975 18343
rect 7009 18340 7021 18343
rect 7653 18343 7711 18349
rect 7653 18340 7665 18343
rect 7009 18312 7665 18340
rect 7009 18309 7021 18312
rect 6972 18303 7021 18309
rect 7653 18309 7665 18312
rect 7699 18309 7711 18343
rect 7653 18303 7711 18309
rect 6972 18300 6978 18303
rect 5902 18232 5908 18284
rect 5960 18272 5966 18284
rect 8662 18272 8668 18284
rect 5960 18244 6935 18272
rect 8623 18244 8668 18272
rect 5960 18232 5966 18244
rect 1210 18164 1216 18216
rect 1268 18204 1274 18216
rect 1432 18207 1490 18213
rect 1432 18204 1444 18207
rect 1268 18176 1444 18204
rect 1268 18164 1274 18176
rect 1432 18173 1444 18176
rect 1478 18204 1490 18207
rect 1857 18207 1915 18213
rect 1857 18204 1869 18207
rect 1478 18176 1869 18204
rect 1478 18173 1490 18176
rect 1432 18167 1490 18173
rect 1857 18173 1869 18176
rect 1903 18173 1915 18207
rect 1857 18167 1915 18173
rect 5788 18207 5846 18213
rect 5788 18173 5800 18207
rect 5834 18204 5846 18207
rect 6178 18204 6184 18216
rect 5834 18176 6184 18204
rect 5834 18173 5846 18176
rect 5788 18167 5846 18173
rect 6178 18164 6184 18176
rect 6236 18164 6242 18216
rect 6907 18213 6935 18244
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18272 11575 18275
rect 11698 18272 11704 18284
rect 11563 18244 11704 18272
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 11698 18232 11704 18244
rect 11756 18232 11762 18284
rect 13630 18232 13636 18284
rect 13688 18272 13694 18284
rect 14553 18275 14611 18281
rect 14553 18272 14565 18275
rect 13688 18244 14565 18272
rect 13688 18232 13694 18244
rect 14553 18241 14565 18244
rect 14599 18241 14611 18275
rect 14553 18235 14611 18241
rect 6892 18207 6950 18213
rect 6892 18173 6904 18207
rect 6938 18204 6950 18207
rect 7285 18207 7343 18213
rect 7285 18204 7297 18207
rect 6938 18176 7297 18204
rect 6938 18173 6950 18176
rect 6892 18167 6950 18173
rect 7285 18173 7297 18176
rect 7331 18173 7343 18207
rect 15140 18207 15198 18213
rect 15140 18204 15152 18207
rect 7285 18167 7343 18173
rect 14292 18176 15152 18204
rect 14292 18148 14320 18176
rect 15140 18173 15152 18176
rect 15186 18204 15198 18207
rect 15565 18207 15623 18213
rect 15565 18204 15577 18207
rect 15186 18176 15577 18204
rect 15186 18173 15198 18176
rect 15140 18167 15198 18173
rect 15565 18173 15577 18176
rect 15611 18173 15623 18207
rect 15565 18167 15623 18173
rect 8386 18136 8392 18148
rect 8347 18108 8392 18136
rect 8386 18096 8392 18108
rect 8444 18096 8450 18148
rect 8481 18139 8539 18145
rect 8481 18105 8493 18139
rect 8527 18105 8539 18139
rect 8481 18099 8539 18105
rect 10321 18139 10379 18145
rect 10321 18105 10333 18139
rect 10367 18136 10379 18139
rect 10870 18136 10876 18148
rect 10367 18108 10876 18136
rect 10367 18105 10379 18108
rect 10321 18099 10379 18105
rect 1535 18071 1593 18077
rect 1535 18037 1547 18071
rect 1581 18068 1593 18071
rect 2498 18068 2504 18080
rect 1581 18040 2504 18068
rect 1581 18037 1593 18040
rect 1535 18031 1593 18037
rect 2498 18028 2504 18040
rect 2556 18028 2562 18080
rect 5859 18071 5917 18077
rect 5859 18037 5871 18071
rect 5905 18068 5917 18071
rect 7926 18068 7932 18080
rect 5905 18040 7932 18068
rect 5905 18037 5917 18040
rect 5859 18031 5917 18037
rect 7926 18028 7932 18040
rect 7984 18028 7990 18080
rect 8202 18068 8208 18080
rect 8163 18040 8208 18068
rect 8202 18028 8208 18040
rect 8260 18068 8266 18080
rect 8496 18068 8524 18099
rect 10870 18096 10876 18108
rect 10928 18096 10934 18148
rect 10962 18096 10968 18148
rect 11020 18136 11026 18148
rect 12529 18139 12587 18145
rect 11020 18108 11065 18136
rect 11020 18096 11026 18108
rect 12529 18105 12541 18139
rect 12575 18136 12587 18139
rect 13081 18139 13139 18145
rect 13081 18136 13093 18139
rect 12575 18108 13093 18136
rect 12575 18105 12587 18108
rect 12529 18099 12587 18105
rect 13081 18105 13093 18108
rect 13127 18136 13139 18139
rect 13633 18139 13691 18145
rect 13633 18136 13645 18139
rect 13127 18108 13645 18136
rect 13127 18105 13139 18108
rect 13081 18099 13139 18105
rect 13633 18105 13645 18108
rect 13679 18105 13691 18139
rect 13633 18099 13691 18105
rect 13725 18139 13783 18145
rect 13725 18105 13737 18139
rect 13771 18105 13783 18139
rect 14274 18136 14280 18148
rect 14235 18108 14280 18136
rect 13725 18099 13783 18105
rect 8260 18040 8524 18068
rect 8260 18028 8266 18040
rect 13354 18028 13360 18080
rect 13412 18068 13418 18080
rect 13740 18068 13768 18099
rect 14274 18096 14280 18108
rect 14332 18096 14338 18148
rect 13412 18040 13768 18068
rect 13412 18028 13418 18040
rect 1104 17978 22816 18000
rect 1104 17926 8982 17978
rect 9034 17926 9046 17978
rect 9098 17926 9110 17978
rect 9162 17926 9174 17978
rect 9226 17926 16982 17978
rect 17034 17926 17046 17978
rect 17098 17926 17110 17978
rect 17162 17926 17174 17978
rect 17226 17926 22816 17978
rect 1104 17904 22816 17926
rect 2866 17824 2872 17876
rect 2924 17864 2930 17876
rect 8846 17864 8852 17876
rect 2924 17836 8852 17864
rect 2924 17824 2930 17836
rect 8846 17824 8852 17836
rect 8904 17824 8910 17876
rect 10244 17836 11744 17864
rect 10244 17808 10272 17836
rect 5721 17799 5779 17805
rect 5721 17765 5733 17799
rect 5767 17796 5779 17799
rect 5994 17796 6000 17808
rect 5767 17768 6000 17796
rect 5767 17765 5779 17768
rect 5721 17759 5779 17765
rect 5994 17756 6000 17768
rect 6052 17756 6058 17808
rect 8018 17796 8024 17808
rect 7979 17768 8024 17796
rect 8018 17756 8024 17768
rect 8076 17756 8082 17808
rect 10226 17796 10232 17808
rect 10139 17768 10232 17796
rect 10226 17756 10232 17768
rect 10284 17756 10290 17808
rect 10781 17799 10839 17805
rect 10781 17765 10793 17799
rect 10827 17796 10839 17799
rect 10870 17796 10876 17808
rect 10827 17768 10876 17796
rect 10827 17765 10839 17768
rect 10781 17759 10839 17765
rect 10870 17756 10876 17768
rect 10928 17756 10934 17808
rect 11716 17740 11744 17836
rect 13630 17796 13636 17808
rect 13591 17768 13636 17796
rect 13630 17756 13636 17768
rect 13688 17756 13694 17808
rect 14185 17799 14243 17805
rect 14185 17765 14197 17799
rect 14231 17796 14243 17799
rect 14274 17796 14280 17808
rect 14231 17768 14280 17796
rect 14231 17765 14243 17768
rect 14185 17759 14243 17765
rect 14274 17756 14280 17768
rect 14332 17756 14338 17808
rect 106 17688 112 17740
rect 164 17728 170 17740
rect 1432 17731 1490 17737
rect 1432 17728 1444 17731
rect 164 17700 1444 17728
rect 164 17688 170 17700
rect 1432 17697 1444 17700
rect 1478 17728 1490 17731
rect 1854 17728 1860 17740
rect 1478 17700 1860 17728
rect 1478 17697 1490 17700
rect 1432 17691 1490 17697
rect 1854 17688 1860 17700
rect 1912 17688 1918 17740
rect 2774 17728 2780 17740
rect 2735 17700 2780 17728
rect 2774 17688 2780 17700
rect 2832 17688 2838 17740
rect 11698 17728 11704 17740
rect 11659 17700 11704 17728
rect 11698 17688 11704 17700
rect 11756 17688 11762 17740
rect 15378 17737 15384 17740
rect 15356 17731 15384 17737
rect 15356 17728 15368 17731
rect 15291 17700 15368 17728
rect 15356 17697 15368 17700
rect 15436 17728 15442 17740
rect 20070 17728 20076 17740
rect 15436 17700 20076 17728
rect 15356 17691 15384 17697
rect 15378 17688 15384 17691
rect 15436 17688 15442 17700
rect 20070 17688 20076 17700
rect 20128 17688 20134 17740
rect 20968 17731 21026 17737
rect 20968 17697 20980 17731
rect 21014 17728 21026 17731
rect 21266 17728 21272 17740
rect 21014 17700 21272 17728
rect 21014 17697 21026 17700
rect 20968 17691 21026 17697
rect 21266 17688 21272 17700
rect 21324 17688 21330 17740
rect 5626 17660 5632 17672
rect 5587 17632 5632 17660
rect 5626 17620 5632 17632
rect 5684 17620 5690 17672
rect 5902 17660 5908 17672
rect 5863 17632 5908 17660
rect 5902 17620 5908 17632
rect 5960 17620 5966 17672
rect 7926 17660 7932 17672
rect 7887 17632 7932 17660
rect 7926 17620 7932 17632
rect 7984 17620 7990 17672
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17660 8631 17663
rect 8662 17660 8668 17672
rect 8619 17632 8668 17660
rect 8619 17629 8631 17632
rect 8573 17623 8631 17629
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 10134 17660 10140 17672
rect 10095 17632 10140 17660
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 10778 17620 10784 17672
rect 10836 17660 10842 17672
rect 11609 17663 11667 17669
rect 11609 17660 11621 17663
rect 10836 17632 11621 17660
rect 10836 17620 10842 17632
rect 11609 17629 11621 17632
rect 11655 17629 11667 17663
rect 13538 17660 13544 17672
rect 13499 17632 13544 17660
rect 11609 17623 11667 17629
rect 13538 17620 13544 17632
rect 13596 17620 13602 17672
rect 13262 17592 13268 17604
rect 13223 17564 13268 17592
rect 13262 17552 13268 17564
rect 13320 17592 13326 17604
rect 13320 17564 13814 17592
rect 13320 17552 13326 17564
rect 1535 17527 1593 17533
rect 1535 17493 1547 17527
rect 1581 17524 1593 17527
rect 1670 17524 1676 17536
rect 1581 17496 1676 17524
rect 1581 17493 1593 17496
rect 1535 17487 1593 17493
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 2682 17524 2688 17536
rect 2643 17496 2688 17524
rect 2682 17484 2688 17496
rect 2740 17484 2746 17536
rect 5261 17527 5319 17533
rect 5261 17493 5273 17527
rect 5307 17524 5319 17527
rect 5350 17524 5356 17536
rect 5307 17496 5356 17524
rect 5307 17493 5319 17496
rect 5261 17487 5319 17493
rect 5350 17484 5356 17496
rect 5408 17484 5414 17536
rect 13786 17524 13814 17564
rect 15427 17527 15485 17533
rect 15427 17524 15439 17527
rect 13786 17496 15439 17524
rect 15427 17493 15439 17496
rect 15473 17493 15485 17527
rect 15427 17487 15485 17493
rect 19334 17484 19340 17536
rect 19392 17524 19398 17536
rect 21039 17527 21097 17533
rect 21039 17524 21051 17527
rect 19392 17496 21051 17524
rect 19392 17484 19398 17496
rect 21039 17493 21051 17496
rect 21085 17493 21097 17527
rect 21039 17487 21097 17493
rect 1104 17434 22816 17456
rect 1104 17382 4982 17434
rect 5034 17382 5046 17434
rect 5098 17382 5110 17434
rect 5162 17382 5174 17434
rect 5226 17382 12982 17434
rect 13034 17382 13046 17434
rect 13098 17382 13110 17434
rect 13162 17382 13174 17434
rect 13226 17382 20982 17434
rect 21034 17382 21046 17434
rect 21098 17382 21110 17434
rect 21162 17382 21174 17434
rect 21226 17382 22816 17434
rect 1104 17360 22816 17382
rect 1854 17320 1860 17332
rect 1815 17292 1860 17320
rect 1854 17280 1860 17292
rect 1912 17280 1918 17332
rect 8202 17320 8208 17332
rect 8163 17292 8208 17320
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 10045 17323 10103 17329
rect 10045 17289 10057 17323
rect 10091 17320 10103 17323
rect 10226 17320 10232 17332
rect 10091 17292 10232 17320
rect 10091 17289 10103 17292
rect 10045 17283 10103 17289
rect 10226 17280 10232 17292
rect 10284 17320 10290 17332
rect 10502 17320 10508 17332
rect 10284 17292 10508 17320
rect 10284 17280 10290 17292
rect 10502 17280 10508 17292
rect 10560 17280 10566 17332
rect 11698 17320 11704 17332
rect 11659 17292 11704 17320
rect 11698 17280 11704 17292
rect 11756 17280 11762 17332
rect 15378 17320 15384 17332
rect 15339 17292 15384 17320
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 20993 17323 21051 17329
rect 20993 17289 21005 17323
rect 21039 17320 21051 17323
rect 21266 17320 21272 17332
rect 21039 17292 21272 17320
rect 21039 17289 21051 17292
rect 20993 17283 21051 17289
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 7926 17212 7932 17264
rect 7984 17252 7990 17264
rect 8941 17255 8999 17261
rect 8941 17252 8953 17255
rect 7984 17224 8953 17252
rect 7984 17212 7990 17224
rect 8941 17221 8953 17224
rect 8987 17221 8999 17255
rect 8941 17215 8999 17221
rect 2498 17144 2504 17196
rect 2556 17184 2562 17196
rect 2685 17187 2743 17193
rect 2685 17184 2697 17187
rect 2556 17156 2697 17184
rect 2556 17144 2562 17156
rect 2685 17153 2697 17156
rect 2731 17153 2743 17187
rect 3142 17184 3148 17196
rect 3103 17156 3148 17184
rect 2685 17147 2743 17153
rect 3142 17144 3148 17156
rect 3200 17184 3206 17196
rect 4617 17187 4675 17193
rect 4617 17184 4629 17187
rect 3200 17156 4629 17184
rect 3200 17144 3206 17156
rect 4617 17153 4629 17156
rect 4663 17184 4675 17187
rect 5261 17187 5319 17193
rect 5261 17184 5273 17187
rect 4663 17156 5273 17184
rect 4663 17153 4675 17156
rect 4617 17147 4675 17153
rect 5261 17153 5273 17156
rect 5307 17153 5319 17187
rect 5902 17184 5908 17196
rect 5863 17156 5908 17184
rect 5261 17147 5319 17153
rect 5902 17144 5908 17156
rect 5960 17144 5966 17196
rect 8110 17144 8116 17196
rect 8168 17184 8174 17196
rect 9585 17187 9643 17193
rect 9585 17184 9597 17187
rect 8168 17156 9597 17184
rect 8168 17144 8174 17156
rect 9585 17153 9597 17156
rect 9631 17184 9643 17187
rect 10134 17184 10140 17196
rect 9631 17156 10140 17184
rect 9631 17153 9643 17156
rect 9585 17147 9643 17153
rect 10134 17144 10140 17156
rect 10192 17144 10198 17196
rect 10870 17184 10876 17196
rect 10831 17156 10876 17184
rect 10870 17144 10876 17156
rect 10928 17144 10934 17196
rect 13262 17184 13268 17196
rect 13223 17156 13268 17184
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 13538 17184 13544 17196
rect 13499 17156 13544 17184
rect 13538 17144 13544 17156
rect 13596 17144 13602 17196
rect 1461 17116 1467 17128
rect 1422 17088 1467 17116
rect 1461 17076 1467 17088
rect 1519 17116 1525 17128
rect 2225 17119 2283 17125
rect 2225 17116 2237 17119
rect 1519 17088 2237 17116
rect 1519 17076 1525 17088
rect 2225 17085 2237 17088
rect 2271 17085 2283 17119
rect 2225 17079 2283 17085
rect 7469 17119 7527 17125
rect 7469 17085 7481 17119
rect 7515 17116 7527 17119
rect 7837 17119 7895 17125
rect 7837 17116 7849 17119
rect 7515 17088 7849 17116
rect 7515 17085 7527 17088
rect 7469 17079 7527 17085
rect 7837 17085 7849 17088
rect 7883 17116 7895 17119
rect 8018 17116 8024 17128
rect 7883 17088 8024 17116
rect 7883 17085 7895 17088
rect 7837 17079 7895 17085
rect 8018 17076 8024 17088
rect 8076 17116 8082 17128
rect 8386 17116 8392 17128
rect 8076 17088 8392 17116
rect 8076 17076 8082 17088
rect 8386 17076 8392 17088
rect 8444 17076 8450 17128
rect 2774 17008 2780 17060
rect 2832 17048 2838 17060
rect 3605 17051 3663 17057
rect 3605 17048 3617 17051
rect 2832 17020 3617 17048
rect 2832 17008 2838 17020
rect 3605 17017 3617 17020
rect 3651 17048 3663 17051
rect 3786 17048 3792 17060
rect 3651 17020 3792 17048
rect 3651 17017 3663 17020
rect 3605 17011 3663 17017
rect 3786 17008 3792 17020
rect 3844 17048 3850 17060
rect 3973 17051 4031 17057
rect 3973 17048 3985 17051
rect 3844 17020 3985 17048
rect 3844 17008 3850 17020
rect 3973 17017 3985 17020
rect 4019 17017 4031 17051
rect 5350 17048 5356 17060
rect 5311 17020 5356 17048
rect 3973 17011 4031 17017
rect 5350 17008 5356 17020
rect 5408 17008 5414 17060
rect 5626 17008 5632 17060
rect 5684 17048 5690 17060
rect 6825 17051 6883 17057
rect 6825 17048 6837 17051
rect 5684 17020 6837 17048
rect 5684 17008 5690 17020
rect 6825 17017 6837 17020
rect 6871 17017 6883 17051
rect 6825 17011 6883 17017
rect 10318 17008 10324 17060
rect 10376 17048 10382 17060
rect 10597 17051 10655 17057
rect 10597 17048 10609 17051
rect 10376 17020 10609 17048
rect 10376 17008 10382 17020
rect 10597 17017 10609 17020
rect 10643 17017 10655 17051
rect 10597 17011 10655 17017
rect 10689 17051 10747 17057
rect 10689 17017 10701 17051
rect 10735 17048 10747 17051
rect 10778 17048 10784 17060
rect 10735 17020 10784 17048
rect 10735 17017 10747 17020
rect 10689 17011 10747 17017
rect 1535 16983 1593 16989
rect 1535 16949 1547 16983
rect 1581 16980 1593 16983
rect 1854 16980 1860 16992
rect 1581 16952 1860 16980
rect 1581 16949 1593 16952
rect 1535 16943 1593 16949
rect 1854 16940 1860 16952
rect 1912 16940 1918 16992
rect 5077 16983 5135 16989
rect 5077 16949 5089 16983
rect 5123 16980 5135 16983
rect 5644 16980 5672 17008
rect 5123 16952 5672 16980
rect 5123 16949 5135 16952
rect 5077 16943 5135 16949
rect 5994 16940 6000 16992
rect 6052 16980 6058 16992
rect 6181 16983 6239 16989
rect 6181 16980 6193 16983
rect 6052 16952 6193 16980
rect 6052 16940 6058 16952
rect 6181 16949 6193 16952
rect 6227 16949 6239 16983
rect 6181 16943 6239 16949
rect 10413 16983 10471 16989
rect 10413 16949 10425 16983
rect 10459 16980 10471 16983
rect 10704 16980 10732 17011
rect 10778 17008 10784 17020
rect 10836 17008 10842 17060
rect 13357 17051 13415 17057
rect 13357 17017 13369 17051
rect 13403 17017 13415 17051
rect 13357 17011 13415 17017
rect 10459 16952 10732 16980
rect 10459 16949 10471 16952
rect 10413 16943 10471 16949
rect 12802 16940 12808 16992
rect 12860 16980 12866 16992
rect 12989 16983 13047 16989
rect 12989 16980 13001 16983
rect 12860 16952 13001 16980
rect 12860 16940 12866 16952
rect 12989 16949 13001 16952
rect 13035 16980 13047 16983
rect 13372 16980 13400 17011
rect 13035 16952 13400 16980
rect 13035 16949 13047 16952
rect 12989 16943 13047 16949
rect 13446 16940 13452 16992
rect 13504 16980 13510 16992
rect 13630 16980 13636 16992
rect 13504 16952 13636 16980
rect 13504 16940 13510 16952
rect 13630 16940 13636 16952
rect 13688 16980 13694 16992
rect 14185 16983 14243 16989
rect 14185 16980 14197 16983
rect 13688 16952 14197 16980
rect 13688 16940 13694 16952
rect 14185 16949 14197 16952
rect 14231 16949 14243 16983
rect 14185 16943 14243 16949
rect 1104 16890 22816 16912
rect 1104 16838 8982 16890
rect 9034 16838 9046 16890
rect 9098 16838 9110 16890
rect 9162 16838 9174 16890
rect 9226 16838 16982 16890
rect 17034 16838 17046 16890
rect 17098 16838 17110 16890
rect 17162 16838 17174 16890
rect 17226 16838 22816 16890
rect 1104 16816 22816 16838
rect 2498 16736 2504 16788
rect 2556 16776 2562 16788
rect 3421 16779 3479 16785
rect 3421 16776 3433 16779
rect 2556 16748 3433 16776
rect 2556 16736 2562 16748
rect 3421 16745 3433 16748
rect 3467 16745 3479 16779
rect 8386 16776 8392 16788
rect 8347 16748 8392 16776
rect 3421 16739 3479 16745
rect 8386 16736 8392 16748
rect 8444 16736 8450 16788
rect 13538 16776 13544 16788
rect 13372 16748 13544 16776
rect 2593 16711 2651 16717
rect 2593 16677 2605 16711
rect 2639 16708 2651 16711
rect 2682 16708 2688 16720
rect 2639 16680 2688 16708
rect 2639 16677 2651 16680
rect 2593 16671 2651 16677
rect 2682 16668 2688 16680
rect 2740 16668 2746 16720
rect 3142 16708 3148 16720
rect 3103 16680 3148 16708
rect 3142 16668 3148 16680
rect 3200 16668 3206 16720
rect 5994 16708 6000 16720
rect 5955 16680 6000 16708
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 7831 16711 7889 16717
rect 7831 16677 7843 16711
rect 7877 16708 7889 16711
rect 8018 16708 8024 16720
rect 7877 16680 8024 16708
rect 7877 16677 7889 16680
rect 7831 16671 7889 16677
rect 8018 16668 8024 16680
rect 8076 16668 8082 16720
rect 10410 16708 10416 16720
rect 9968 16680 10416 16708
rect 1464 16643 1522 16649
rect 1464 16609 1476 16643
rect 1510 16640 1522 16643
rect 1946 16640 1952 16652
rect 1510 16612 1952 16640
rect 1510 16609 1522 16612
rect 1464 16603 1522 16609
rect 1946 16600 1952 16612
rect 2004 16600 2010 16652
rect 5350 16640 5356 16652
rect 5311 16612 5356 16640
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 9968 16649 9996 16680
rect 10410 16668 10416 16680
rect 10468 16668 10474 16720
rect 11882 16668 11888 16720
rect 11940 16708 11946 16720
rect 13372 16717 13400 16748
rect 13538 16736 13544 16748
rect 13596 16776 13602 16788
rect 13633 16779 13691 16785
rect 13633 16776 13645 16779
rect 13596 16748 13645 16776
rect 13596 16736 13602 16748
rect 13633 16745 13645 16748
rect 13679 16745 13691 16779
rect 13633 16739 13691 16745
rect 12805 16711 12863 16717
rect 12805 16708 12817 16711
rect 11940 16680 12817 16708
rect 11940 16668 11946 16680
rect 12805 16677 12817 16680
rect 12851 16677 12863 16711
rect 12805 16671 12863 16677
rect 13357 16711 13415 16717
rect 13357 16677 13369 16711
rect 13403 16677 13415 16711
rect 13357 16671 13415 16677
rect 9953 16643 10011 16649
rect 9953 16609 9965 16643
rect 9999 16609 10011 16643
rect 10134 16640 10140 16652
rect 10095 16612 10140 16640
rect 9953 16603 10011 16609
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 20968 16643 21026 16649
rect 20968 16609 20980 16643
rect 21014 16640 21026 16643
rect 21266 16640 21272 16652
rect 21014 16612 21272 16640
rect 21014 16609 21026 16612
rect 20968 16603 21026 16609
rect 21266 16600 21272 16612
rect 21324 16600 21330 16652
rect 2222 16532 2228 16584
rect 2280 16572 2286 16584
rect 2501 16575 2559 16581
rect 2501 16572 2513 16575
rect 2280 16544 2513 16572
rect 2280 16532 2286 16544
rect 2501 16541 2513 16544
rect 2547 16541 2559 16575
rect 2501 16535 2559 16541
rect 7469 16575 7527 16581
rect 7469 16541 7481 16575
rect 7515 16572 7527 16575
rect 8386 16572 8392 16584
rect 7515 16544 8392 16572
rect 7515 16541 7527 16544
rect 7469 16535 7527 16541
rect 8386 16532 8392 16544
rect 8444 16532 8450 16584
rect 10226 16572 10232 16584
rect 10187 16544 10232 16572
rect 10226 16532 10232 16544
rect 10284 16532 10290 16584
rect 12710 16572 12716 16584
rect 12671 16544 12716 16572
rect 12710 16532 12716 16544
rect 12768 16532 12774 16584
rect 1535 16439 1593 16445
rect 1535 16405 1547 16439
rect 1581 16436 1593 16439
rect 1762 16436 1768 16448
rect 1581 16408 1768 16436
rect 1581 16405 1593 16408
rect 1535 16399 1593 16405
rect 1762 16396 1768 16408
rect 1820 16396 1826 16448
rect 7098 16436 7104 16448
rect 7059 16408 7104 16436
rect 7098 16396 7104 16408
rect 7156 16396 7162 16448
rect 10318 16396 10324 16448
rect 10376 16436 10382 16448
rect 10689 16439 10747 16445
rect 10689 16436 10701 16439
rect 10376 16408 10701 16436
rect 10376 16396 10382 16408
rect 10689 16405 10701 16408
rect 10735 16405 10747 16439
rect 10689 16399 10747 16405
rect 20438 16396 20444 16448
rect 20496 16436 20502 16448
rect 21039 16439 21097 16445
rect 21039 16436 21051 16439
rect 20496 16408 21051 16436
rect 20496 16396 20502 16408
rect 21039 16405 21051 16408
rect 21085 16405 21097 16439
rect 21039 16399 21097 16405
rect 1104 16346 22816 16368
rect 1104 16294 4982 16346
rect 5034 16294 5046 16346
rect 5098 16294 5110 16346
rect 5162 16294 5174 16346
rect 5226 16294 12982 16346
rect 13034 16294 13046 16346
rect 13098 16294 13110 16346
rect 13162 16294 13174 16346
rect 13226 16294 20982 16346
rect 21034 16294 21046 16346
rect 21098 16294 21110 16346
rect 21162 16294 21174 16346
rect 21226 16294 22816 16346
rect 1104 16272 22816 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 2409 16235 2467 16241
rect 2409 16201 2421 16235
rect 2455 16232 2467 16235
rect 2682 16232 2688 16244
rect 2455 16204 2688 16232
rect 2455 16201 2467 16204
rect 2409 16195 2467 16201
rect 2682 16192 2688 16204
rect 2740 16192 2746 16244
rect 3786 16232 3792 16244
rect 3747 16204 3792 16232
rect 3786 16192 3792 16204
rect 3844 16192 3850 16244
rect 5350 16192 5356 16244
rect 5408 16232 5414 16244
rect 5629 16235 5687 16241
rect 5629 16232 5641 16235
rect 5408 16204 5641 16232
rect 5408 16192 5414 16204
rect 5629 16201 5641 16204
rect 5675 16232 5687 16235
rect 5905 16235 5963 16241
rect 5905 16232 5917 16235
rect 5675 16204 5917 16232
rect 5675 16201 5687 16204
rect 5629 16195 5687 16201
rect 5905 16201 5917 16204
rect 5951 16201 5963 16235
rect 10502 16232 10508 16244
rect 10463 16204 10508 16232
rect 5905 16195 5963 16201
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 11882 16232 11888 16244
rect 11843 16204 11888 16232
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 12802 16192 12808 16244
rect 12860 16232 12866 16244
rect 14001 16235 14059 16241
rect 14001 16232 14013 16235
rect 12860 16204 14013 16232
rect 12860 16192 12866 16204
rect 14001 16201 14013 16204
rect 14047 16201 14059 16235
rect 14001 16195 14059 16201
rect 20993 16235 21051 16241
rect 20993 16201 21005 16235
rect 21039 16232 21051 16235
rect 21266 16232 21272 16244
rect 21039 16204 21272 16232
rect 21039 16201 21051 16204
rect 20993 16195 21051 16201
rect 21266 16192 21272 16204
rect 21324 16192 21330 16244
rect 7374 16096 7380 16108
rect 7335 16068 7380 16096
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 11900 16096 11928 16192
rect 13446 16164 13452 16176
rect 13407 16136 13452 16164
rect 13446 16124 13452 16136
rect 13504 16124 13510 16176
rect 14277 16099 14335 16105
rect 14277 16096 14289 16099
rect 11900 16068 14289 16096
rect 14277 16065 14289 16068
rect 14323 16065 14335 16099
rect 14277 16059 14335 16065
rect 1394 16028 1400 16040
rect 1355 16000 1400 16028
rect 1394 15988 1400 16000
rect 1452 15988 1458 16040
rect 2866 16028 2872 16040
rect 2827 16000 2872 16028
rect 2866 15988 2872 16000
rect 2924 15988 2930 16040
rect 4706 16028 4712 16040
rect 4667 16000 4712 16028
rect 4706 15988 4712 16000
rect 4764 15988 4770 16040
rect 9585 16031 9643 16037
rect 9585 15997 9597 16031
rect 9631 16028 9643 16031
rect 9766 16028 9772 16040
rect 9631 16000 9772 16028
rect 9631 15997 9643 16000
rect 9585 15991 9643 15997
rect 9766 15988 9772 16000
rect 9824 16028 9830 16040
rect 10781 16031 10839 16037
rect 10781 16028 10793 16031
rect 9824 16000 10793 16028
rect 9824 15988 9830 16000
rect 10781 15997 10793 16000
rect 10827 15997 10839 16031
rect 10781 15991 10839 15997
rect 12529 16031 12587 16037
rect 12529 15997 12541 16031
rect 12575 16028 12587 16031
rect 13262 16028 13268 16040
rect 12575 16000 13268 16028
rect 12575 15997 12587 16000
rect 12529 15991 12587 15997
rect 13262 15988 13268 16000
rect 13320 16028 13326 16040
rect 13725 16031 13783 16037
rect 13725 16028 13737 16031
rect 13320 16000 13737 16028
rect 13320 15988 13326 16000
rect 13725 15997 13737 16000
rect 13771 15997 13783 16031
rect 13725 15991 13783 15997
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 16028 14059 16031
rect 14185 16031 14243 16037
rect 14185 16028 14197 16031
rect 14047 16000 14197 16028
rect 14047 15997 14059 16000
rect 14001 15991 14059 15997
rect 14185 15997 14197 16000
rect 14231 16028 14243 16031
rect 14369 16031 14427 16037
rect 14369 16028 14381 16031
rect 14231 16000 14381 16028
rect 14231 15997 14243 16000
rect 14185 15991 14243 15997
rect 14369 15997 14381 16000
rect 14415 15997 14427 16031
rect 14369 15991 14427 15997
rect 2774 15960 2780 15972
rect 2735 15932 2780 15960
rect 2774 15920 2780 15932
rect 2832 15960 2838 15972
rect 3190 15963 3248 15969
rect 3190 15960 3202 15963
rect 2832 15932 3202 15960
rect 2832 15920 2838 15932
rect 3190 15929 3202 15932
rect 3236 15960 3248 15963
rect 4525 15963 4583 15969
rect 4525 15960 4537 15963
rect 3236 15932 4537 15960
rect 3236 15929 3248 15932
rect 3190 15923 3248 15929
rect 4525 15929 4537 15932
rect 4571 15960 4583 15963
rect 5030 15963 5088 15969
rect 5030 15960 5042 15963
rect 4571 15932 5042 15960
rect 4571 15929 4583 15932
rect 4525 15923 4583 15929
rect 5030 15929 5042 15932
rect 5076 15929 5088 15963
rect 7098 15960 7104 15972
rect 7059 15932 7104 15960
rect 5030 15923 5088 15929
rect 7098 15920 7104 15932
rect 7156 15920 7162 15972
rect 7193 15963 7251 15969
rect 7193 15929 7205 15963
rect 7239 15929 7251 15963
rect 9401 15963 9459 15969
rect 9401 15960 9413 15963
rect 7193 15923 7251 15929
rect 8036 15932 9413 15960
rect 1946 15892 1952 15904
rect 1907 15864 1952 15892
rect 1946 15852 1952 15864
rect 2004 15852 2010 15904
rect 2222 15852 2228 15904
rect 2280 15892 2286 15904
rect 4065 15895 4123 15901
rect 4065 15892 4077 15895
rect 2280 15864 4077 15892
rect 2280 15852 2286 15864
rect 4065 15861 4077 15864
rect 4111 15861 4123 15895
rect 6546 15892 6552 15904
rect 6507 15864 6552 15892
rect 4065 15855 4123 15861
rect 6546 15852 6552 15864
rect 6604 15892 6610 15904
rect 7208 15892 7236 15923
rect 8036 15904 8064 15932
rect 9401 15929 9413 15932
rect 9447 15960 9459 15963
rect 9906 15963 9964 15969
rect 9906 15960 9918 15963
rect 9447 15932 9918 15960
rect 9447 15929 9459 15932
rect 9401 15923 9459 15929
rect 9906 15929 9918 15932
rect 9952 15960 9964 15963
rect 10042 15960 10048 15972
rect 9952 15932 10048 15960
rect 9952 15929 9964 15932
rect 9906 15923 9964 15929
rect 10042 15920 10048 15932
rect 10100 15920 10106 15972
rect 12850 15963 12908 15969
rect 12850 15929 12862 15963
rect 12896 15929 12908 15963
rect 12850 15923 12908 15929
rect 8018 15892 8024 15904
rect 6604 15864 7236 15892
rect 7979 15864 8024 15892
rect 6604 15852 6610 15864
rect 8018 15852 8024 15864
rect 8076 15852 8082 15904
rect 8386 15892 8392 15904
rect 8347 15864 8392 15892
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 9125 15895 9183 15901
rect 9125 15861 9137 15895
rect 9171 15892 9183 15895
rect 10410 15892 10416 15904
rect 9171 15864 10416 15892
rect 9171 15861 9183 15864
rect 9125 15855 9183 15861
rect 10410 15852 10416 15864
rect 10468 15852 10474 15904
rect 12250 15892 12256 15904
rect 12211 15864 12256 15892
rect 12250 15852 12256 15864
rect 12308 15892 12314 15904
rect 12865 15892 12893 15923
rect 12308 15864 12893 15892
rect 12308 15852 12314 15864
rect 1104 15802 22816 15824
rect 1104 15750 8982 15802
rect 9034 15750 9046 15802
rect 9098 15750 9110 15802
rect 9162 15750 9174 15802
rect 9226 15750 16982 15802
rect 17034 15750 17046 15802
rect 17098 15750 17110 15802
rect 17162 15750 17174 15802
rect 17226 15750 22816 15802
rect 1104 15728 22816 15750
rect 1394 15648 1400 15700
rect 1452 15688 1458 15700
rect 1535 15691 1593 15697
rect 1535 15688 1547 15691
rect 1452 15660 1547 15688
rect 1452 15648 1458 15660
rect 1535 15657 1547 15660
rect 1581 15688 1593 15691
rect 1857 15691 1915 15697
rect 1857 15688 1869 15691
rect 1581 15660 1869 15688
rect 1581 15657 1593 15660
rect 1535 15651 1593 15657
rect 1857 15657 1869 15660
rect 1903 15657 1915 15691
rect 1857 15651 1915 15657
rect 2685 15691 2743 15697
rect 2685 15657 2697 15691
rect 2731 15688 2743 15691
rect 2866 15688 2872 15700
rect 2731 15660 2872 15688
rect 2731 15657 2743 15660
rect 2685 15651 2743 15657
rect 2866 15648 2872 15660
rect 2924 15688 2930 15700
rect 3421 15691 3479 15697
rect 3421 15688 3433 15691
rect 2924 15660 3433 15688
rect 2924 15648 2930 15660
rect 3421 15657 3433 15660
rect 3467 15657 3479 15691
rect 3421 15651 3479 15657
rect 7098 15648 7104 15700
rect 7156 15688 7162 15700
rect 8573 15691 8631 15697
rect 8573 15688 8585 15691
rect 7156 15660 8585 15688
rect 7156 15648 7162 15660
rect 8573 15657 8585 15660
rect 8619 15657 8631 15691
rect 8573 15651 8631 15657
rect 9953 15691 10011 15697
rect 9953 15657 9965 15691
rect 9999 15688 10011 15691
rect 10134 15688 10140 15700
rect 9999 15660 10140 15688
rect 9999 15657 10011 15660
rect 9953 15651 10011 15657
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 10962 15688 10968 15700
rect 10923 15660 10968 15688
rect 10962 15648 10968 15660
rect 11020 15648 11026 15700
rect 12802 15648 12808 15700
rect 12860 15688 12866 15700
rect 13081 15691 13139 15697
rect 13081 15688 13093 15691
rect 12860 15660 13093 15688
rect 12860 15648 12866 15660
rect 13081 15657 13093 15660
rect 13127 15657 13139 15691
rect 13081 15651 13139 15657
rect 6181 15623 6239 15629
rect 6181 15589 6193 15623
rect 6227 15620 6239 15623
rect 6546 15620 6552 15632
rect 6227 15592 6552 15620
rect 6227 15589 6239 15592
rect 6181 15583 6239 15589
rect 6546 15580 6552 15592
rect 6604 15580 6610 15632
rect 7190 15620 7196 15632
rect 7151 15592 7196 15620
rect 7190 15580 7196 15592
rect 7248 15580 7254 15632
rect 10407 15623 10465 15629
rect 10407 15589 10419 15623
rect 10453 15589 10465 15623
rect 10407 15583 10465 15589
rect 1464 15555 1522 15561
rect 1464 15521 1476 15555
rect 1510 15521 1522 15555
rect 2682 15552 2688 15564
rect 2643 15524 2688 15552
rect 1464 15515 1522 15521
rect 1479 15484 1507 15515
rect 2682 15512 2688 15524
rect 2740 15512 2746 15564
rect 2958 15552 2964 15564
rect 2919 15524 2964 15552
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 6086 15552 6092 15564
rect 6047 15524 6092 15552
rect 6086 15512 6092 15524
rect 6144 15512 6150 15564
rect 10045 15555 10103 15561
rect 10045 15521 10057 15555
rect 10091 15552 10103 15555
rect 10226 15552 10232 15564
rect 10091 15524 10232 15552
rect 10091 15521 10103 15524
rect 10045 15515 10103 15521
rect 10226 15512 10232 15524
rect 10284 15512 10290 15564
rect 1578 15484 1584 15496
rect 1479 15456 1584 15484
rect 1578 15444 1584 15456
rect 1636 15484 1642 15496
rect 7098 15484 7104 15496
rect 1636 15456 4154 15484
rect 7059 15456 7104 15484
rect 1636 15444 1642 15456
rect 4126 15416 4154 15456
rect 7098 15444 7104 15456
rect 7156 15444 7162 15496
rect 7374 15484 7380 15496
rect 7287 15456 7380 15484
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 7392 15416 7420 15444
rect 4126 15388 7420 15416
rect 10042 15376 10048 15428
rect 10100 15416 10106 15428
rect 10422 15416 10450 15583
rect 12250 15580 12256 15632
rect 12308 15620 12314 15632
rect 12482 15623 12540 15629
rect 12482 15620 12494 15623
rect 12308 15592 12494 15620
rect 12308 15580 12314 15592
rect 12482 15589 12494 15592
rect 12528 15589 12540 15623
rect 12482 15583 12540 15589
rect 12158 15484 12164 15496
rect 12119 15456 12164 15484
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 10100 15388 10450 15416
rect 10100 15376 10106 15388
rect 4706 15348 4712 15360
rect 4667 15320 4712 15348
rect 4706 15308 4712 15320
rect 4764 15308 4770 15360
rect 6822 15348 6828 15360
rect 6783 15320 6828 15348
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 11146 15308 11152 15360
rect 11204 15348 11210 15360
rect 12710 15348 12716 15360
rect 11204 15320 12716 15348
rect 11204 15308 11210 15320
rect 12710 15308 12716 15320
rect 12768 15348 12774 15360
rect 13357 15351 13415 15357
rect 13357 15348 13369 15351
rect 12768 15320 13369 15348
rect 12768 15308 12774 15320
rect 13357 15317 13369 15320
rect 13403 15317 13415 15351
rect 13357 15311 13415 15317
rect 1104 15258 22816 15280
rect 1104 15206 4982 15258
rect 5034 15206 5046 15258
rect 5098 15206 5110 15258
rect 5162 15206 5174 15258
rect 5226 15206 12982 15258
rect 13034 15206 13046 15258
rect 13098 15206 13110 15258
rect 13162 15206 13174 15258
rect 13226 15206 20982 15258
rect 21034 15206 21046 15258
rect 21098 15206 21110 15258
rect 21162 15206 21174 15258
rect 21226 15206 22816 15258
rect 1104 15184 22816 15206
rect 2958 15104 2964 15156
rect 3016 15144 3022 15156
rect 3145 15147 3203 15153
rect 3145 15144 3157 15147
rect 3016 15116 3157 15144
rect 3016 15104 3022 15116
rect 3145 15113 3157 15116
rect 3191 15144 3203 15147
rect 3605 15147 3663 15153
rect 3605 15144 3617 15147
rect 3191 15116 3617 15144
rect 3191 15113 3203 15116
rect 3145 15107 3203 15113
rect 3605 15113 3617 15116
rect 3651 15113 3663 15147
rect 3605 15107 3663 15113
rect 5537 15147 5595 15153
rect 5537 15113 5549 15147
rect 5583 15144 5595 15147
rect 6086 15144 6092 15156
rect 5583 15116 6092 15144
rect 5583 15113 5595 15116
rect 5537 15107 5595 15113
rect 1673 14943 1731 14949
rect 1673 14909 1685 14943
rect 1719 14940 1731 14943
rect 1857 14943 1915 14949
rect 1857 14940 1869 14943
rect 1719 14912 1869 14940
rect 1719 14909 1731 14912
rect 1673 14903 1731 14909
rect 1857 14909 1869 14912
rect 1903 14940 1915 14943
rect 2130 14940 2136 14952
rect 1903 14912 2136 14940
rect 1903 14909 1915 14912
rect 1857 14903 1915 14909
rect 2130 14900 2136 14912
rect 2188 14900 2194 14952
rect 3620 14872 3648 15107
rect 6086 15104 6092 15116
rect 6144 15144 6150 15156
rect 6273 15147 6331 15153
rect 6273 15144 6285 15147
rect 6144 15116 6285 15144
rect 6144 15104 6150 15116
rect 6273 15113 6285 15116
rect 6319 15144 6331 15147
rect 7190 15144 7196 15156
rect 6319 15116 7196 15144
rect 6319 15113 6331 15116
rect 6273 15107 6331 15113
rect 7190 15104 7196 15116
rect 7248 15144 7254 15156
rect 7745 15147 7803 15153
rect 7745 15144 7757 15147
rect 7248 15116 7757 15144
rect 7248 15104 7254 15116
rect 7745 15113 7757 15116
rect 7791 15113 7803 15147
rect 7745 15107 7803 15113
rect 8938 15104 8944 15156
rect 8996 15144 9002 15156
rect 15611 15147 15669 15153
rect 15611 15144 15623 15147
rect 8996 15116 15623 15144
rect 8996 15104 9002 15116
rect 15611 15113 15623 15116
rect 15657 15113 15669 15147
rect 15611 15107 15669 15113
rect 10226 15036 10232 15088
rect 10284 15076 10290 15088
rect 10597 15079 10655 15085
rect 10597 15076 10609 15079
rect 10284 15048 10609 15076
rect 10284 15036 10290 15048
rect 10597 15045 10609 15048
rect 10643 15045 10655 15079
rect 14550 15076 14556 15088
rect 14511 15048 14556 15076
rect 10597 15039 10655 15045
rect 14550 15036 14556 15048
rect 14608 15036 14614 15088
rect 4706 15008 4712 15020
rect 4667 14980 4712 15008
rect 4706 14968 4712 14980
rect 4764 14968 4770 15020
rect 9766 15008 9772 15020
rect 9727 14980 9772 15008
rect 9766 14968 9772 14980
rect 9824 14968 9830 15020
rect 10042 14968 10048 15020
rect 10100 15008 10106 15020
rect 10321 15011 10379 15017
rect 10321 15008 10333 15011
rect 10100 14980 10333 15008
rect 10100 14968 10106 14980
rect 10321 14977 10333 14980
rect 10367 15008 10379 15011
rect 12250 15008 12256 15020
rect 10367 14980 12256 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 12250 14968 12256 14980
rect 12308 14968 12314 15020
rect 13173 15011 13231 15017
rect 13173 14977 13185 15011
rect 13219 15008 13231 15011
rect 13262 15008 13268 15020
rect 13219 14980 13268 15008
rect 13219 14977 13231 14980
rect 13173 14971 13231 14977
rect 13262 14968 13268 14980
rect 13320 14968 13326 15020
rect 4065 14943 4123 14949
rect 4065 14909 4077 14943
rect 4111 14940 4123 14943
rect 4430 14940 4436 14952
rect 4111 14912 4436 14940
rect 4111 14909 4123 14912
rect 4065 14903 4123 14909
rect 4430 14900 4436 14912
rect 4488 14900 4494 14952
rect 4614 14940 4620 14952
rect 4575 14912 4620 14940
rect 4614 14900 4620 14912
rect 4672 14900 4678 14952
rect 5626 14900 5632 14952
rect 5684 14940 5690 14952
rect 6822 14940 6828 14952
rect 5684 14912 6828 14940
rect 5684 14900 5690 14912
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 9217 14943 9275 14949
rect 9217 14909 9229 14943
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 4632 14872 4660 14900
rect 3620 14844 4660 14872
rect 7146 14875 7204 14881
rect 7146 14841 7158 14875
rect 7192 14872 7204 14875
rect 8018 14872 8024 14884
rect 7192 14844 8024 14872
rect 7192 14841 7204 14844
rect 7146 14835 7204 14841
rect 2038 14804 2044 14816
rect 1999 14776 2044 14804
rect 2038 14764 2044 14776
rect 2096 14764 2102 14816
rect 2682 14764 2688 14816
rect 2740 14804 2746 14816
rect 2777 14807 2835 14813
rect 2777 14804 2789 14807
rect 2740 14776 2789 14804
rect 2740 14764 2746 14776
rect 2777 14773 2789 14776
rect 2823 14773 2835 14807
rect 2777 14767 2835 14773
rect 6270 14764 6276 14816
rect 6328 14804 6334 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 6328 14776 6561 14804
rect 6328 14764 6334 14776
rect 6549 14773 6561 14776
rect 6595 14804 6607 14807
rect 7161 14804 7189 14835
rect 8018 14832 8024 14844
rect 8076 14832 8082 14884
rect 6595 14776 7189 14804
rect 9125 14807 9183 14813
rect 6595 14773 6607 14776
rect 6549 14767 6607 14773
rect 9125 14773 9137 14807
rect 9171 14804 9183 14807
rect 9232 14804 9260 14903
rect 9306 14900 9312 14952
rect 9364 14940 9370 14952
rect 9677 14943 9735 14949
rect 9677 14940 9689 14943
rect 9364 14912 9689 14940
rect 9364 14900 9370 14912
rect 9677 14909 9689 14912
rect 9723 14940 9735 14943
rect 10134 14940 10140 14952
rect 9723 14912 10140 14940
rect 9723 14909 9735 14912
rect 9677 14903 9735 14909
rect 10134 14900 10140 14912
rect 10192 14900 10198 14952
rect 11517 14943 11575 14949
rect 11517 14909 11529 14943
rect 11563 14940 11575 14943
rect 12158 14940 12164 14952
rect 11563 14912 12164 14940
rect 11563 14909 11575 14912
rect 11517 14903 11575 14909
rect 12158 14900 12164 14912
rect 12216 14900 12222 14952
rect 12434 14940 12440 14952
rect 12395 14912 12440 14940
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 12544 14912 12909 14940
rect 11885 14875 11943 14881
rect 11885 14841 11897 14875
rect 11931 14872 11943 14875
rect 11974 14872 11980 14884
rect 11931 14844 11980 14872
rect 11931 14841 11943 14844
rect 11885 14835 11943 14841
rect 11974 14832 11980 14844
rect 12032 14872 12038 14884
rect 12544 14872 12572 14912
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 14366 14940 14372 14952
rect 14279 14912 14372 14940
rect 12897 14903 12955 14909
rect 14366 14900 14372 14912
rect 14424 14940 14430 14952
rect 14921 14943 14979 14949
rect 14921 14940 14933 14943
rect 14424 14912 14933 14940
rect 14424 14900 14430 14912
rect 14921 14909 14933 14912
rect 14967 14909 14979 14943
rect 14921 14903 14979 14909
rect 15540 14943 15598 14949
rect 15540 14909 15552 14943
rect 15586 14940 15598 14943
rect 15654 14940 15660 14952
rect 15586 14912 15660 14940
rect 15586 14909 15598 14912
rect 15540 14903 15598 14909
rect 15654 14900 15660 14912
rect 15712 14940 15718 14952
rect 15933 14943 15991 14949
rect 15933 14940 15945 14943
rect 15712 14912 15945 14940
rect 15712 14900 15718 14912
rect 15933 14909 15945 14912
rect 15979 14909 15991 14943
rect 15933 14903 15991 14909
rect 12032 14844 12572 14872
rect 12032 14832 12038 14844
rect 9398 14804 9404 14816
rect 9171 14776 9404 14804
rect 9171 14773 9183 14776
rect 9125 14767 9183 14773
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 1104 14714 22816 14736
rect 1104 14662 8982 14714
rect 9034 14662 9046 14714
rect 9098 14662 9110 14714
rect 9162 14662 9174 14714
rect 9226 14662 16982 14714
rect 17034 14662 17046 14714
rect 17098 14662 17110 14714
rect 17162 14662 17174 14714
rect 17226 14662 22816 14714
rect 1104 14640 22816 14662
rect 1578 14600 1584 14612
rect 1539 14572 1584 14600
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 8754 14560 8760 14612
rect 8812 14600 8818 14612
rect 9306 14600 9312 14612
rect 8812 14572 9312 14600
rect 8812 14560 8818 14572
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 10502 14560 10508 14612
rect 10560 14600 10566 14612
rect 12434 14600 12440 14612
rect 10560 14572 12440 14600
rect 10560 14560 10566 14572
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 13311 14603 13369 14609
rect 13311 14569 13323 14603
rect 13357 14600 13369 14603
rect 14366 14600 14372 14612
rect 13357 14572 14372 14600
rect 13357 14569 13369 14572
rect 13311 14563 13369 14569
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 1854 14532 1860 14544
rect 1815 14504 1860 14532
rect 1854 14492 1860 14504
rect 1912 14492 1918 14544
rect 1949 14535 2007 14541
rect 1949 14501 1961 14535
rect 1995 14532 2007 14535
rect 2038 14532 2044 14544
rect 1995 14504 2044 14532
rect 1995 14501 2007 14504
rect 1949 14495 2007 14501
rect 2038 14492 2044 14504
rect 2096 14492 2102 14544
rect 5626 14532 5632 14544
rect 5587 14504 5632 14532
rect 5626 14492 5632 14504
rect 5684 14492 5690 14544
rect 5810 14492 5816 14544
rect 5868 14532 5874 14544
rect 6549 14535 6607 14541
rect 6549 14532 6561 14535
rect 5868 14504 6561 14532
rect 5868 14492 5874 14504
rect 6549 14501 6561 14504
rect 6595 14501 6607 14535
rect 6549 14495 6607 14501
rect 6641 14535 6699 14541
rect 6641 14501 6653 14535
rect 6687 14532 6699 14535
rect 6822 14532 6828 14544
rect 6687 14504 6828 14532
rect 6687 14501 6699 14504
rect 6641 14495 6699 14501
rect 6822 14492 6828 14504
rect 6880 14492 6886 14544
rect 9398 14492 9404 14544
rect 9456 14532 9462 14544
rect 12158 14532 12164 14544
rect 9456 14504 11468 14532
rect 12119 14504 12164 14532
rect 9456 14492 9462 14504
rect 4430 14424 4436 14476
rect 4488 14464 4494 14476
rect 5169 14467 5227 14473
rect 5169 14464 5181 14467
rect 4488 14436 5181 14464
rect 4488 14424 4494 14436
rect 5169 14433 5181 14436
rect 5215 14433 5227 14467
rect 5169 14427 5227 14433
rect 5445 14467 5503 14473
rect 5445 14433 5457 14467
rect 5491 14464 5503 14467
rect 5718 14464 5724 14476
rect 5491 14436 5724 14464
rect 5491 14433 5503 14436
rect 5445 14427 5503 14433
rect 2501 14399 2559 14405
rect 2501 14365 2513 14399
rect 2547 14396 2559 14399
rect 2590 14396 2596 14408
rect 2547 14368 2596 14396
rect 2547 14365 2559 14368
rect 2501 14359 2559 14365
rect 2590 14356 2596 14368
rect 2648 14356 2654 14408
rect 5184 14396 5212 14427
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 10042 14464 10048 14476
rect 10003 14436 10048 14464
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 11440 14473 11468 14504
rect 12158 14492 12164 14504
rect 12216 14492 12222 14544
rect 15470 14532 15476 14544
rect 15431 14504 15476 14532
rect 15470 14492 15476 14504
rect 15528 14492 15534 14544
rect 11425 14467 11483 14473
rect 11425 14433 11437 14467
rect 11471 14464 11483 14467
rect 11790 14464 11796 14476
rect 11471 14436 11796 14464
rect 11471 14433 11483 14436
rect 11425 14427 11483 14433
rect 11790 14424 11796 14436
rect 11848 14424 11854 14476
rect 11974 14464 11980 14476
rect 11935 14436 11980 14464
rect 11974 14424 11980 14436
rect 12032 14424 12038 14476
rect 13240 14467 13298 14473
rect 13240 14433 13252 14467
rect 13286 14464 13298 14467
rect 13446 14464 13452 14476
rect 13286 14436 13452 14464
rect 13286 14433 13298 14436
rect 13240 14427 13298 14433
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 5350 14396 5356 14408
rect 5184 14368 5356 14396
rect 5350 14356 5356 14368
rect 5408 14396 5414 14408
rect 10502 14396 10508 14408
rect 5408 14368 10508 14396
rect 5408 14356 5414 14368
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 14185 14399 14243 14405
rect 14185 14365 14197 14399
rect 14231 14396 14243 14399
rect 14734 14396 14740 14408
rect 14231 14368 14740 14396
rect 14231 14365 14243 14368
rect 14185 14359 14243 14365
rect 14734 14356 14740 14368
rect 14792 14396 14798 14408
rect 15381 14399 15439 14405
rect 15381 14396 15393 14399
rect 14792 14368 15393 14396
rect 14792 14356 14798 14368
rect 15381 14365 15393 14368
rect 15427 14365 15439 14399
rect 15654 14396 15660 14408
rect 15615 14368 15660 14396
rect 15381 14359 15439 14365
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 7098 14328 7104 14340
rect 7011 14300 7104 14328
rect 7098 14288 7104 14300
rect 7156 14328 7162 14340
rect 7156 14300 7604 14328
rect 7156 14288 7162 14300
rect 3786 14260 3792 14272
rect 3747 14232 3792 14260
rect 3786 14220 3792 14232
rect 3844 14220 3850 14272
rect 7576 14269 7604 14300
rect 7561 14263 7619 14269
rect 7561 14229 7573 14263
rect 7607 14260 7619 14263
rect 8018 14260 8024 14272
rect 7607 14232 8024 14260
rect 7607 14229 7619 14232
rect 7561 14223 7619 14229
rect 8018 14220 8024 14232
rect 8076 14220 8082 14272
rect 9766 14220 9772 14272
rect 9824 14260 9830 14272
rect 9953 14263 10011 14269
rect 9953 14260 9965 14263
rect 9824 14232 9965 14260
rect 9824 14220 9830 14232
rect 9953 14229 9965 14232
rect 9999 14229 10011 14263
rect 14918 14260 14924 14272
rect 14879 14232 14924 14260
rect 9953 14223 10011 14229
rect 14918 14220 14924 14232
rect 14976 14220 14982 14272
rect 1104 14170 22816 14192
rect 1104 14118 4982 14170
rect 5034 14118 5046 14170
rect 5098 14118 5110 14170
rect 5162 14118 5174 14170
rect 5226 14118 12982 14170
rect 13034 14118 13046 14170
rect 13098 14118 13110 14170
rect 13162 14118 13174 14170
rect 13226 14118 20982 14170
rect 21034 14118 21046 14170
rect 21098 14118 21110 14170
rect 21162 14118 21174 14170
rect 21226 14118 22816 14170
rect 1104 14096 22816 14118
rect 1765 14059 1823 14065
rect 1765 14025 1777 14059
rect 1811 14056 1823 14059
rect 2038 14056 2044 14068
rect 1811 14028 2044 14056
rect 1811 14025 1823 14028
rect 1765 14019 1823 14025
rect 2038 14016 2044 14028
rect 2096 14016 2102 14068
rect 2130 14016 2136 14068
rect 2188 14056 2194 14068
rect 2869 14059 2927 14065
rect 2869 14056 2881 14059
rect 2188 14028 2881 14056
rect 2188 14016 2194 14028
rect 2869 14025 2881 14028
rect 2915 14025 2927 14059
rect 2869 14019 2927 14025
rect 5077 14059 5135 14065
rect 5077 14025 5089 14059
rect 5123 14056 5135 14059
rect 5350 14056 5356 14068
rect 5123 14028 5356 14056
rect 5123 14025 5135 14028
rect 5077 14019 5135 14025
rect 1854 13948 1860 14000
rect 1912 13988 1918 14000
rect 2884 13988 2912 14019
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 5810 14056 5816 14068
rect 5771 14028 5816 14056
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 10042 14056 10048 14068
rect 10003 14028 10048 14056
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 11790 14056 11796 14068
rect 11751 14028 11796 14056
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 14734 14056 14740 14068
rect 14695 14028 14740 14056
rect 14734 14016 14740 14028
rect 14792 14016 14798 14068
rect 15470 14016 15476 14068
rect 15528 14056 15534 14068
rect 15841 14059 15899 14065
rect 15841 14056 15853 14059
rect 15528 14028 15853 14056
rect 15528 14016 15534 14028
rect 15841 14025 15853 14028
rect 15887 14025 15899 14059
rect 15841 14019 15899 14025
rect 4709 13991 4767 13997
rect 4709 13988 4721 13991
rect 1912 13960 2820 13988
rect 2884 13960 4721 13988
rect 1912 13948 1918 13960
rect 1762 13880 1768 13932
rect 1820 13920 1826 13932
rect 1949 13923 2007 13929
rect 1949 13920 1961 13923
rect 1820 13892 1961 13920
rect 1820 13880 1826 13892
rect 1949 13889 1961 13892
rect 1995 13889 2007 13923
rect 2792 13920 2820 13960
rect 4709 13957 4721 13960
rect 4755 13957 4767 13991
rect 4709 13951 4767 13957
rect 14936 13960 16804 13988
rect 14936 13932 14964 13960
rect 3237 13923 3295 13929
rect 3237 13920 3249 13923
rect 2792 13892 3249 13920
rect 1949 13883 2007 13889
rect 3237 13889 3249 13892
rect 3283 13889 3295 13923
rect 3786 13920 3792 13932
rect 3747 13892 3792 13920
rect 3237 13883 3295 13889
rect 3786 13880 3792 13892
rect 3844 13880 3850 13932
rect 8846 13880 8852 13932
rect 8904 13920 8910 13932
rect 9125 13923 9183 13929
rect 9125 13920 9137 13923
rect 8904 13892 9137 13920
rect 8904 13880 8910 13892
rect 9125 13889 9137 13892
rect 9171 13889 9183 13923
rect 14918 13920 14924 13932
rect 14879 13892 14924 13920
rect 9125 13883 9183 13889
rect 14918 13880 14924 13892
rect 14976 13880 14982 13932
rect 15565 13923 15623 13929
rect 15565 13889 15577 13923
rect 15611 13920 15623 13923
rect 15654 13920 15660 13932
rect 15611 13892 15660 13920
rect 15611 13889 15623 13892
rect 15565 13883 15623 13889
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 16482 13920 16488 13932
rect 16443 13892 16488 13920
rect 16482 13880 16488 13892
rect 16540 13880 16546 13932
rect 16776 13929 16804 13960
rect 16761 13923 16819 13929
rect 16761 13889 16773 13923
rect 16807 13920 16819 13923
rect 17310 13920 17316 13932
rect 16807 13892 17316 13920
rect 16807 13889 16819 13892
rect 16761 13883 16819 13889
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 6181 13855 6239 13861
rect 6181 13821 6193 13855
rect 6227 13852 6239 13855
rect 6549 13855 6607 13861
rect 6549 13852 6561 13855
rect 6227 13824 6561 13852
rect 6227 13821 6239 13824
rect 6181 13815 6239 13821
rect 6549 13821 6561 13824
rect 6595 13852 6607 13855
rect 6822 13852 6828 13864
rect 6595 13824 6828 13852
rect 6595 13821 6607 13824
rect 6549 13815 6607 13821
rect 6822 13812 6828 13824
rect 6880 13852 6886 13864
rect 6917 13855 6975 13861
rect 6917 13852 6929 13855
rect 6880 13824 6929 13852
rect 6880 13812 6886 13824
rect 6917 13821 6929 13824
rect 6963 13821 6975 13855
rect 6917 13815 6975 13821
rect 2041 13787 2099 13793
rect 2041 13753 2053 13787
rect 2087 13784 2099 13787
rect 2130 13784 2136 13796
rect 2087 13756 2136 13784
rect 2087 13753 2099 13756
rect 2041 13747 2099 13753
rect 2130 13744 2136 13756
rect 2188 13744 2194 13796
rect 2590 13784 2596 13796
rect 2503 13756 2596 13784
rect 2590 13744 2596 13756
rect 2648 13784 2654 13796
rect 3142 13784 3148 13796
rect 2648 13756 3148 13784
rect 2648 13744 2654 13756
rect 3142 13744 3148 13756
rect 3200 13744 3206 13796
rect 4111 13787 4169 13793
rect 4111 13753 4123 13787
rect 4157 13753 4169 13787
rect 7558 13784 7564 13796
rect 7519 13756 7564 13784
rect 4111 13747 4169 13753
rect 2774 13676 2780 13728
rect 2832 13716 2838 13728
rect 3697 13719 3755 13725
rect 3697 13716 3709 13719
rect 2832 13688 3709 13716
rect 2832 13676 2838 13688
rect 3697 13685 3709 13688
rect 3743 13716 3755 13719
rect 4126 13716 4154 13747
rect 7558 13744 7564 13756
rect 7616 13744 7622 13796
rect 8941 13787 8999 13793
rect 8941 13753 8953 13787
rect 8987 13784 8999 13787
rect 9217 13787 9275 13793
rect 9217 13784 9229 13787
rect 8987 13756 9229 13784
rect 8987 13753 8999 13756
rect 8941 13747 8999 13753
rect 9217 13753 9229 13756
rect 9263 13784 9275 13787
rect 9306 13784 9312 13796
rect 9263 13756 9312 13784
rect 9263 13753 9275 13756
rect 9217 13747 9275 13753
rect 9306 13744 9312 13756
rect 9364 13744 9370 13796
rect 9769 13787 9827 13793
rect 9769 13753 9781 13787
rect 9815 13784 9827 13787
rect 9858 13784 9864 13796
rect 9815 13756 9864 13784
rect 9815 13753 9827 13756
rect 9769 13747 9827 13753
rect 9858 13744 9864 13756
rect 9916 13784 9922 13796
rect 12526 13784 12532 13796
rect 9916 13756 12532 13784
rect 9916 13744 9922 13756
rect 12526 13744 12532 13756
rect 12584 13744 12590 13796
rect 12621 13787 12679 13793
rect 12621 13753 12633 13787
rect 12667 13753 12679 13787
rect 12621 13747 12679 13753
rect 13173 13787 13231 13793
rect 13173 13753 13185 13787
rect 13219 13753 13231 13787
rect 15010 13784 15016 13796
rect 14971 13756 15016 13784
rect 13173 13747 13231 13753
rect 4430 13716 4436 13728
rect 3743 13688 4436 13716
rect 3743 13685 3755 13688
rect 3697 13679 3755 13685
rect 4430 13676 4436 13688
rect 4488 13676 4494 13728
rect 5445 13719 5503 13725
rect 5445 13685 5457 13719
rect 5491 13716 5503 13719
rect 5718 13716 5724 13728
rect 5491 13688 5724 13716
rect 5491 13685 5503 13688
rect 5445 13679 5503 13685
rect 5718 13676 5724 13688
rect 5776 13676 5782 13728
rect 11333 13719 11391 13725
rect 11333 13685 11345 13719
rect 11379 13716 11391 13719
rect 11606 13716 11612 13728
rect 11379 13688 11612 13716
rect 11379 13685 11391 13688
rect 11333 13679 11391 13685
rect 11606 13676 11612 13688
rect 11664 13676 11670 13728
rect 11698 13676 11704 13728
rect 11756 13716 11762 13728
rect 12158 13716 12164 13728
rect 11756 13688 12164 13716
rect 11756 13676 11762 13688
rect 12158 13676 12164 13688
rect 12216 13676 12222 13728
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12636 13716 12664 13747
rect 12492 13688 12664 13716
rect 13188 13716 13216 13747
rect 15010 13744 15016 13756
rect 15068 13744 15074 13796
rect 16301 13787 16359 13793
rect 16301 13753 16313 13787
rect 16347 13784 16359 13787
rect 16574 13784 16580 13796
rect 16347 13756 16580 13784
rect 16347 13753 16359 13756
rect 16301 13747 16359 13753
rect 16574 13744 16580 13756
rect 16632 13744 16638 13796
rect 13446 13716 13452 13728
rect 13188 13688 13452 13716
rect 12492 13676 12498 13688
rect 13446 13676 13452 13688
rect 13504 13676 13510 13728
rect 1104 13626 22816 13648
rect 1104 13574 8982 13626
rect 9034 13574 9046 13626
rect 9098 13574 9110 13626
rect 9162 13574 9174 13626
rect 9226 13574 16982 13626
rect 17034 13574 17046 13626
rect 17098 13574 17110 13626
rect 17162 13574 17174 13626
rect 17226 13574 22816 13626
rect 1104 13552 22816 13574
rect 1762 13472 1768 13524
rect 1820 13512 1826 13524
rect 2593 13515 2651 13521
rect 2593 13512 2605 13515
rect 1820 13484 2605 13512
rect 1820 13472 1826 13484
rect 2593 13481 2605 13484
rect 2639 13481 2651 13515
rect 2593 13475 2651 13481
rect 3786 13472 3792 13524
rect 3844 13512 3850 13524
rect 4157 13515 4215 13521
rect 4157 13512 4169 13515
rect 3844 13484 4169 13512
rect 3844 13472 3850 13484
rect 4157 13481 4169 13484
rect 4203 13481 4215 13515
rect 6270 13512 6276 13524
rect 6231 13484 6276 13512
rect 4157 13475 4215 13481
rect 6270 13472 6276 13484
rect 6328 13472 6334 13524
rect 6822 13512 6828 13524
rect 6783 13484 6828 13512
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 8846 13472 8852 13524
rect 8904 13512 8910 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 8904 13484 9045 13512
rect 8904 13472 8910 13484
rect 9033 13481 9045 13484
rect 9079 13481 9091 13515
rect 9033 13475 9091 13481
rect 11514 13472 11520 13524
rect 11572 13512 11578 13524
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 11572 13484 11621 13512
rect 11572 13472 11578 13484
rect 11609 13481 11621 13484
rect 11655 13481 11667 13515
rect 11609 13475 11667 13481
rect 12526 13472 12532 13524
rect 12584 13512 12590 13524
rect 12805 13515 12863 13521
rect 12805 13512 12817 13515
rect 12584 13484 12817 13512
rect 12584 13472 12590 13484
rect 12805 13481 12817 13484
rect 12851 13481 12863 13515
rect 12805 13475 12863 13481
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 15565 13515 15623 13521
rect 15565 13512 15577 13515
rect 15528 13484 15577 13512
rect 15528 13472 15534 13484
rect 15565 13481 15577 13484
rect 15611 13481 15623 13515
rect 16482 13512 16488 13524
rect 16443 13484 16488 13512
rect 15565 13475 15623 13481
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 7558 13404 7564 13456
rect 7616 13444 7622 13456
rect 7837 13447 7895 13453
rect 7837 13444 7849 13447
rect 7616 13416 7849 13444
rect 7616 13404 7622 13416
rect 7837 13413 7849 13416
rect 7883 13413 7895 13447
rect 7837 13407 7895 13413
rect 9766 13404 9772 13456
rect 9824 13444 9830 13456
rect 9861 13447 9919 13453
rect 9861 13444 9873 13447
rect 9824 13416 9873 13444
rect 9824 13404 9830 13416
rect 9861 13413 9873 13416
rect 9907 13444 9919 13447
rect 10226 13444 10232 13456
rect 9907 13416 10232 13444
rect 9907 13413 9919 13416
rect 9861 13407 9919 13413
rect 10226 13404 10232 13416
rect 10284 13404 10290 13456
rect 13173 13447 13231 13453
rect 13173 13413 13185 13447
rect 13219 13444 13231 13447
rect 13262 13444 13268 13456
rect 13219 13416 13268 13444
rect 13219 13413 13231 13416
rect 13173 13407 13231 13413
rect 13262 13404 13268 13416
rect 13320 13404 13326 13456
rect 17034 13444 17040 13456
rect 16995 13416 17040 13444
rect 17034 13404 17040 13416
rect 17092 13404 17098 13456
rect 1762 13376 1768 13388
rect 1723 13348 1768 13376
rect 1762 13336 1768 13348
rect 1820 13336 1826 13388
rect 4062 13376 4068 13388
rect 4023 13348 4068 13376
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 4246 13336 4252 13388
rect 4304 13376 4310 13388
rect 4525 13379 4583 13385
rect 4525 13376 4537 13379
rect 4304 13348 4537 13376
rect 4304 13336 4310 13348
rect 4525 13345 4537 13348
rect 4571 13345 4583 13379
rect 4525 13339 4583 13345
rect 14921 13379 14979 13385
rect 14921 13345 14933 13379
rect 14967 13376 14979 13379
rect 15010 13376 15016 13388
rect 14967 13348 15016 13376
rect 14967 13345 14979 13348
rect 14921 13339 14979 13345
rect 15010 13336 15016 13348
rect 15068 13376 15074 13388
rect 15470 13376 15476 13388
rect 15068 13348 15476 13376
rect 15068 13336 15074 13348
rect 15470 13336 15476 13348
rect 15528 13336 15534 13388
rect 20968 13379 21026 13385
rect 20968 13345 20980 13379
rect 21014 13376 21026 13379
rect 21450 13376 21456 13388
rect 21014 13348 21456 13376
rect 21014 13345 21026 13348
rect 20968 13339 21026 13345
rect 21450 13336 21456 13348
rect 21508 13336 21514 13388
rect 5902 13308 5908 13320
rect 5863 13280 5908 13308
rect 5902 13268 5908 13280
rect 5960 13268 5966 13320
rect 7745 13311 7803 13317
rect 7745 13277 7757 13311
rect 7791 13277 7803 13311
rect 8018 13308 8024 13320
rect 7979 13280 8024 13308
rect 7745 13271 7803 13277
rect 7760 13240 7788 13271
rect 8018 13268 8024 13280
rect 8076 13268 8082 13320
rect 9766 13308 9772 13320
rect 9727 13280 9772 13308
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 9858 13268 9864 13320
rect 9916 13308 9922 13320
rect 10045 13311 10103 13317
rect 10045 13308 10057 13311
rect 9916 13280 10057 13308
rect 9916 13268 9922 13280
rect 10045 13277 10057 13280
rect 10091 13277 10103 13311
rect 10045 13271 10103 13277
rect 11241 13311 11299 13317
rect 11241 13277 11253 13311
rect 11287 13308 11299 13311
rect 11330 13308 11336 13320
rect 11287 13280 11336 13308
rect 11287 13277 11299 13280
rect 11241 13271 11299 13277
rect 11330 13268 11336 13280
rect 11388 13268 11394 13320
rect 11606 13268 11612 13320
rect 11664 13308 11670 13320
rect 12802 13308 12808 13320
rect 11664 13280 12808 13308
rect 11664 13268 11670 13280
rect 12802 13268 12808 13280
rect 12860 13308 12866 13320
rect 13081 13311 13139 13317
rect 13081 13308 13093 13311
rect 12860 13280 13093 13308
rect 12860 13268 12866 13280
rect 13081 13277 13093 13280
rect 13127 13277 13139 13311
rect 13446 13308 13452 13320
rect 13407 13280 13452 13308
rect 13081 13271 13139 13277
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 16945 13311 17003 13317
rect 16945 13277 16957 13311
rect 16991 13277 17003 13311
rect 17310 13308 17316 13320
rect 17271 13280 17316 13308
rect 16945 13271 17003 13277
rect 8110 13240 8116 13252
rect 7760 13212 8116 13240
rect 8110 13200 8116 13212
rect 8168 13200 8174 13252
rect 16850 13200 16856 13252
rect 16908 13240 16914 13252
rect 16960 13240 16988 13271
rect 17310 13268 17316 13280
rect 17368 13268 17374 13320
rect 16908 13212 16988 13240
rect 16908 13200 16914 13212
rect 1854 13172 1860 13184
rect 1815 13144 1860 13172
rect 1854 13132 1860 13144
rect 1912 13132 1918 13184
rect 2958 13172 2964 13184
rect 2919 13144 2964 13172
rect 2958 13132 2964 13144
rect 3016 13132 3022 13184
rect 3694 13172 3700 13184
rect 3655 13144 3700 13172
rect 3694 13132 3700 13144
rect 3752 13132 3758 13184
rect 5261 13175 5319 13181
rect 5261 13141 5273 13175
rect 5307 13172 5319 13175
rect 5718 13172 5724 13184
rect 5307 13144 5724 13172
rect 5307 13141 5319 13144
rect 5261 13135 5319 13141
rect 5718 13132 5724 13144
rect 5776 13132 5782 13184
rect 6730 13132 6736 13184
rect 6788 13172 6794 13184
rect 7101 13175 7159 13181
rect 7101 13172 7113 13175
rect 6788 13144 7113 13172
rect 6788 13132 6794 13144
rect 7101 13141 7113 13144
rect 7147 13141 7159 13175
rect 7101 13135 7159 13141
rect 10134 13132 10140 13184
rect 10192 13172 10198 13184
rect 10781 13175 10839 13181
rect 10781 13172 10793 13175
rect 10192 13144 10793 13172
rect 10192 13132 10198 13144
rect 10781 13141 10793 13144
rect 10827 13172 10839 13175
rect 11238 13172 11244 13184
rect 10827 13144 11244 13172
rect 10827 13141 10839 13144
rect 10781 13135 10839 13141
rect 11238 13132 11244 13144
rect 11296 13132 11302 13184
rect 12161 13175 12219 13181
rect 12161 13141 12173 13175
rect 12207 13172 12219 13175
rect 12434 13172 12440 13184
rect 12207 13144 12440 13172
rect 12207 13141 12219 13144
rect 12161 13135 12219 13141
rect 12434 13132 12440 13144
rect 12492 13132 12498 13184
rect 14274 13172 14280 13184
rect 14235 13144 14280 13172
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 20806 13132 20812 13184
rect 20864 13172 20870 13184
rect 21039 13175 21097 13181
rect 21039 13172 21051 13175
rect 20864 13144 21051 13172
rect 20864 13132 20870 13144
rect 21039 13141 21051 13144
rect 21085 13141 21097 13175
rect 21039 13135 21097 13141
rect 1104 13082 22816 13104
rect 1104 13030 4982 13082
rect 5034 13030 5046 13082
rect 5098 13030 5110 13082
rect 5162 13030 5174 13082
rect 5226 13030 12982 13082
rect 13034 13030 13046 13082
rect 13098 13030 13110 13082
rect 13162 13030 13174 13082
rect 13226 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 22816 13082
rect 1104 13008 22816 13030
rect 2682 12928 2688 12980
rect 2740 12968 2746 12980
rect 3421 12971 3479 12977
rect 3421 12968 3433 12971
rect 2740 12940 3433 12968
rect 2740 12928 2746 12940
rect 3421 12937 3433 12940
rect 3467 12968 3479 12971
rect 4062 12968 4068 12980
rect 3467 12940 4068 12968
rect 3467 12937 3479 12940
rect 3421 12931 3479 12937
rect 1762 12860 1768 12912
rect 1820 12900 1826 12912
rect 3050 12900 3056 12912
rect 1820 12872 3056 12900
rect 1820 12860 1826 12872
rect 3050 12860 3056 12872
rect 3108 12860 3114 12912
rect 1670 12832 1676 12844
rect 1583 12804 1676 12832
rect 1670 12792 1676 12804
rect 1728 12832 1734 12844
rect 2958 12832 2964 12844
rect 1728 12804 2964 12832
rect 1728 12792 1734 12804
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 3436 12764 3464 12931
rect 4062 12928 4068 12940
rect 4120 12968 4126 12980
rect 4525 12971 4583 12977
rect 4525 12968 4537 12971
rect 4120 12940 4537 12968
rect 4120 12928 4126 12940
rect 4525 12937 4537 12940
rect 4571 12937 4583 12971
rect 4525 12931 4583 12937
rect 7558 12928 7564 12980
rect 7616 12968 7622 12980
rect 7653 12971 7711 12977
rect 7653 12968 7665 12971
rect 7616 12940 7665 12968
rect 7616 12928 7622 12940
rect 7653 12937 7665 12940
rect 7699 12937 7711 12971
rect 7653 12931 7711 12937
rect 9306 12928 9312 12980
rect 9364 12968 9370 12980
rect 9953 12971 10011 12977
rect 9953 12968 9965 12971
rect 9364 12940 9965 12968
rect 9364 12928 9370 12940
rect 9953 12937 9965 12940
rect 9999 12968 10011 12971
rect 10042 12968 10048 12980
rect 9999 12940 10048 12968
rect 9999 12937 10011 12940
rect 9953 12931 10011 12937
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 10226 12968 10232 12980
rect 10187 12940 10232 12968
rect 10226 12928 10232 12940
rect 10284 12928 10290 12980
rect 15197 12971 15255 12977
rect 15197 12937 15209 12971
rect 15243 12968 15255 12971
rect 15470 12968 15476 12980
rect 15243 12940 15476 12968
rect 15243 12937 15255 12940
rect 15197 12931 15255 12937
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 16574 12928 16580 12980
rect 16632 12968 16638 12980
rect 16669 12971 16727 12977
rect 16669 12968 16681 12971
rect 16632 12940 16681 12968
rect 16632 12928 16638 12940
rect 16669 12937 16681 12940
rect 16715 12937 16727 12971
rect 21450 12968 21456 12980
rect 21411 12940 21456 12968
rect 16669 12931 16727 12937
rect 21450 12928 21456 12940
rect 21508 12928 21514 12980
rect 4430 12860 4436 12912
rect 4488 12900 4494 12912
rect 6181 12903 6239 12909
rect 6181 12900 6193 12903
rect 4488 12872 6193 12900
rect 4488 12860 4494 12872
rect 6181 12869 6193 12872
rect 6227 12900 6239 12903
rect 6270 12900 6276 12912
rect 6227 12872 6276 12900
rect 6227 12869 6239 12872
rect 6181 12863 6239 12869
rect 6270 12860 6276 12872
rect 6328 12860 6334 12912
rect 6362 12860 6368 12912
rect 6420 12900 6426 12912
rect 6641 12903 6699 12909
rect 6641 12900 6653 12903
rect 6420 12872 6653 12900
rect 6420 12860 6426 12872
rect 6641 12869 6653 12872
rect 6687 12900 6699 12903
rect 11422 12900 11428 12912
rect 6687 12872 11428 12900
rect 6687 12869 6699 12872
rect 6641 12863 6699 12869
rect 11422 12860 11428 12872
rect 11480 12860 11486 12912
rect 5902 12832 5908 12844
rect 5815 12804 5908 12832
rect 5902 12792 5908 12804
rect 5960 12832 5966 12844
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 5960 12804 7297 12832
rect 5960 12792 5966 12804
rect 7285 12801 7297 12804
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12832 9091 12835
rect 9306 12832 9312 12844
rect 9079 12804 9312 12832
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 11330 12832 11336 12844
rect 11291 12804 11336 12832
rect 11330 12792 11336 12804
rect 11388 12792 11394 12844
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12832 13231 12835
rect 13262 12832 13268 12844
rect 13219 12804 13268 12832
rect 13219 12801 13231 12804
rect 13173 12795 13231 12801
rect 13262 12792 13268 12804
rect 13320 12832 13326 12844
rect 13449 12835 13507 12841
rect 13449 12832 13461 12835
rect 13320 12804 13461 12832
rect 13320 12792 13326 12804
rect 13449 12801 13461 12804
rect 13495 12801 13507 12835
rect 14274 12832 14280 12844
rect 14235 12804 14280 12832
rect 13449 12795 13507 12801
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 20438 12832 20444 12844
rect 20399 12804 20444 12832
rect 20438 12792 20444 12804
rect 20496 12792 20502 12844
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 3436 12736 3617 12764
rect 3605 12733 3617 12736
rect 3651 12733 3663 12767
rect 3605 12727 3663 12733
rect 3694 12724 3700 12776
rect 3752 12764 3758 12776
rect 4157 12767 4215 12773
rect 4157 12764 4169 12767
rect 3752 12736 4169 12764
rect 3752 12724 3758 12736
rect 4157 12733 4169 12736
rect 4203 12764 4215 12767
rect 4522 12764 4528 12776
rect 4203 12736 4528 12764
rect 4203 12733 4215 12736
rect 4157 12727 4215 12733
rect 4522 12724 4528 12736
rect 4580 12764 4586 12776
rect 5074 12764 5080 12776
rect 4580 12736 5080 12764
rect 4580 12724 4586 12736
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 5442 12764 5448 12776
rect 5403 12736 5448 12764
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 5718 12764 5724 12776
rect 5631 12736 5724 12764
rect 5718 12724 5724 12736
rect 5776 12764 5782 12776
rect 6546 12764 6552 12776
rect 5776 12736 6552 12764
rect 5776 12724 5782 12736
rect 6546 12724 6552 12736
rect 6604 12724 6610 12776
rect 6730 12724 6736 12776
rect 6788 12764 6794 12776
rect 6860 12767 6918 12773
rect 6860 12764 6872 12767
rect 6788 12736 6872 12764
rect 6788 12724 6794 12736
rect 6860 12733 6872 12736
rect 6906 12733 6918 12767
rect 6860 12727 6918 12733
rect 10502 12724 10508 12776
rect 10560 12764 10566 12776
rect 10781 12767 10839 12773
rect 10781 12764 10793 12767
rect 10560 12736 10793 12764
rect 10560 12724 10566 12736
rect 10781 12733 10793 12736
rect 10827 12733 10839 12767
rect 11238 12764 11244 12776
rect 11199 12736 11244 12764
rect 10781 12727 10839 12733
rect 11238 12724 11244 12736
rect 11296 12724 11302 12776
rect 12253 12767 12311 12773
rect 12253 12733 12265 12767
rect 12299 12764 12311 12767
rect 12434 12764 12440 12776
rect 12299 12736 12440 12764
rect 12299 12733 12311 12736
rect 12253 12727 12311 12733
rect 12434 12724 12440 12736
rect 12492 12764 12498 12776
rect 12529 12767 12587 12773
rect 12529 12764 12541 12767
rect 12492 12736 12541 12764
rect 12492 12724 12498 12736
rect 12529 12733 12541 12736
rect 12575 12733 12587 12767
rect 12529 12727 12587 12733
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 16574 12764 16580 12776
rect 16347 12736 16580 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 16574 12724 16580 12736
rect 16632 12764 16638 12776
rect 17034 12764 17040 12776
rect 16632 12736 17040 12764
rect 16632 12724 16638 12736
rect 17034 12724 17040 12736
rect 17092 12764 17098 12776
rect 17405 12767 17463 12773
rect 17405 12764 17417 12767
rect 17092 12736 17417 12764
rect 17092 12724 17098 12736
rect 17405 12733 17417 12736
rect 17451 12733 17463 12767
rect 17405 12727 17463 12733
rect 1765 12699 1823 12705
rect 1765 12665 1777 12699
rect 1811 12696 1823 12699
rect 1854 12696 1860 12708
rect 1811 12668 1860 12696
rect 1811 12665 1823 12668
rect 1765 12659 1823 12665
rect 1854 12656 1860 12668
rect 1912 12656 1918 12708
rect 2038 12656 2044 12708
rect 2096 12696 2102 12708
rect 2317 12699 2375 12705
rect 2317 12696 2329 12699
rect 2096 12668 2329 12696
rect 2096 12656 2102 12668
rect 2317 12665 2329 12668
rect 2363 12665 2375 12699
rect 2317 12659 2375 12665
rect 6270 12656 6276 12708
rect 6328 12696 6334 12708
rect 8849 12699 8907 12705
rect 8849 12696 8861 12699
rect 6328 12668 8861 12696
rect 6328 12656 6334 12668
rect 8849 12665 8861 12668
rect 8895 12696 8907 12699
rect 9354 12699 9412 12705
rect 9354 12696 9366 12699
rect 8895 12668 9366 12696
rect 8895 12665 8907 12668
rect 8849 12659 8907 12665
rect 9354 12665 9366 12668
rect 9400 12696 9412 12699
rect 11514 12696 11520 12708
rect 9400 12668 11520 12696
rect 9400 12665 9412 12668
rect 9354 12659 9412 12665
rect 11514 12656 11520 12668
rect 11572 12696 11578 12708
rect 11793 12699 11851 12705
rect 11793 12696 11805 12699
rect 11572 12668 11805 12696
rect 11572 12656 11578 12668
rect 11793 12665 11805 12668
rect 11839 12696 11851 12699
rect 13446 12696 13452 12708
rect 11839 12668 13452 12696
rect 11839 12665 11851 12668
rect 11793 12659 11851 12665
rect 13446 12656 13452 12668
rect 13504 12696 13510 12708
rect 14185 12699 14243 12705
rect 14185 12696 14197 12699
rect 13504 12668 14197 12696
rect 13504 12656 13510 12668
rect 14185 12665 14197 12668
rect 14231 12696 14243 12699
rect 14639 12699 14697 12705
rect 14639 12696 14651 12699
rect 14231 12668 14651 12696
rect 14231 12665 14243 12668
rect 14185 12659 14243 12665
rect 14639 12665 14651 12668
rect 14685 12696 14697 12699
rect 16206 12696 16212 12708
rect 14685 12668 16212 12696
rect 14685 12665 14697 12668
rect 14639 12659 14697 12665
rect 16206 12656 16212 12668
rect 16264 12656 16270 12708
rect 20533 12699 20591 12705
rect 20533 12665 20545 12699
rect 20579 12665 20591 12699
rect 21082 12696 21088 12708
rect 21043 12668 21088 12696
rect 20533 12659 20591 12665
rect 1872 12628 1900 12656
rect 2593 12631 2651 12637
rect 2593 12628 2605 12631
rect 1872 12600 2605 12628
rect 2593 12597 2605 12600
rect 2639 12597 2651 12631
rect 2593 12591 2651 12597
rect 3881 12631 3939 12637
rect 3881 12597 3893 12631
rect 3927 12628 3939 12631
rect 4062 12628 4068 12640
rect 3927 12600 4068 12628
rect 3927 12597 3939 12600
rect 3881 12591 3939 12597
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 4525 12631 4583 12637
rect 4525 12597 4537 12631
rect 4571 12628 4583 12631
rect 4709 12631 4767 12637
rect 4709 12628 4721 12631
rect 4571 12600 4721 12628
rect 4571 12597 4583 12600
rect 4525 12591 4583 12597
rect 4709 12597 4721 12600
rect 4755 12628 4767 12631
rect 5077 12631 5135 12637
rect 5077 12628 5089 12631
rect 4755 12600 5089 12628
rect 4755 12597 4767 12600
rect 4709 12591 4767 12597
rect 5077 12597 5089 12600
rect 5123 12628 5135 12631
rect 5442 12628 5448 12640
rect 5123 12600 5448 12628
rect 5123 12597 5135 12600
rect 5077 12591 5135 12597
rect 5442 12588 5448 12600
rect 5500 12628 5506 12640
rect 6454 12628 6460 12640
rect 5500 12600 6460 12628
rect 5500 12588 5506 12600
rect 6454 12588 6460 12600
rect 6512 12588 6518 12640
rect 6638 12588 6644 12640
rect 6696 12628 6702 12640
rect 6963 12631 7021 12637
rect 6963 12628 6975 12631
rect 6696 12600 6975 12628
rect 6696 12588 6702 12600
rect 6963 12597 6975 12600
rect 7009 12597 7021 12631
rect 8110 12628 8116 12640
rect 8071 12600 8116 12628
rect 6963 12591 7021 12597
rect 8110 12588 8116 12600
rect 8168 12588 8174 12640
rect 10502 12588 10508 12640
rect 10560 12628 10566 12640
rect 10597 12631 10655 12637
rect 10597 12628 10609 12631
rect 10560 12600 10609 12628
rect 10560 12588 10566 12600
rect 10597 12597 10609 12600
rect 10643 12597 10655 12631
rect 20162 12628 20168 12640
rect 20123 12600 20168 12628
rect 10597 12591 10655 12597
rect 20162 12588 20168 12600
rect 20220 12628 20226 12640
rect 20548 12628 20576 12659
rect 21082 12656 21088 12668
rect 21140 12656 21146 12708
rect 20220 12600 20576 12628
rect 20220 12588 20226 12600
rect 1104 12538 22816 12560
rect 1104 12486 8982 12538
rect 9034 12486 9046 12538
rect 9098 12486 9110 12538
rect 9162 12486 9174 12538
rect 9226 12486 16982 12538
rect 17034 12486 17046 12538
rect 17098 12486 17110 12538
rect 17162 12486 17174 12538
rect 17226 12486 22816 12538
rect 1104 12464 22816 12486
rect 3050 12384 3056 12436
rect 3108 12424 3114 12436
rect 4985 12427 5043 12433
rect 4985 12424 4997 12427
rect 3108 12396 4997 12424
rect 3108 12384 3114 12396
rect 4985 12393 4997 12396
rect 5031 12393 5043 12427
rect 4985 12387 5043 12393
rect 5074 12384 5080 12436
rect 5132 12424 5138 12436
rect 6457 12427 6515 12433
rect 6457 12424 6469 12427
rect 5132 12396 6469 12424
rect 5132 12384 5138 12396
rect 6457 12393 6469 12396
rect 6503 12393 6515 12427
rect 6457 12387 6515 12393
rect 9125 12427 9183 12433
rect 9125 12393 9137 12427
rect 9171 12424 9183 12427
rect 9306 12424 9312 12436
rect 9171 12396 9312 12424
rect 9171 12393 9183 12396
rect 9125 12387 9183 12393
rect 9306 12384 9312 12396
rect 9364 12424 9370 12436
rect 9769 12427 9827 12433
rect 9769 12424 9781 12427
rect 9364 12396 9781 12424
rect 9364 12384 9370 12396
rect 9769 12393 9781 12396
rect 9815 12393 9827 12427
rect 9769 12387 9827 12393
rect 11149 12427 11207 12433
rect 11149 12393 11161 12427
rect 11195 12424 11207 12427
rect 11330 12424 11336 12436
rect 11195 12396 11336 12424
rect 11195 12393 11207 12396
rect 11149 12387 11207 12393
rect 11330 12384 11336 12396
rect 11388 12384 11394 12436
rect 12802 12384 12808 12436
rect 12860 12424 12866 12436
rect 12989 12427 13047 12433
rect 12989 12424 13001 12427
rect 12860 12396 13001 12424
rect 12860 12384 12866 12396
rect 12989 12393 13001 12396
rect 13035 12393 13047 12427
rect 16574 12424 16580 12436
rect 16535 12396 16580 12424
rect 12989 12387 13047 12393
rect 16574 12384 16580 12396
rect 16632 12384 16638 12436
rect 20438 12424 20444 12436
rect 20399 12396 20444 12424
rect 20438 12384 20444 12396
rect 20496 12384 20502 12436
rect 20548 12396 21128 12424
rect 1762 12356 1768 12368
rect 1723 12328 1768 12356
rect 1762 12316 1768 12328
rect 1820 12316 1826 12368
rect 3881 12359 3939 12365
rect 3881 12325 3893 12359
rect 3927 12356 3939 12359
rect 4246 12356 4252 12368
rect 3927 12328 4252 12356
rect 3927 12325 3939 12328
rect 3881 12319 3939 12325
rect 4246 12316 4252 12328
rect 4304 12316 4310 12368
rect 4430 12365 4436 12368
rect 4427 12356 4436 12365
rect 4391 12328 4436 12356
rect 4427 12319 4436 12328
rect 4430 12316 4436 12319
rect 4488 12316 4494 12368
rect 11241 12359 11299 12365
rect 11241 12325 11253 12359
rect 11287 12356 11299 12359
rect 11514 12356 11520 12368
rect 11287 12328 11520 12356
rect 11287 12325 11299 12328
rect 11241 12319 11299 12325
rect 11514 12316 11520 12328
rect 11572 12316 11578 12368
rect 14274 12316 14280 12368
rect 14332 12356 14338 12368
rect 14369 12359 14427 12365
rect 14369 12356 14381 12359
rect 14332 12328 14381 12356
rect 14332 12316 14338 12328
rect 14369 12325 14381 12328
rect 14415 12325 14427 12359
rect 14369 12319 14427 12325
rect 16019 12359 16077 12365
rect 16019 12325 16031 12359
rect 16065 12356 16077 12359
rect 16206 12356 16212 12368
rect 16065 12328 16212 12356
rect 16065 12325 16077 12328
rect 16019 12319 16077 12325
rect 16206 12316 16212 12328
rect 16264 12316 16270 12368
rect 19981 12359 20039 12365
rect 19981 12325 19993 12359
rect 20027 12356 20039 12359
rect 20162 12356 20168 12368
rect 20027 12328 20168 12356
rect 20027 12325 20039 12328
rect 19981 12319 20039 12325
rect 20162 12316 20168 12328
rect 20220 12316 20226 12368
rect 4062 12288 4068 12300
rect 4023 12260 4068 12288
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 5813 12291 5871 12297
rect 5813 12288 5825 12291
rect 5592 12260 5825 12288
rect 5592 12248 5598 12260
rect 5813 12257 5825 12260
rect 5859 12288 5871 12291
rect 7374 12288 7380 12300
rect 5859 12260 6960 12288
rect 7335 12260 7380 12288
rect 5859 12257 5871 12260
rect 5813 12251 5871 12257
rect 1670 12220 1676 12232
rect 1631 12192 1676 12220
rect 1670 12180 1676 12192
rect 1728 12180 1734 12232
rect 2038 12220 2044 12232
rect 1999 12192 2044 12220
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 6181 12223 6239 12229
rect 5684 12192 5994 12220
rect 5684 12180 5690 12192
rect 5966 12161 5994 12192
rect 6181 12189 6193 12223
rect 6227 12220 6239 12223
rect 6270 12220 6276 12232
rect 6227 12192 6276 12220
rect 6227 12189 6239 12192
rect 6181 12183 6239 12189
rect 6270 12180 6276 12192
rect 6328 12180 6334 12232
rect 5966 12155 6036 12161
rect 5966 12124 5990 12155
rect 5978 12121 5990 12124
rect 6024 12152 6036 12155
rect 6362 12152 6368 12164
rect 6024 12124 6368 12152
rect 6024 12121 6036 12124
rect 5978 12115 6036 12121
rect 6362 12112 6368 12124
rect 6420 12112 6426 12164
rect 6932 12161 6960 12260
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 9674 12288 9680 12300
rect 9635 12260 9680 12288
rect 9674 12248 9680 12260
rect 9732 12248 9738 12300
rect 10042 12248 10048 12300
rect 10100 12288 10106 12300
rect 11422 12297 11428 12300
rect 10137 12291 10195 12297
rect 10137 12288 10149 12291
rect 10100 12260 10149 12288
rect 10100 12248 10106 12260
rect 10137 12257 10149 12260
rect 10183 12257 10195 12291
rect 11388 12291 11428 12297
rect 11388 12288 11400 12291
rect 11335 12260 11400 12288
rect 10137 12251 10195 12257
rect 11388 12257 11400 12260
rect 11480 12288 11486 12300
rect 12710 12288 12716 12300
rect 11480 12260 12716 12288
rect 11388 12251 11428 12257
rect 11422 12248 11428 12251
rect 11480 12248 11486 12260
rect 12710 12248 12716 12260
rect 12768 12248 12774 12300
rect 13354 12248 13360 12300
rect 13412 12288 13418 12300
rect 13633 12291 13691 12297
rect 13633 12288 13645 12291
rect 13412 12260 13645 12288
rect 13412 12248 13418 12260
rect 13633 12257 13645 12260
rect 13679 12257 13691 12291
rect 14182 12288 14188 12300
rect 14143 12260 14188 12288
rect 13633 12251 13691 12257
rect 14182 12248 14188 12260
rect 14240 12248 14246 12300
rect 19610 12248 19616 12300
rect 19668 12288 19674 12300
rect 19889 12291 19947 12297
rect 19889 12288 19901 12291
rect 19668 12260 19901 12288
rect 19668 12248 19674 12260
rect 19889 12257 19901 12260
rect 19935 12288 19947 12291
rect 20548 12288 20576 12396
rect 20806 12316 20812 12368
rect 20864 12356 20870 12368
rect 21100 12365 21128 12396
rect 20993 12359 21051 12365
rect 20993 12356 21005 12359
rect 20864 12328 21005 12356
rect 20864 12316 20870 12328
rect 20993 12325 21005 12328
rect 21039 12325 21051 12359
rect 20993 12319 21051 12325
rect 21085 12359 21143 12365
rect 21085 12325 21097 12359
rect 21131 12356 21143 12359
rect 21726 12356 21732 12368
rect 21131 12328 21732 12356
rect 21131 12325 21143 12328
rect 21085 12319 21143 12325
rect 21726 12316 21732 12328
rect 21784 12316 21790 12368
rect 19935 12260 20576 12288
rect 19935 12257 19947 12260
rect 19889 12251 19947 12257
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 11609 12223 11667 12229
rect 11609 12220 11621 12223
rect 11020 12192 11621 12220
rect 11020 12180 11026 12192
rect 11609 12189 11621 12192
rect 11655 12189 11667 12223
rect 15654 12220 15660 12232
rect 15615 12192 15660 12220
rect 11609 12183 11667 12189
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 15746 12180 15752 12232
rect 15804 12220 15810 12232
rect 21082 12220 21088 12232
rect 15804 12192 21088 12220
rect 15804 12180 15810 12192
rect 21082 12180 21088 12192
rect 21140 12220 21146 12232
rect 21269 12223 21327 12229
rect 21269 12220 21281 12223
rect 21140 12192 21281 12220
rect 21140 12180 21146 12192
rect 21269 12189 21281 12192
rect 21315 12189 21327 12223
rect 21269 12183 21327 12189
rect 6917 12155 6975 12161
rect 6917 12121 6929 12155
rect 6963 12152 6975 12155
rect 6963 12124 10732 12152
rect 6963 12121 6975 12124
rect 6917 12115 6975 12121
rect 10704 12096 10732 12124
rect 11238 12112 11244 12164
rect 11296 12152 11302 12164
rect 11517 12155 11575 12161
rect 11517 12152 11529 12155
rect 11296 12124 11529 12152
rect 11296 12112 11302 12124
rect 11517 12121 11529 12124
rect 11563 12121 11575 12155
rect 11517 12115 11575 12121
rect 2774 12084 2780 12096
rect 2735 12056 2780 12084
rect 2774 12044 2780 12056
rect 2832 12044 2838 12096
rect 5350 12084 5356 12096
rect 5311 12056 5356 12084
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 5718 12084 5724 12096
rect 5679 12056 5724 12084
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 6086 12084 6092 12096
rect 6047 12056 6092 12084
rect 6086 12044 6092 12056
rect 6144 12044 6150 12096
rect 7282 12084 7288 12096
rect 7243 12056 7288 12084
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 7515 12087 7573 12093
rect 7515 12053 7527 12087
rect 7561 12084 7573 12087
rect 7650 12084 7656 12096
rect 7561 12056 7656 12084
rect 7561 12053 7573 12056
rect 7515 12047 7573 12053
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 8478 12044 8484 12096
rect 8536 12084 8542 12096
rect 9401 12087 9459 12093
rect 9401 12084 9413 12087
rect 8536 12056 9413 12084
rect 8536 12044 8542 12056
rect 9401 12053 9413 12056
rect 9447 12084 9459 12087
rect 9766 12084 9772 12096
rect 9447 12056 9772 12084
rect 9447 12053 9459 12056
rect 9401 12047 9459 12053
rect 9766 12044 9772 12056
rect 9824 12044 9830 12096
rect 10686 12084 10692 12096
rect 10647 12056 10692 12084
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 11882 12084 11888 12096
rect 11843 12056 11888 12084
rect 11882 12044 11888 12056
rect 11940 12044 11946 12096
rect 16942 12084 16948 12096
rect 16903 12056 16948 12084
rect 16942 12044 16948 12056
rect 17000 12044 17006 12096
rect 18322 12084 18328 12096
rect 18283 12056 18328 12084
rect 18322 12044 18328 12056
rect 18380 12044 18386 12096
rect 1104 11994 22816 12016
rect 1104 11942 4982 11994
rect 5034 11942 5046 11994
rect 5098 11942 5110 11994
rect 5162 11942 5174 11994
rect 5226 11942 12982 11994
rect 13034 11942 13046 11994
rect 13098 11942 13110 11994
rect 13162 11942 13174 11994
rect 13226 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 22816 11994
rect 1104 11920 22816 11942
rect 4614 11840 4620 11892
rect 4672 11880 4678 11892
rect 5629 11883 5687 11889
rect 5629 11880 5641 11883
rect 4672 11852 5641 11880
rect 4672 11840 4678 11852
rect 5629 11849 5641 11852
rect 5675 11849 5687 11883
rect 5629 11843 5687 11849
rect 8113 11883 8171 11889
rect 8113 11849 8125 11883
rect 8159 11880 8171 11883
rect 8386 11880 8392 11892
rect 8159 11852 8392 11880
rect 8159 11849 8171 11852
rect 8113 11843 8171 11849
rect 8386 11840 8392 11852
rect 8444 11840 8450 11892
rect 9033 11883 9091 11889
rect 9033 11849 9045 11883
rect 9079 11880 9091 11883
rect 10042 11880 10048 11892
rect 9079 11852 10048 11880
rect 9079 11849 9091 11852
rect 9033 11843 9091 11849
rect 10042 11840 10048 11852
rect 10100 11880 10106 11892
rect 10505 11883 10563 11889
rect 10505 11880 10517 11883
rect 10100 11852 10517 11880
rect 10100 11840 10106 11852
rect 10505 11849 10517 11852
rect 10551 11849 10563 11883
rect 10505 11843 10563 11849
rect 11882 11840 11888 11892
rect 11940 11880 11946 11892
rect 12989 11883 13047 11889
rect 12989 11880 13001 11883
rect 11940 11852 13001 11880
rect 11940 11840 11946 11852
rect 12989 11849 13001 11852
rect 13035 11880 13047 11883
rect 19245 11883 19303 11889
rect 13035 11852 14228 11880
rect 13035 11849 13047 11852
rect 12989 11843 13047 11849
rect 14200 11824 14228 11852
rect 19245 11849 19257 11883
rect 19291 11880 19303 11883
rect 19610 11880 19616 11892
rect 19291 11852 19616 11880
rect 19291 11849 19303 11852
rect 19245 11843 19303 11849
rect 19610 11840 19616 11852
rect 19668 11840 19674 11892
rect 20806 11880 20812 11892
rect 20767 11852 20812 11880
rect 20806 11840 20812 11852
rect 20864 11840 20870 11892
rect 21726 11880 21732 11892
rect 21687 11852 21732 11880
rect 21726 11840 21732 11852
rect 21784 11840 21790 11892
rect 4798 11772 4804 11824
rect 4856 11812 4862 11824
rect 5077 11815 5135 11821
rect 5077 11812 5089 11815
rect 4856 11784 5089 11812
rect 4856 11772 4862 11784
rect 5077 11781 5089 11784
rect 5123 11812 5135 11815
rect 5445 11815 5503 11821
rect 5445 11812 5457 11815
rect 5123 11784 5457 11812
rect 5123 11781 5135 11784
rect 5077 11775 5135 11781
rect 5445 11781 5457 11784
rect 5491 11812 5503 11815
rect 5491 11784 7420 11812
rect 5491 11781 5503 11784
rect 5445 11775 5503 11781
rect 1118 11704 1124 11756
rect 1176 11744 1182 11756
rect 1857 11747 1915 11753
rect 1857 11744 1869 11747
rect 1176 11716 1869 11744
rect 1176 11704 1182 11716
rect 1479 11685 1507 11716
rect 1857 11713 1869 11716
rect 1903 11713 1915 11747
rect 1857 11707 1915 11713
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 5537 11747 5595 11753
rect 5537 11744 5549 11747
rect 4764 11716 5549 11744
rect 4764 11704 4770 11716
rect 5537 11713 5549 11716
rect 5583 11713 5595 11747
rect 7392 11744 7420 11784
rect 10226 11772 10232 11824
rect 10284 11812 10290 11824
rect 10321 11815 10379 11821
rect 10321 11812 10333 11815
rect 10284 11784 10333 11812
rect 10284 11772 10290 11784
rect 10321 11781 10333 11784
rect 10367 11781 10379 11815
rect 10321 11775 10379 11781
rect 10336 11744 10364 11775
rect 14182 11772 14188 11824
rect 14240 11812 14246 11824
rect 14645 11815 14703 11821
rect 14645 11812 14657 11815
rect 14240 11784 14657 11812
rect 14240 11772 14246 11784
rect 14645 11781 14657 11784
rect 14691 11812 14703 11815
rect 14691 11784 15608 11812
rect 14691 11781 14703 11784
rect 14645 11775 14703 11781
rect 7392 11716 10364 11744
rect 5537 11707 5595 11713
rect 10410 11704 10416 11756
rect 10468 11744 10474 11756
rect 10468 11716 10513 11744
rect 10468 11704 10474 11716
rect 1464 11679 1522 11685
rect 1464 11645 1476 11679
rect 1510 11645 1522 11679
rect 1464 11639 1522 11645
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11676 2743 11679
rect 2774 11676 2780 11688
rect 2731 11648 2780 11676
rect 2731 11645 2743 11648
rect 2685 11639 2743 11645
rect 2774 11636 2780 11648
rect 2832 11676 2838 11688
rect 4154 11676 4160 11688
rect 2832 11648 4160 11676
rect 2832 11636 2838 11648
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 5350 11685 5356 11688
rect 5316 11679 5356 11685
rect 5316 11676 5328 11679
rect 5263 11648 5328 11676
rect 5316 11645 5328 11648
rect 5408 11676 5414 11688
rect 6362 11676 6368 11688
rect 5408 11648 6368 11676
rect 5316 11639 5356 11645
rect 5350 11636 5356 11639
rect 5408 11636 5414 11648
rect 6362 11636 6368 11648
rect 6420 11636 6426 11688
rect 7098 11676 7104 11688
rect 7059 11648 7104 11676
rect 7098 11636 7104 11648
rect 7156 11636 7162 11688
rect 7282 11636 7288 11688
rect 7340 11676 7346 11688
rect 7469 11679 7527 11685
rect 7469 11676 7481 11679
rect 7340 11648 7481 11676
rect 7340 11636 7346 11648
rect 7469 11645 7481 11648
rect 7515 11645 7527 11679
rect 7834 11676 7840 11688
rect 7747 11648 7840 11676
rect 7469 11639 7527 11645
rect 7834 11636 7840 11648
rect 7892 11676 7898 11688
rect 9674 11676 9680 11688
rect 7892 11648 9680 11676
rect 7892 11636 7898 11648
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 10192 11679 10250 11685
rect 10192 11645 10204 11679
rect 10238 11676 10250 11679
rect 10778 11676 10784 11688
rect 10238 11648 10784 11676
rect 10238 11645 10250 11648
rect 10192 11639 10250 11645
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 11238 11636 11244 11688
rect 11296 11676 11302 11688
rect 11609 11679 11667 11685
rect 11609 11676 11621 11679
rect 11296 11648 11621 11676
rect 11296 11636 11302 11648
rect 11609 11645 11621 11648
rect 11655 11645 11667 11679
rect 13998 11676 14004 11688
rect 13959 11648 14004 11676
rect 11609 11639 11667 11645
rect 13998 11636 14004 11648
rect 14056 11636 14062 11688
rect 15580 11685 15608 11784
rect 16942 11772 16948 11824
rect 17000 11812 17006 11824
rect 21039 11815 21097 11821
rect 21039 11812 21051 11815
rect 17000 11784 21051 11812
rect 17000 11772 17006 11784
rect 21039 11781 21051 11784
rect 21085 11781 21097 11815
rect 21450 11812 21456 11824
rect 21411 11784 21456 11812
rect 21039 11775 21097 11781
rect 21450 11772 21456 11784
rect 21508 11772 21514 11824
rect 15654 11704 15660 11756
rect 15712 11744 15718 11756
rect 15841 11747 15899 11753
rect 15841 11744 15853 11747
rect 15712 11716 15853 11744
rect 15712 11704 15718 11716
rect 15841 11713 15853 11716
rect 15887 11744 15899 11747
rect 16485 11747 16543 11753
rect 16485 11744 16497 11747
rect 15887 11716 16497 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 16485 11713 16497 11716
rect 16531 11713 16543 11747
rect 16485 11707 16543 11713
rect 15381 11679 15439 11685
rect 15381 11645 15393 11679
rect 15427 11645 15439 11679
rect 15381 11639 15439 11645
rect 15565 11679 15623 11685
rect 15565 11645 15577 11679
rect 15611 11645 15623 11679
rect 15565 11639 15623 11645
rect 2593 11611 2651 11617
rect 2593 11577 2605 11611
rect 2639 11608 2651 11611
rect 3047 11611 3105 11617
rect 3047 11608 3059 11611
rect 2639 11580 3059 11608
rect 2639 11577 2651 11580
rect 2593 11571 2651 11577
rect 3047 11577 3059 11580
rect 3093 11608 3105 11611
rect 5169 11611 5227 11617
rect 3093 11580 4200 11608
rect 3093 11577 3105 11580
rect 3047 11571 3105 11577
rect 1535 11543 1593 11549
rect 1535 11509 1547 11543
rect 1581 11540 1593 11543
rect 1670 11540 1676 11552
rect 1581 11512 1676 11540
rect 1581 11509 1593 11512
rect 1535 11503 1593 11509
rect 1670 11500 1676 11512
rect 1728 11500 1734 11552
rect 3602 11540 3608 11552
rect 3563 11512 3608 11540
rect 3602 11500 3608 11512
rect 3660 11500 3666 11552
rect 4172 11549 4200 11580
rect 5169 11577 5181 11611
rect 5215 11608 5227 11611
rect 5718 11608 5724 11620
rect 5215 11580 5724 11608
rect 5215 11577 5227 11580
rect 5169 11571 5227 11577
rect 5718 11568 5724 11580
rect 5776 11568 5782 11620
rect 9309 11611 9367 11617
rect 9309 11608 9321 11611
rect 6288 11580 9321 11608
rect 6288 11552 6316 11580
rect 9309 11577 9321 11580
rect 9355 11608 9367 11611
rect 10042 11608 10048 11620
rect 9355 11580 9904 11608
rect 10003 11580 10048 11608
rect 9355 11577 9367 11580
rect 9309 11571 9367 11577
rect 4157 11543 4215 11549
rect 4157 11509 4169 11543
rect 4203 11540 4215 11543
rect 4430 11540 4436 11552
rect 4203 11512 4436 11540
rect 4203 11509 4215 11512
rect 4157 11503 4215 11509
rect 4430 11500 4436 11512
rect 4488 11500 4494 11552
rect 4706 11540 4712 11552
rect 4667 11512 4712 11540
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 6270 11540 6276 11552
rect 6231 11512 6276 11540
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 6454 11500 6460 11552
rect 6512 11540 6518 11552
rect 6641 11543 6699 11549
rect 6641 11540 6653 11543
rect 6512 11512 6653 11540
rect 6512 11500 6518 11512
rect 6641 11509 6653 11512
rect 6687 11540 6699 11543
rect 7834 11540 7840 11552
rect 6687 11512 7840 11540
rect 6687 11509 6699 11512
rect 6641 11503 6699 11509
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 9674 11540 9680 11552
rect 9635 11512 9680 11540
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 9876 11540 9904 11580
rect 10042 11568 10048 11580
rect 10100 11568 10106 11620
rect 13538 11568 13544 11620
rect 13596 11608 13602 11620
rect 13596 11580 15056 11608
rect 13596 11568 13602 11580
rect 10410 11540 10416 11552
rect 9876 11512 10416 11540
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 10962 11500 10968 11552
rect 11020 11540 11026 11552
rect 11241 11543 11299 11549
rect 11241 11540 11253 11543
rect 11020 11512 11253 11540
rect 11020 11500 11026 11512
rect 11241 11509 11253 11512
rect 11287 11509 11299 11543
rect 11241 11503 11299 11509
rect 11514 11500 11520 11552
rect 11572 11540 11578 11552
rect 11977 11543 12035 11549
rect 11977 11540 11989 11543
rect 11572 11512 11989 11540
rect 11572 11500 11578 11512
rect 11977 11509 11989 11512
rect 12023 11509 12035 11543
rect 12710 11540 12716 11552
rect 12671 11512 12716 11540
rect 11977 11503 12035 11509
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 13354 11540 13360 11552
rect 13315 11512 13360 11540
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 15028 11549 15056 11580
rect 15013 11543 15071 11549
rect 13872 11512 13917 11540
rect 13872 11500 13878 11512
rect 15013 11509 15025 11543
rect 15059 11540 15071 11543
rect 15396 11540 15424 11639
rect 17862 11636 17868 11688
rect 17920 11676 17926 11688
rect 18322 11676 18328 11688
rect 17920 11648 18328 11676
rect 17920 11636 17926 11648
rect 18322 11636 18328 11648
rect 18380 11636 18386 11688
rect 20968 11679 21026 11685
rect 20968 11645 20980 11679
rect 21014 11676 21026 11679
rect 21468 11676 21496 11772
rect 21014 11648 21496 11676
rect 21014 11645 21026 11648
rect 20968 11639 21026 11645
rect 16206 11608 16212 11620
rect 16119 11580 16212 11608
rect 16206 11568 16212 11580
rect 16264 11608 16270 11620
rect 18414 11608 18420 11620
rect 16264 11580 18420 11608
rect 16264 11568 16270 11580
rect 18414 11568 18420 11580
rect 18472 11608 18478 11620
rect 18646 11611 18704 11617
rect 18646 11608 18658 11611
rect 18472 11580 18658 11608
rect 18472 11568 18478 11580
rect 18646 11577 18658 11580
rect 18692 11577 18704 11611
rect 18646 11571 18704 11577
rect 15059 11512 15424 11540
rect 15059 11509 15071 11512
rect 15013 11503 15071 11509
rect 1104 11450 22816 11472
rect 1104 11398 8982 11450
rect 9034 11398 9046 11450
rect 9098 11398 9110 11450
rect 9162 11398 9174 11450
rect 9226 11398 16982 11450
rect 17034 11398 17046 11450
rect 17098 11398 17110 11450
rect 17162 11398 17174 11450
rect 17226 11398 22816 11450
rect 1104 11376 22816 11398
rect 1670 11296 1676 11348
rect 1728 11336 1734 11348
rect 2777 11339 2835 11345
rect 2777 11336 2789 11339
rect 1728 11308 2789 11336
rect 1728 11296 1734 11308
rect 2777 11305 2789 11308
rect 2823 11305 2835 11339
rect 2777 11299 2835 11305
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 4212 11308 4257 11336
rect 4212 11296 4218 11308
rect 4706 11296 4712 11348
rect 4764 11336 4770 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 4764 11308 5181 11336
rect 4764 11296 4770 11308
rect 5169 11305 5181 11308
rect 5215 11336 5227 11339
rect 5350 11336 5356 11348
rect 5215 11308 5356 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 5350 11296 5356 11308
rect 5408 11296 5414 11348
rect 6546 11336 6552 11348
rect 6507 11308 6552 11336
rect 6546 11296 6552 11308
rect 6604 11296 6610 11348
rect 7374 11336 7380 11348
rect 7335 11308 7380 11336
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 10226 11336 10232 11348
rect 10187 11308 10232 11336
rect 10226 11296 10232 11308
rect 10284 11296 10290 11348
rect 12989 11339 13047 11345
rect 12989 11305 13001 11339
rect 13035 11336 13047 11339
rect 15381 11339 15439 11345
rect 15381 11336 15393 11339
rect 13035 11308 15393 11336
rect 13035 11305 13047 11308
rect 12989 11299 13047 11305
rect 1854 11228 1860 11280
rect 1912 11268 1918 11280
rect 1949 11271 2007 11277
rect 1949 11268 1961 11271
rect 1912 11240 1961 11268
rect 1912 11228 1918 11240
rect 1949 11237 1961 11240
rect 1995 11237 2007 11271
rect 1949 11231 2007 11237
rect 3881 11271 3939 11277
rect 3881 11237 3893 11271
rect 3927 11268 3939 11271
rect 4062 11268 4068 11280
rect 3927 11240 4068 11268
rect 3927 11237 3939 11240
rect 3881 11231 3939 11237
rect 4062 11228 4068 11240
rect 4120 11228 4126 11280
rect 5718 11228 5724 11280
rect 5776 11268 5782 11280
rect 5905 11271 5963 11277
rect 5905 11268 5917 11271
rect 5776 11240 5917 11268
rect 5776 11228 5782 11240
rect 5905 11237 5917 11240
rect 5951 11268 5963 11271
rect 7098 11268 7104 11280
rect 5951 11240 7104 11268
rect 5951 11237 5963 11240
rect 5905 11231 5963 11237
rect 7098 11228 7104 11240
rect 7156 11228 7162 11280
rect 8754 11268 8760 11280
rect 8715 11240 8760 11268
rect 8754 11228 8760 11240
rect 8812 11228 8818 11280
rect 11514 11268 11520 11280
rect 9324 11240 11520 11268
rect 4338 11200 4344 11212
rect 4299 11172 4344 11200
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 4522 11200 4528 11212
rect 4483 11172 4528 11200
rect 4522 11160 4528 11172
rect 4580 11160 4586 11212
rect 6052 11203 6110 11209
rect 6052 11169 6064 11203
rect 6098 11200 6110 11203
rect 6362 11200 6368 11212
rect 6098 11172 6368 11200
rect 6098 11169 6110 11172
rect 6052 11163 6110 11169
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 7834 11160 7840 11212
rect 7892 11200 7898 11212
rect 8021 11203 8079 11209
rect 8021 11200 8033 11203
rect 7892 11172 8033 11200
rect 7892 11160 7898 11172
rect 8021 11169 8033 11172
rect 8067 11200 8079 11203
rect 9324 11200 9352 11240
rect 11514 11228 11520 11240
rect 11572 11228 11578 11280
rect 11698 11268 11704 11280
rect 11659 11240 11704 11268
rect 11698 11228 11704 11240
rect 11756 11228 11762 11280
rect 8067 11172 9352 11200
rect 8067 11169 8079 11172
rect 8021 11163 8079 11169
rect 9398 11160 9404 11212
rect 9456 11200 9462 11212
rect 9712 11203 9770 11209
rect 9712 11200 9724 11203
rect 9456 11172 9724 11200
rect 9456 11160 9462 11172
rect 9712 11169 9724 11172
rect 9758 11169 9770 11203
rect 9712 11163 9770 11169
rect 10042 11160 10048 11212
rect 10100 11200 10106 11212
rect 10686 11200 10692 11212
rect 10100 11172 10692 11200
rect 10100 11160 10106 11172
rect 10686 11160 10692 11172
rect 10744 11200 10750 11212
rect 10965 11203 11023 11209
rect 10965 11200 10977 11203
rect 10744 11172 10977 11200
rect 10744 11160 10750 11172
rect 10965 11169 10977 11172
rect 11011 11169 11023 11203
rect 11532 11200 11560 11228
rect 12437 11203 12495 11209
rect 12437 11200 12449 11203
rect 11532 11172 12449 11200
rect 10965 11163 11023 11169
rect 12437 11169 12449 11172
rect 12483 11200 12495 11203
rect 12526 11200 12532 11212
rect 12483 11172 12532 11200
rect 12483 11169 12495 11172
rect 12437 11163 12495 11169
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11132 1915 11135
rect 1946 11132 1952 11144
rect 1903 11104 1952 11132
rect 1903 11101 1915 11104
rect 1857 11095 1915 11101
rect 1946 11092 1952 11104
rect 2004 11092 2010 11144
rect 6270 11132 6276 11144
rect 6231 11104 6276 11132
rect 6270 11092 6276 11104
rect 6328 11092 6334 11144
rect 7926 11092 7932 11144
rect 7984 11132 7990 11144
rect 8389 11135 8447 11141
rect 8389 11132 8401 11135
rect 7984 11104 8401 11132
rect 7984 11092 7990 11104
rect 8389 11101 8401 11104
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 1673 11067 1731 11073
rect 1673 11033 1685 11067
rect 1719 11064 1731 11067
rect 1762 11064 1768 11076
rect 1719 11036 1768 11064
rect 1719 11033 1731 11036
rect 1673 11027 1731 11033
rect 1762 11024 1768 11036
rect 1820 11024 1826 11076
rect 2409 11067 2467 11073
rect 2409 11033 2421 11067
rect 2455 11064 2467 11067
rect 2590 11064 2596 11076
rect 2455 11036 2596 11064
rect 2455 11033 2467 11036
rect 2409 11027 2467 11033
rect 2590 11024 2596 11036
rect 2648 11064 2654 11076
rect 6730 11064 6736 11076
rect 2648 11036 6736 11064
rect 2648 11024 2654 11036
rect 6730 11024 6736 11036
rect 6788 11024 6794 11076
rect 6914 11024 6920 11076
rect 6972 11064 6978 11076
rect 9815 11067 9873 11073
rect 9815 11064 9827 11067
rect 6972 11036 9827 11064
rect 6972 11024 6978 11036
rect 9815 11033 9827 11036
rect 9861 11033 9873 11067
rect 10980 11064 11008 11163
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 13096 11209 13124 11308
rect 15381 11305 15393 11308
rect 15427 11305 15439 11339
rect 18414 11336 18420 11348
rect 18375 11308 18420 11336
rect 15381 11299 15439 11305
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 13334 11271 13392 11277
rect 13334 11237 13346 11271
rect 13380 11268 13392 11271
rect 13446 11268 13452 11280
rect 13380 11240 13452 11268
rect 13380 11237 13392 11240
rect 13334 11231 13392 11237
rect 13446 11228 13452 11240
rect 13504 11228 13510 11280
rect 17862 11268 17868 11280
rect 17823 11240 17868 11268
rect 17862 11228 17868 11240
rect 17920 11228 17926 11280
rect 13081 11203 13139 11209
rect 13081 11169 13093 11203
rect 13127 11169 13139 11203
rect 13998 11200 14004 11212
rect 13959 11172 14004 11200
rect 13081 11163 13139 11169
rect 13998 11160 14004 11172
rect 14056 11200 14062 11212
rect 14277 11203 14335 11209
rect 14277 11200 14289 11203
rect 14056 11172 14289 11200
rect 14056 11160 14062 11172
rect 14277 11169 14289 11172
rect 14323 11169 14335 11203
rect 15378 11200 15384 11212
rect 15339 11172 15384 11200
rect 14277 11163 14335 11169
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 15838 11200 15844 11212
rect 15799 11172 15844 11200
rect 15838 11160 15844 11172
rect 15896 11160 15902 11212
rect 17405 11203 17463 11209
rect 17405 11169 17417 11203
rect 17451 11169 17463 11203
rect 17586 11200 17592 11212
rect 17547 11172 17592 11200
rect 17405 11163 17463 11169
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 11333 11135 11391 11141
rect 11333 11132 11345 11135
rect 11112 11104 11345 11132
rect 11112 11092 11118 11104
rect 11333 11101 11345 11104
rect 11379 11101 11391 11135
rect 17420 11132 17448 11163
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 17494 11132 17500 11144
rect 17420 11104 17500 11132
rect 11333 11095 11391 11101
rect 17494 11092 17500 11104
rect 17552 11092 17558 11144
rect 10980 11036 11376 11064
rect 9815 11027 9873 11033
rect 11348 11008 11376 11036
rect 5442 10956 5448 11008
rect 5500 10996 5506 11008
rect 5721 10999 5779 11005
rect 5721 10996 5733 10999
rect 5500 10968 5733 10996
rect 5500 10956 5506 10968
rect 5721 10965 5733 10968
rect 5767 10996 5779 10999
rect 6086 10996 6092 11008
rect 5767 10968 6092 10996
rect 5767 10965 5779 10968
rect 5721 10959 5779 10965
rect 6086 10956 6092 10968
rect 6144 10996 6150 11008
rect 6181 10999 6239 11005
rect 6181 10996 6193 10999
rect 6144 10968 6193 10996
rect 6144 10956 6150 10968
rect 6181 10965 6193 10968
rect 6227 10996 6239 10999
rect 6546 10996 6552 11008
rect 6227 10968 6552 10996
rect 6227 10965 6239 10968
rect 6181 10959 6239 10965
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 7098 10996 7104 11008
rect 7059 10968 7104 10996
rect 7098 10956 7104 10968
rect 7156 10956 7162 11008
rect 7837 10999 7895 11005
rect 7837 10965 7849 10999
rect 7883 10996 7895 10999
rect 8018 10996 8024 11008
rect 7883 10968 8024 10996
rect 7883 10965 7895 10968
rect 7837 10959 7895 10965
rect 8018 10956 8024 10968
rect 8076 10956 8082 11008
rect 8202 11005 8208 11008
rect 8186 10999 8208 11005
rect 8186 10965 8198 10999
rect 8186 10959 8208 10965
rect 8202 10956 8208 10959
rect 8260 10956 8266 11008
rect 8297 10999 8355 11005
rect 8297 10965 8309 10999
rect 8343 10996 8355 10999
rect 8478 10996 8484 11008
rect 8343 10968 8484 10996
rect 8343 10965 8355 10968
rect 8297 10959 8355 10965
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 9398 10996 9404 11008
rect 9359 10968 9404 10996
rect 9398 10956 9404 10968
rect 9456 10956 9462 11008
rect 10505 10999 10563 11005
rect 10505 10965 10517 10999
rect 10551 10996 10563 10999
rect 10778 10996 10784 11008
rect 10551 10968 10784 10996
rect 10551 10965 10563 10968
rect 10505 10959 10563 10965
rect 10778 10956 10784 10968
rect 10836 10996 10842 11008
rect 11103 10999 11161 11005
rect 11103 10996 11115 10999
rect 10836 10968 11115 10996
rect 10836 10956 10842 10968
rect 11103 10965 11115 10968
rect 11149 10965 11161 10999
rect 11238 10996 11244 11008
rect 11199 10968 11244 10996
rect 11103 10959 11161 10965
rect 11238 10956 11244 10968
rect 11296 10956 11302 11008
rect 11330 10956 11336 11008
rect 11388 10996 11394 11008
rect 11977 10999 12035 11005
rect 11977 10996 11989 10999
rect 11388 10968 11989 10996
rect 11388 10956 11394 10968
rect 11977 10965 11989 10968
rect 12023 10965 12035 10999
rect 11977 10959 12035 10965
rect 1104 10906 22816 10928
rect 1104 10854 4982 10906
rect 5034 10854 5046 10906
rect 5098 10854 5110 10906
rect 5162 10854 5174 10906
rect 5226 10854 12982 10906
rect 13034 10854 13046 10906
rect 13098 10854 13110 10906
rect 13162 10854 13174 10906
rect 13226 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 22816 10906
rect 1104 10832 22816 10854
rect 3421 10795 3479 10801
rect 3421 10761 3433 10795
rect 3467 10792 3479 10795
rect 4522 10792 4528 10804
rect 3467 10764 4528 10792
rect 3467 10761 3479 10764
rect 3421 10755 3479 10761
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 4985 10795 5043 10801
rect 4985 10792 4997 10795
rect 4856 10764 4997 10792
rect 4856 10752 4862 10764
rect 4985 10761 4997 10764
rect 5031 10761 5043 10795
rect 4985 10755 5043 10761
rect 5334 10795 5392 10801
rect 5334 10761 5346 10795
rect 5380 10792 5392 10795
rect 5626 10792 5632 10804
rect 5380 10764 5632 10792
rect 5380 10761 5392 10764
rect 5334 10755 5392 10761
rect 2590 10724 2596 10736
rect 2551 10696 2596 10724
rect 2590 10684 2596 10696
rect 2648 10684 2654 10736
rect 5000 10724 5028 10755
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 6546 10792 6552 10804
rect 6507 10764 6552 10792
rect 6546 10752 6552 10764
rect 6604 10792 6610 10804
rect 7193 10795 7251 10801
rect 7193 10792 7205 10795
rect 6604 10764 7205 10792
rect 6604 10752 6610 10764
rect 7193 10761 7205 10764
rect 7239 10792 7251 10795
rect 8478 10792 8484 10804
rect 7239 10764 8484 10792
rect 7239 10761 7251 10764
rect 7193 10755 7251 10761
rect 8478 10752 8484 10764
rect 8536 10752 8542 10804
rect 13446 10792 13452 10804
rect 13407 10764 13452 10792
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 13909 10795 13967 10801
rect 13909 10761 13921 10795
rect 13955 10792 13967 10795
rect 13998 10792 14004 10804
rect 13955 10764 14004 10792
rect 13955 10761 13967 10764
rect 13909 10755 13967 10761
rect 13998 10752 14004 10764
rect 14056 10752 14062 10804
rect 14182 10752 14188 10804
rect 14240 10792 14246 10804
rect 15289 10795 15347 10801
rect 15289 10792 15301 10795
rect 14240 10764 15301 10792
rect 14240 10752 14246 10764
rect 15289 10761 15301 10764
rect 15335 10792 15347 10795
rect 15378 10792 15384 10804
rect 15335 10764 15384 10792
rect 15335 10761 15347 10764
rect 15289 10755 15347 10761
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 5445 10727 5503 10733
rect 5445 10724 5457 10727
rect 5000 10696 5457 10724
rect 5445 10693 5457 10696
rect 5491 10693 5503 10727
rect 7561 10727 7619 10733
rect 7561 10724 7573 10727
rect 5445 10687 5503 10693
rect 5552 10696 7573 10724
rect 1854 10656 1860 10668
rect 1767 10628 1860 10656
rect 1854 10616 1860 10628
rect 1912 10656 1918 10668
rect 3513 10659 3571 10665
rect 3513 10656 3525 10659
rect 1912 10628 3525 10656
rect 1912 10616 1918 10628
rect 3513 10625 3525 10628
rect 3559 10625 3571 10659
rect 3513 10619 3571 10625
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 4525 10659 4583 10665
rect 4525 10656 4537 10659
rect 4396 10628 4537 10656
rect 4396 10616 4402 10628
rect 4525 10625 4537 10628
rect 4571 10625 4583 10659
rect 4525 10619 4583 10625
rect 5350 10616 5356 10668
rect 5408 10656 5414 10668
rect 5552 10665 5580 10696
rect 7561 10693 7573 10696
rect 7607 10724 7619 10727
rect 7926 10724 7932 10736
rect 7607 10696 7932 10724
rect 7607 10693 7619 10696
rect 7561 10687 7619 10693
rect 7926 10684 7932 10696
rect 7984 10724 7990 10736
rect 10962 10724 10968 10736
rect 7984 10696 10968 10724
rect 7984 10684 7990 10696
rect 10962 10684 10968 10696
rect 11020 10684 11026 10736
rect 12713 10727 12771 10733
rect 12713 10724 12725 10727
rect 12360 10696 12725 10724
rect 5537 10659 5595 10665
rect 5537 10656 5549 10659
rect 5408 10628 5549 10656
rect 5408 10616 5414 10628
rect 5537 10625 5549 10628
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 3053 10591 3111 10597
rect 3053 10557 3065 10591
rect 3099 10588 3111 10591
rect 3602 10588 3608 10600
rect 3099 10560 3608 10588
rect 3099 10557 3111 10560
rect 3053 10551 3111 10557
rect 2038 10520 2044 10532
rect 1999 10492 2044 10520
rect 2038 10480 2044 10492
rect 2096 10480 2102 10532
rect 2133 10523 2191 10529
rect 2133 10489 2145 10523
rect 2179 10520 2191 10523
rect 3068 10520 3096 10551
rect 3602 10548 3608 10560
rect 3660 10548 3666 10600
rect 4246 10548 4252 10600
rect 4304 10588 4310 10600
rect 5644 10588 5672 10619
rect 9398 10616 9404 10668
rect 9456 10656 9462 10668
rect 9861 10659 9919 10665
rect 9861 10656 9873 10659
rect 9456 10628 9873 10656
rect 9456 10616 9462 10628
rect 9861 10625 9873 10628
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 7742 10588 7748 10600
rect 4304 10560 5672 10588
rect 7703 10560 7748 10588
rect 4304 10548 4310 10560
rect 7742 10548 7748 10560
rect 7800 10548 7806 10600
rect 8665 10591 8723 10597
rect 8665 10557 8677 10591
rect 8711 10588 8723 10591
rect 9309 10591 9367 10597
rect 9309 10588 9321 10591
rect 8711 10560 9321 10588
rect 8711 10557 8723 10560
rect 8665 10551 8723 10557
rect 9309 10557 9321 10560
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 11400 10591 11458 10597
rect 11400 10557 11412 10591
rect 11446 10588 11458 10591
rect 12158 10588 12164 10600
rect 11446 10560 12164 10588
rect 11446 10557 11458 10560
rect 11400 10551 11458 10557
rect 2179 10492 3096 10520
rect 5169 10523 5227 10529
rect 2179 10489 2191 10492
rect 2133 10483 2191 10489
rect 5169 10489 5181 10523
rect 5215 10520 5227 10523
rect 5534 10520 5540 10532
rect 5215 10492 5540 10520
rect 5215 10489 5227 10492
rect 5169 10483 5227 10489
rect 5534 10480 5540 10492
rect 5592 10480 5598 10532
rect 7834 10480 7840 10532
rect 7892 10520 7898 10532
rect 8941 10523 8999 10529
rect 8941 10520 8953 10523
rect 7892 10492 8953 10520
rect 7892 10480 7898 10492
rect 8941 10489 8953 10492
rect 8987 10489 8999 10523
rect 8941 10483 8999 10489
rect 6270 10452 6276 10464
rect 6231 10424 6276 10452
rect 6270 10412 6276 10424
rect 6328 10412 6334 10464
rect 8018 10412 8024 10464
rect 8076 10452 8082 10464
rect 8113 10455 8171 10461
rect 8113 10452 8125 10455
rect 8076 10424 8125 10452
rect 8076 10412 8082 10424
rect 8113 10421 8125 10424
rect 8159 10421 8171 10455
rect 9324 10452 9352 10551
rect 12158 10548 12164 10560
rect 12216 10548 12222 10600
rect 9582 10520 9588 10532
rect 9543 10492 9588 10520
rect 9582 10480 9588 10492
rect 9640 10480 9646 10532
rect 9677 10523 9735 10529
rect 9677 10489 9689 10523
rect 9723 10489 9735 10523
rect 9677 10483 9735 10489
rect 9692 10452 9720 10483
rect 11238 10480 11244 10532
rect 11296 10520 11302 10532
rect 11793 10523 11851 10529
rect 11793 10520 11805 10523
rect 11296 10492 11805 10520
rect 11296 10480 11302 10492
rect 11793 10489 11805 10492
rect 11839 10489 11851 10523
rect 11793 10483 11851 10489
rect 9766 10452 9772 10464
rect 9324 10424 9772 10452
rect 8113 10415 8171 10421
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 10689 10455 10747 10461
rect 10689 10421 10701 10455
rect 10735 10452 10747 10455
rect 10778 10452 10784 10464
rect 10735 10424 10784 10452
rect 10735 10421 10747 10424
rect 10689 10415 10747 10421
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 11471 10455 11529 10461
rect 11471 10421 11483 10455
rect 11517 10452 11529 10455
rect 11698 10452 11704 10464
rect 11517 10424 11704 10452
rect 11517 10421 11529 10424
rect 11471 10415 11529 10421
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 11882 10412 11888 10464
rect 11940 10452 11946 10464
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 11940 10424 12173 10452
rect 11940 10412 11946 10424
rect 12161 10421 12173 10424
rect 12207 10452 12219 10455
rect 12360 10452 12388 10696
rect 12713 10693 12725 10696
rect 12759 10693 12771 10727
rect 12713 10687 12771 10693
rect 13081 10727 13139 10733
rect 13081 10693 13093 10727
rect 13127 10724 13139 10727
rect 15838 10724 15844 10736
rect 13127 10696 15844 10724
rect 13127 10693 13139 10696
rect 13081 10687 13139 10693
rect 15838 10684 15844 10696
rect 15896 10724 15902 10736
rect 16025 10727 16083 10733
rect 16025 10724 16037 10727
rect 15896 10696 16037 10724
rect 15896 10684 15902 10696
rect 16025 10693 16037 10696
rect 16071 10724 16083 10727
rect 17497 10727 17555 10733
rect 17497 10724 17509 10727
rect 16071 10696 17509 10724
rect 16071 10693 16083 10696
rect 16025 10687 16083 10693
rect 17497 10693 17509 10696
rect 17543 10724 17555 10727
rect 17586 10724 17592 10736
rect 17543 10696 17592 10724
rect 17543 10693 17555 10696
rect 17497 10687 17555 10693
rect 17586 10684 17592 10696
rect 17644 10684 17650 10736
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 12805 10659 12863 10665
rect 12805 10656 12817 10659
rect 12492 10628 12817 10656
rect 12492 10616 12498 10628
rect 12805 10625 12817 10628
rect 12851 10625 12863 10659
rect 12805 10619 12863 10625
rect 13354 10616 13360 10668
rect 13412 10656 13418 10668
rect 14182 10656 14188 10668
rect 13412 10628 14188 10656
rect 13412 10616 13418 10628
rect 14182 10616 14188 10628
rect 14240 10616 14246 10668
rect 14366 10656 14372 10668
rect 14327 10628 14372 10656
rect 14366 10616 14372 10628
rect 14424 10616 14430 10668
rect 12584 10591 12642 10597
rect 12584 10557 12596 10591
rect 12630 10588 12642 10591
rect 12710 10588 12716 10600
rect 12630 10560 12716 10588
rect 12630 10557 12642 10560
rect 12584 10551 12642 10557
rect 12710 10548 12716 10560
rect 12768 10548 12774 10600
rect 19150 10548 19156 10600
rect 19208 10588 19214 10600
rect 19889 10591 19947 10597
rect 19889 10588 19901 10591
rect 19208 10560 19901 10588
rect 19208 10548 19214 10560
rect 19889 10557 19901 10560
rect 19935 10588 19947 10591
rect 20622 10588 20628 10600
rect 19935 10560 20628 10588
rect 19935 10557 19947 10560
rect 19889 10551 19947 10557
rect 20622 10548 20628 10560
rect 20680 10548 20686 10600
rect 21612 10591 21670 10597
rect 21612 10557 21624 10591
rect 21658 10588 21670 10591
rect 22094 10588 22100 10600
rect 21658 10560 22100 10588
rect 21658 10557 21670 10560
rect 21612 10551 21670 10557
rect 22094 10548 22100 10560
rect 22152 10548 22158 10600
rect 12437 10523 12495 10529
rect 12437 10489 12449 10523
rect 12483 10489 12495 10523
rect 14090 10520 14096 10532
rect 14051 10492 14096 10520
rect 12437 10483 12495 10489
rect 12207 10424 12388 10452
rect 12452 10452 12480 10483
rect 14090 10480 14096 10492
rect 14148 10480 14154 10532
rect 14185 10523 14243 10529
rect 14185 10489 14197 10523
rect 14231 10489 14243 10523
rect 14185 10483 14243 10489
rect 12526 10452 12532 10464
rect 12452 10424 12532 10452
rect 12207 10421 12219 10424
rect 12161 10415 12219 10421
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 13998 10412 14004 10464
rect 14056 10452 14062 10464
rect 14200 10452 14228 10483
rect 14056 10424 14228 10452
rect 14056 10412 14062 10424
rect 14458 10412 14464 10464
rect 14516 10452 14522 10464
rect 15565 10455 15623 10461
rect 15565 10452 15577 10455
rect 14516 10424 15577 10452
rect 14516 10412 14522 10424
rect 15565 10421 15577 10424
rect 15611 10421 15623 10455
rect 15565 10415 15623 10421
rect 17221 10455 17279 10461
rect 17221 10421 17233 10455
rect 17267 10452 17279 10455
rect 17494 10452 17500 10464
rect 17267 10424 17500 10452
rect 17267 10421 17279 10424
rect 17221 10415 17279 10421
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 20254 10452 20260 10464
rect 20215 10424 20260 10452
rect 20254 10412 20260 10424
rect 20312 10412 20318 10464
rect 20530 10412 20536 10464
rect 20588 10452 20594 10464
rect 21683 10455 21741 10461
rect 21683 10452 21695 10455
rect 20588 10424 21695 10452
rect 20588 10412 20594 10424
rect 21683 10421 21695 10424
rect 21729 10421 21741 10455
rect 22094 10452 22100 10464
rect 22055 10424 22100 10452
rect 21683 10415 21741 10421
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 1104 10362 22816 10384
rect 1104 10310 8982 10362
rect 9034 10310 9046 10362
rect 9098 10310 9110 10362
rect 9162 10310 9174 10362
rect 9226 10310 16982 10362
rect 17034 10310 17046 10362
rect 17098 10310 17110 10362
rect 17162 10310 17174 10362
rect 17226 10310 22816 10362
rect 1104 10288 22816 10310
rect 2038 10208 2044 10260
rect 2096 10248 2102 10260
rect 3145 10251 3203 10257
rect 3145 10248 3157 10251
rect 2096 10220 3157 10248
rect 2096 10208 2102 10220
rect 3145 10217 3157 10220
rect 3191 10217 3203 10251
rect 3602 10248 3608 10260
rect 3563 10220 3608 10248
rect 3145 10211 3203 10217
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 4341 10251 4399 10257
rect 4341 10248 4353 10251
rect 4120 10220 4353 10248
rect 4120 10208 4126 10220
rect 4341 10217 4353 10220
rect 4387 10217 4399 10251
rect 4341 10211 4399 10217
rect 5353 10251 5411 10257
rect 5353 10217 5365 10251
rect 5399 10248 5411 10251
rect 5534 10248 5540 10260
rect 5399 10220 5540 10248
rect 5399 10217 5411 10220
rect 5353 10211 5411 10217
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 5626 10208 5632 10260
rect 5684 10248 5690 10260
rect 5684 10220 5729 10248
rect 5684 10208 5690 10220
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 7800 10220 7941 10248
rect 7800 10208 7806 10220
rect 7929 10217 7941 10220
rect 7975 10248 7987 10251
rect 8757 10251 8815 10257
rect 8757 10248 8769 10251
rect 7975 10220 8769 10248
rect 7975 10217 7987 10220
rect 7929 10211 7987 10217
rect 8757 10217 8769 10220
rect 8803 10217 8815 10251
rect 8757 10211 8815 10217
rect 12710 10208 12716 10260
rect 12768 10248 12774 10260
rect 12805 10251 12863 10257
rect 12805 10248 12817 10251
rect 12768 10220 12817 10248
rect 12768 10208 12774 10220
rect 12805 10217 12817 10220
rect 12851 10217 12863 10251
rect 12805 10211 12863 10217
rect 13446 10208 13452 10260
rect 13504 10248 13510 10260
rect 13906 10248 13912 10260
rect 13504 10220 13912 10248
rect 13504 10208 13510 10220
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 14090 10208 14096 10260
rect 14148 10248 14154 10260
rect 14737 10251 14795 10257
rect 14737 10248 14749 10251
rect 14148 10220 14749 10248
rect 14148 10208 14154 10220
rect 14737 10217 14749 10220
rect 14783 10248 14795 10251
rect 15746 10248 15752 10260
rect 14783 10220 15752 10248
rect 14783 10217 14795 10220
rect 14737 10211 14795 10217
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 3786 10140 3792 10192
rect 3844 10180 3850 10192
rect 4154 10180 4160 10192
rect 3844 10152 4160 10180
rect 3844 10140 3850 10152
rect 4154 10140 4160 10152
rect 4212 10180 4218 10192
rect 4212 10152 4752 10180
rect 4212 10140 4218 10152
rect 2038 10072 2044 10124
rect 2096 10112 2102 10124
rect 2225 10115 2283 10121
rect 2225 10112 2237 10115
rect 2096 10084 2237 10112
rect 2096 10072 2102 10084
rect 2225 10081 2237 10084
rect 2271 10081 2283 10115
rect 4338 10112 4344 10124
rect 4299 10084 4344 10112
rect 2225 10075 2283 10081
rect 4338 10072 4344 10084
rect 4396 10072 4402 10124
rect 4724 10121 4752 10152
rect 7208 10152 7788 10180
rect 4709 10115 4767 10121
rect 4709 10081 4721 10115
rect 4755 10081 4767 10115
rect 5810 10112 5816 10124
rect 5771 10084 5816 10112
rect 4709 10075 4767 10081
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 6733 10115 6791 10121
rect 6733 10081 6745 10115
rect 6779 10112 6791 10115
rect 7098 10112 7104 10124
rect 6779 10084 7104 10112
rect 6779 10081 6791 10084
rect 6733 10075 6791 10081
rect 7098 10072 7104 10084
rect 7156 10112 7162 10124
rect 7208 10121 7236 10152
rect 7760 10124 7788 10152
rect 8662 10140 8668 10192
rect 8720 10180 8726 10192
rect 9401 10183 9459 10189
rect 9401 10180 9413 10183
rect 8720 10152 9413 10180
rect 8720 10140 8726 10152
rect 9401 10149 9413 10152
rect 9447 10180 9459 10183
rect 9582 10180 9588 10192
rect 9447 10152 9588 10180
rect 9447 10149 9459 10152
rect 9401 10143 9459 10149
rect 9582 10140 9588 10152
rect 9640 10140 9646 10192
rect 13814 10140 13820 10192
rect 13872 10180 13878 10192
rect 14366 10180 14372 10192
rect 13872 10152 13917 10180
rect 14327 10152 14372 10180
rect 13872 10140 13878 10152
rect 14366 10140 14372 10152
rect 14424 10140 14430 10192
rect 20622 10140 20628 10192
rect 20680 10180 20686 10192
rect 21085 10183 21143 10189
rect 21085 10180 21097 10183
rect 20680 10152 21097 10180
rect 20680 10140 20686 10152
rect 21085 10149 21097 10152
rect 21131 10180 21143 10183
rect 21450 10180 21456 10192
rect 21131 10152 21456 10180
rect 21131 10149 21143 10152
rect 21085 10143 21143 10149
rect 21450 10140 21456 10152
rect 21508 10140 21514 10192
rect 7193 10115 7251 10121
rect 7193 10112 7205 10115
rect 7156 10084 7205 10112
rect 7156 10072 7162 10084
rect 7193 10081 7205 10084
rect 7239 10081 7251 10115
rect 7193 10075 7251 10081
rect 7282 10072 7288 10124
rect 7340 10112 7346 10124
rect 7469 10115 7527 10121
rect 7469 10112 7481 10115
rect 7340 10084 7481 10112
rect 7340 10072 7346 10084
rect 7469 10081 7481 10084
rect 7515 10081 7527 10115
rect 7469 10075 7527 10081
rect 7742 10072 7748 10124
rect 7800 10072 7806 10124
rect 7837 10115 7895 10121
rect 7837 10081 7849 10115
rect 7883 10112 7895 10115
rect 7926 10112 7932 10124
rect 7883 10084 7932 10112
rect 7883 10081 7895 10084
rect 7837 10075 7895 10081
rect 7926 10072 7932 10084
rect 7984 10072 7990 10124
rect 9766 10112 9772 10124
rect 9727 10084 9772 10112
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 10226 10072 10232 10124
rect 10284 10112 10290 10124
rect 11333 10115 11391 10121
rect 11333 10112 11345 10115
rect 10284 10084 11345 10112
rect 10284 10072 10290 10084
rect 11333 10081 11345 10084
rect 11379 10112 11391 10115
rect 11790 10112 11796 10124
rect 11379 10084 11796 10112
rect 11379 10081 11391 10084
rect 11333 10075 11391 10081
rect 11790 10072 11796 10084
rect 11848 10072 11854 10124
rect 15930 10112 15936 10124
rect 15891 10084 15936 10112
rect 15930 10072 15936 10084
rect 15988 10072 15994 10124
rect 17405 10115 17463 10121
rect 17405 10081 17417 10115
rect 17451 10081 17463 10115
rect 17586 10112 17592 10124
rect 17547 10084 17592 10112
rect 17405 10075 17463 10081
rect 2130 10044 2136 10056
rect 2091 10016 2136 10044
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 6362 10004 6368 10056
rect 6420 10044 6426 10056
rect 8202 10044 8208 10056
rect 6420 10016 8208 10044
rect 6420 10004 6426 10016
rect 8202 10004 8208 10016
rect 8260 10044 8266 10056
rect 8389 10047 8447 10053
rect 8389 10044 8401 10047
rect 8260 10016 8401 10044
rect 8260 10004 8266 10016
rect 8389 10013 8401 10016
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8570 10004 8576 10056
rect 8628 10044 8634 10056
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 8628 10016 9689 10044
rect 8628 10004 8634 10016
rect 9677 10013 9689 10016
rect 9723 10013 9735 10047
rect 11054 10044 11060 10056
rect 9677 10007 9735 10013
rect 10796 10016 11060 10044
rect 1857 9979 1915 9985
rect 1857 9945 1869 9979
rect 1903 9976 1915 9979
rect 1946 9976 1952 9988
rect 1903 9948 1952 9976
rect 1903 9945 1915 9948
rect 1857 9939 1915 9945
rect 1946 9936 1952 9948
rect 2004 9976 2010 9988
rect 6822 9976 6828 9988
rect 2004 9948 6828 9976
rect 2004 9936 2010 9948
rect 6822 9936 6828 9948
rect 6880 9936 6886 9988
rect 8478 9936 8484 9988
rect 8536 9976 8542 9988
rect 10796 9985 10824 10016
rect 11054 10004 11060 10016
rect 11112 10044 11118 10056
rect 11238 10044 11244 10056
rect 11112 10016 11244 10044
rect 11112 10004 11118 10016
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 12158 10004 12164 10056
rect 12216 10044 12222 10056
rect 13725 10047 13783 10053
rect 12216 10016 13486 10044
rect 12216 10004 12222 10016
rect 10781 9979 10839 9985
rect 10781 9976 10793 9979
rect 8536 9948 10793 9976
rect 8536 9936 8542 9948
rect 10781 9945 10793 9948
rect 10827 9945 10839 9979
rect 10781 9939 10839 9945
rect 11422 9936 11428 9988
rect 11480 9976 11486 9988
rect 13173 9979 13231 9985
rect 13173 9976 13185 9979
rect 11480 9948 13185 9976
rect 11480 9936 11486 9948
rect 13173 9945 13185 9948
rect 13219 9945 13231 9979
rect 13458 9976 13486 10016
rect 13725 10013 13737 10047
rect 13771 10044 13783 10047
rect 14458 10044 14464 10056
rect 13771 10016 14464 10044
rect 13771 10013 13783 10016
rect 13725 10007 13783 10013
rect 14458 10004 14464 10016
rect 14516 10004 14522 10056
rect 15378 10044 15384 10056
rect 15339 10016 15384 10044
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 17420 10044 17448 10075
rect 17586 10072 17592 10084
rect 17644 10072 17650 10124
rect 17494 10044 17500 10056
rect 17420 10016 17500 10044
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 17862 10044 17868 10056
rect 17823 10016 17868 10044
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 20993 10047 21051 10053
rect 20993 10013 21005 10047
rect 21039 10044 21051 10047
rect 21818 10044 21824 10056
rect 21039 10016 21824 10044
rect 21039 10013 21051 10016
rect 20993 10007 21051 10013
rect 21818 10004 21824 10016
rect 21876 10004 21882 10056
rect 14366 9976 14372 9988
rect 13458 9948 14372 9976
rect 13173 9939 13231 9945
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 5951 9911 6009 9917
rect 5951 9908 5963 9911
rect 5776 9880 5963 9908
rect 5776 9868 5782 9880
rect 5951 9877 5963 9880
rect 5997 9877 6009 9911
rect 6362 9908 6368 9920
rect 6323 9880 6368 9908
rect 5951 9871 6009 9877
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 12434 9908 12440 9920
rect 12395 9880 12440 9908
rect 12434 9868 12440 9880
rect 12492 9868 12498 9920
rect 13188 9908 13216 9939
rect 14366 9936 14372 9948
rect 14424 9936 14430 9988
rect 21542 9976 21548 9988
rect 21503 9948 21548 9976
rect 21542 9936 21548 9948
rect 21600 9936 21606 9988
rect 13630 9908 13636 9920
rect 13188 9880 13636 9908
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 1104 9818 22816 9840
rect 1104 9766 4982 9818
rect 5034 9766 5046 9818
rect 5098 9766 5110 9818
rect 5162 9766 5174 9818
rect 5226 9766 12982 9818
rect 13034 9766 13046 9818
rect 13098 9766 13110 9818
rect 13162 9766 13174 9818
rect 13226 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 22816 9818
rect 1104 9744 22816 9766
rect 2130 9704 2136 9716
rect 2091 9676 2136 9704
rect 2130 9664 2136 9676
rect 2188 9664 2194 9716
rect 3786 9704 3792 9716
rect 3747 9676 3792 9704
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 4157 9707 4215 9713
rect 4157 9673 4169 9707
rect 4203 9704 4215 9707
rect 4338 9704 4344 9716
rect 4203 9676 4344 9704
rect 4203 9673 4215 9676
rect 4157 9667 4215 9673
rect 4338 9664 4344 9676
rect 4396 9664 4402 9716
rect 5810 9704 5816 9716
rect 5771 9676 5816 9704
rect 5810 9664 5816 9676
rect 5868 9664 5874 9716
rect 6641 9707 6699 9713
rect 6641 9673 6653 9707
rect 6687 9704 6699 9707
rect 7282 9704 7288 9716
rect 6687 9676 7288 9704
rect 6687 9673 6699 9676
rect 6641 9667 6699 9673
rect 7282 9664 7288 9676
rect 7340 9664 7346 9716
rect 9585 9707 9643 9713
rect 9585 9673 9597 9707
rect 9631 9704 9643 9707
rect 9766 9704 9772 9716
rect 9631 9676 9772 9704
rect 9631 9673 9643 9676
rect 9585 9667 9643 9673
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 10410 9664 10416 9716
rect 10468 9704 10474 9716
rect 10597 9707 10655 9713
rect 10597 9704 10609 9707
rect 10468 9676 10609 9704
rect 10468 9664 10474 9676
rect 10597 9673 10609 9676
rect 10643 9673 10655 9707
rect 11054 9704 11060 9716
rect 11015 9676 11060 9704
rect 10597 9667 10655 9673
rect 2314 9596 2320 9648
rect 2372 9636 2378 9648
rect 2961 9639 3019 9645
rect 2961 9636 2973 9639
rect 2372 9608 2973 9636
rect 2372 9596 2378 9608
rect 2961 9605 2973 9608
rect 3007 9605 3019 9639
rect 4356 9636 4384 9664
rect 7377 9639 7435 9645
rect 7377 9636 7389 9639
rect 4356 9608 7389 9636
rect 2961 9599 3019 9605
rect 7377 9605 7389 9608
rect 7423 9636 7435 9639
rect 7558 9636 7564 9648
rect 7423 9608 7564 9636
rect 7423 9605 7435 9608
rect 7377 9599 7435 9605
rect 7558 9596 7564 9608
rect 7616 9636 7622 9648
rect 7926 9636 7932 9648
rect 7616 9608 7932 9636
rect 7616 9596 7622 9608
rect 7926 9596 7932 9608
rect 7984 9596 7990 9648
rect 10612 9636 10640 9667
rect 11054 9664 11060 9676
rect 11112 9664 11118 9716
rect 11422 9704 11428 9716
rect 11383 9676 11428 9704
rect 11422 9664 11428 9676
rect 11480 9664 11486 9716
rect 11790 9704 11796 9716
rect 11751 9676 11796 9704
rect 11790 9664 11796 9676
rect 11848 9664 11854 9716
rect 12158 9704 12164 9716
rect 12119 9676 12164 9704
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 14185 9707 14243 9713
rect 14185 9704 14197 9707
rect 13872 9676 14197 9704
rect 13872 9664 13878 9676
rect 14185 9673 14197 9676
rect 14231 9673 14243 9707
rect 19150 9704 19156 9716
rect 19111 9676 19156 9704
rect 14185 9667 14243 9673
rect 19150 9664 19156 9676
rect 19208 9664 19214 9716
rect 20254 9704 20260 9716
rect 20215 9676 20260 9704
rect 20254 9664 20260 9676
rect 20312 9664 20318 9716
rect 21450 9704 21456 9716
rect 21411 9676 21456 9704
rect 21450 9664 21456 9676
rect 21508 9664 21514 9716
rect 21818 9704 21824 9716
rect 21779 9676 21824 9704
rect 21818 9664 21824 9676
rect 21876 9664 21882 9716
rect 12434 9636 12440 9648
rect 10612 9608 12440 9636
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9568 2467 9571
rect 3418 9568 3424 9580
rect 2455 9540 3424 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 6822 9568 6828 9580
rect 4120 9540 4200 9568
rect 6783 9540 6828 9568
rect 4120 9528 4126 9540
rect 4172 9500 4200 9540
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 9125 9571 9183 9577
rect 9125 9537 9137 9571
rect 9171 9568 9183 9571
rect 9398 9568 9404 9580
rect 9171 9540 9404 9568
rect 9171 9537 9183 9540
rect 9125 9531 9183 9537
rect 9398 9528 9404 9540
rect 9456 9528 9462 9580
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9568 10379 9571
rect 10778 9568 10784 9580
rect 10367 9540 10784 9568
rect 10367 9537 10379 9540
rect 10321 9531 10379 9537
rect 10778 9528 10784 9540
rect 10836 9568 10842 9580
rect 11164 9577 11192 9608
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 13906 9596 13912 9648
rect 13964 9636 13970 9648
rect 14461 9639 14519 9645
rect 14461 9636 14473 9639
rect 13964 9608 14473 9636
rect 13964 9596 13970 9608
rect 14461 9605 14473 9608
rect 14507 9636 14519 9639
rect 14553 9639 14611 9645
rect 14553 9636 14565 9639
rect 14507 9608 14565 9636
rect 14507 9605 14519 9608
rect 14461 9599 14519 9605
rect 14553 9605 14565 9608
rect 14599 9605 14611 9639
rect 14553 9599 14611 9605
rect 15838 9596 15844 9648
rect 15896 9636 15902 9648
rect 15896 9608 21220 9636
rect 15896 9596 15902 9608
rect 10928 9571 10986 9577
rect 10928 9568 10940 9571
rect 10836 9540 10940 9568
rect 10836 9528 10842 9540
rect 10928 9537 10940 9540
rect 10974 9537 10986 9571
rect 10928 9531 10986 9537
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9537 11207 9571
rect 17586 9568 17592 9580
rect 11149 9531 11207 9537
rect 13786 9540 17592 9568
rect 4614 9500 4620 9512
rect 4172 9472 4620 9500
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 13173 9503 13231 9509
rect 13173 9500 13185 9503
rect 13004 9472 13185 9500
rect 2501 9435 2559 9441
rect 2501 9401 2513 9435
rect 2547 9401 2559 9435
rect 2501 9395 2559 9401
rect 4938 9435 4996 9441
rect 4938 9401 4950 9435
rect 4984 9401 4996 9435
rect 8478 9432 8484 9444
rect 8439 9404 8484 9432
rect 4938 9395 4996 9401
rect 1857 9367 1915 9373
rect 1857 9333 1869 9367
rect 1903 9364 1915 9367
rect 2038 9364 2044 9376
rect 1903 9336 2044 9364
rect 1903 9333 1915 9336
rect 1857 9327 1915 9333
rect 2038 9324 2044 9336
rect 2096 9324 2102 9376
rect 2130 9324 2136 9376
rect 2188 9364 2194 9376
rect 2516 9364 2544 9395
rect 3418 9364 3424 9376
rect 2188 9336 2544 9364
rect 3379 9336 3424 9364
rect 2188 9324 2194 9336
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 4430 9364 4436 9376
rect 4391 9336 4436 9364
rect 4430 9324 4436 9336
rect 4488 9364 4494 9376
rect 4953 9364 4981 9395
rect 8478 9392 8484 9404
rect 8536 9392 8542 9444
rect 8570 9392 8576 9444
rect 8628 9432 8634 9444
rect 9953 9435 10011 9441
rect 8628 9404 8673 9432
rect 8628 9392 8634 9404
rect 9953 9401 9965 9435
rect 9999 9432 10011 9435
rect 10781 9435 10839 9441
rect 10781 9432 10793 9435
rect 9999 9404 10793 9432
rect 9999 9401 10011 9404
rect 9953 9395 10011 9401
rect 10781 9401 10793 9404
rect 10827 9432 10839 9435
rect 11238 9432 11244 9444
rect 10827 9404 11244 9432
rect 10827 9401 10839 9404
rect 10781 9395 10839 9401
rect 11238 9392 11244 9404
rect 11296 9392 11302 9444
rect 4488 9336 4981 9364
rect 4488 9324 4494 9336
rect 5258 9324 5264 9376
rect 5316 9364 5322 9376
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 5316 9336 5549 9364
rect 5316 9324 5322 9336
rect 5537 9333 5549 9336
rect 5583 9333 5595 9367
rect 7742 9364 7748 9376
rect 7703 9336 7748 9364
rect 5537 9327 5595 9333
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 8297 9367 8355 9373
rect 8297 9333 8309 9367
rect 8343 9364 8355 9367
rect 8588 9364 8616 9392
rect 8343 9336 8616 9364
rect 8343 9333 8355 9336
rect 8297 9327 8355 9333
rect 10502 9324 10508 9376
rect 10560 9364 10566 9376
rect 13004 9373 13032 9472
rect 13173 9469 13185 9472
rect 13219 9500 13231 9503
rect 13354 9500 13360 9512
rect 13219 9472 13360 9500
rect 13219 9469 13231 9472
rect 13173 9463 13231 9469
rect 13354 9460 13360 9472
rect 13412 9460 13418 9512
rect 13630 9500 13636 9512
rect 13591 9472 13636 9500
rect 13630 9460 13636 9472
rect 13688 9500 13694 9512
rect 13786 9500 13814 9540
rect 17586 9528 17592 9540
rect 17644 9528 17650 9580
rect 17862 9528 17868 9580
rect 17920 9568 17926 9580
rect 18230 9568 18236 9580
rect 17920 9540 18236 9568
rect 17920 9528 17926 9540
rect 18230 9528 18236 9540
rect 18288 9528 18294 9580
rect 20530 9568 20536 9580
rect 20491 9540 20536 9568
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 21192 9577 21220 9608
rect 21177 9571 21235 9577
rect 21177 9537 21189 9571
rect 21223 9568 21235 9571
rect 21542 9568 21548 9580
rect 21223 9540 21548 9568
rect 21223 9537 21235 9540
rect 21177 9531 21235 9537
rect 21542 9528 21548 9540
rect 21600 9528 21606 9580
rect 13688 9472 13814 9500
rect 13909 9503 13967 9509
rect 13688 9460 13694 9472
rect 13909 9469 13921 9503
rect 13955 9500 13967 9503
rect 14734 9500 14740 9512
rect 13955 9472 14740 9500
rect 13955 9469 13967 9472
rect 13909 9463 13967 9469
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 14461 9435 14519 9441
rect 14461 9401 14473 9435
rect 14507 9432 14519 9435
rect 14826 9432 14832 9444
rect 14507 9404 14832 9432
rect 14507 9401 14519 9404
rect 14461 9395 14519 9401
rect 14826 9392 14832 9404
rect 14884 9432 14890 9444
rect 15058 9435 15116 9441
rect 15058 9432 15070 9435
rect 14884 9404 15070 9432
rect 14884 9392 14890 9404
rect 15058 9401 15070 9404
rect 15104 9432 15116 9435
rect 17773 9435 17831 9441
rect 17773 9432 17785 9435
rect 15104 9404 17785 9432
rect 15104 9401 15116 9404
rect 15058 9395 15116 9401
rect 17773 9401 17785 9404
rect 17819 9432 17831 9435
rect 18554 9435 18612 9441
rect 18554 9432 18566 9435
rect 17819 9404 18566 9432
rect 17819 9401 17831 9404
rect 17773 9395 17831 9401
rect 18554 9401 18566 9404
rect 18600 9432 18612 9435
rect 18782 9432 18788 9444
rect 18600 9404 18788 9432
rect 18600 9401 18612 9404
rect 18554 9395 18612 9401
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 20625 9435 20683 9441
rect 20625 9401 20637 9435
rect 20671 9401 20683 9435
rect 20625 9395 20683 9401
rect 12989 9367 13047 9373
rect 12989 9364 13001 9367
rect 10560 9336 13001 9364
rect 10560 9324 10566 9336
rect 12989 9333 13001 9336
rect 13035 9333 13047 9367
rect 12989 9327 13047 9333
rect 15657 9367 15715 9373
rect 15657 9333 15669 9367
rect 15703 9364 15715 9367
rect 15930 9364 15936 9376
rect 15703 9336 15936 9364
rect 15703 9333 15715 9336
rect 15657 9327 15715 9333
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 16482 9364 16488 9376
rect 16443 9336 16488 9364
rect 16482 9324 16488 9336
rect 16540 9324 16546 9376
rect 17221 9367 17279 9373
rect 17221 9333 17233 9367
rect 17267 9364 17279 9367
rect 17494 9364 17500 9376
rect 17267 9336 17500 9364
rect 17267 9333 17279 9336
rect 17221 9327 17279 9333
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 20254 9324 20260 9376
rect 20312 9364 20318 9376
rect 20640 9364 20668 9395
rect 20312 9336 20668 9364
rect 20312 9324 20318 9336
rect 1104 9274 22816 9296
rect 1104 9222 8982 9274
rect 9034 9222 9046 9274
rect 9098 9222 9110 9274
rect 9162 9222 9174 9274
rect 9226 9222 16982 9274
rect 17034 9222 17046 9274
rect 17098 9222 17110 9274
rect 17162 9222 17174 9274
rect 17226 9222 22816 9274
rect 1104 9200 22816 9222
rect 106 9120 112 9172
rect 164 9160 170 9172
rect 4249 9163 4307 9169
rect 4249 9160 4261 9163
rect 164 9132 4261 9160
rect 164 9120 170 9132
rect 4249 9129 4261 9132
rect 4295 9129 4307 9163
rect 4614 9160 4620 9172
rect 4575 9132 4620 9160
rect 4249 9123 4307 9129
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 5258 9160 5264 9172
rect 5219 9132 5264 9160
rect 5258 9120 5264 9132
rect 5316 9120 5322 9172
rect 6914 9160 6920 9172
rect 5644 9132 6920 9160
rect 2038 9092 2044 9104
rect 1999 9064 2044 9092
rect 2038 9052 2044 9064
rect 2096 9052 2102 9104
rect 5644 9092 5672 9132
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 8205 9163 8263 9169
rect 8205 9129 8217 9163
rect 8251 9160 8263 9163
rect 8478 9160 8484 9172
rect 8251 9132 8484 9160
rect 8251 9129 8263 9132
rect 8205 9123 8263 9129
rect 8478 9120 8484 9132
rect 8536 9160 8542 9172
rect 8665 9163 8723 9169
rect 8665 9160 8677 9163
rect 8536 9132 8677 9160
rect 8536 9120 8542 9132
rect 8665 9129 8677 9132
rect 8711 9129 8723 9163
rect 8665 9123 8723 9129
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 12023 9163 12081 9169
rect 12023 9160 12035 9163
rect 10928 9132 12035 9160
rect 10928 9120 10934 9132
rect 12023 9129 12035 9132
rect 12069 9129 12081 9163
rect 12023 9123 12081 9129
rect 14277 9163 14335 9169
rect 14277 9129 14289 9163
rect 14323 9160 14335 9163
rect 14458 9160 14464 9172
rect 14323 9132 14464 9160
rect 14323 9129 14335 9132
rect 14277 9123 14335 9129
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 14734 9160 14740 9172
rect 14695 9132 14740 9160
rect 14734 9120 14740 9132
rect 14792 9120 14798 9172
rect 15654 9160 15660 9172
rect 15567 9132 15660 9160
rect 15654 9120 15660 9132
rect 15712 9160 15718 9172
rect 16482 9160 16488 9172
rect 15712 9132 16488 9160
rect 15712 9120 15718 9132
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 17221 9163 17279 9169
rect 17221 9129 17233 9163
rect 17267 9160 17279 9163
rect 17586 9160 17592 9172
rect 17267 9132 17592 9160
rect 17267 9129 17279 9132
rect 17221 9123 17279 9129
rect 17586 9120 17592 9132
rect 17644 9120 17650 9172
rect 18230 9160 18236 9172
rect 18191 9132 18236 9160
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 20530 9160 20536 9172
rect 20491 9132 20536 9160
rect 20530 9120 20536 9132
rect 20588 9120 20594 9172
rect 4080 9064 5672 9092
rect 5721 9095 5779 9101
rect 3878 8984 3884 9036
rect 3936 9024 3942 9036
rect 4080 9033 4108 9064
rect 5721 9061 5733 9095
rect 5767 9092 5779 9095
rect 6086 9092 6092 9104
rect 5767 9064 6092 9092
rect 5767 9061 5779 9064
rect 5721 9055 5779 9061
rect 6086 9052 6092 9064
rect 6144 9052 6150 9104
rect 13354 9092 13360 9104
rect 13315 9064 13360 9092
rect 13354 9052 13360 9064
rect 13412 9052 13418 9104
rect 15930 9092 15936 9104
rect 15843 9064 15936 9092
rect 15930 9052 15936 9064
rect 15988 9092 15994 9104
rect 16574 9092 16580 9104
rect 15988 9064 16580 9092
rect 15988 9052 15994 9064
rect 16574 9052 16580 9064
rect 16632 9052 16638 9104
rect 4053 9027 4111 9033
rect 4053 9024 4065 9027
rect 3936 8996 4065 9024
rect 3936 8984 3942 8996
rect 4053 8993 4065 8996
rect 4099 8993 4111 9027
rect 4053 8987 4111 8993
rect 7926 8984 7932 9036
rect 7984 9024 7990 9036
rect 9674 9024 9680 9036
rect 7984 8996 9680 9024
rect 7984 8984 7990 8996
rect 9674 8984 9680 8996
rect 9732 9024 9738 9036
rect 10594 9024 10600 9036
rect 9732 8996 10600 9024
rect 9732 8984 9738 8996
rect 10594 8984 10600 8996
rect 10652 9024 10658 9036
rect 10965 9027 11023 9033
rect 10965 9024 10977 9027
rect 10652 8996 10977 9024
rect 10652 8984 10658 8996
rect 10965 8993 10977 8996
rect 11011 9024 11023 9027
rect 11885 9027 11943 9033
rect 11011 8996 11284 9024
rect 11011 8993 11023 8996
rect 10965 8987 11023 8993
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8956 2007 8959
rect 5626 8956 5632 8968
rect 1995 8928 2912 8956
rect 5539 8928 5632 8956
rect 1995 8925 2007 8928
rect 1949 8919 2007 8925
rect 2884 8900 2912 8928
rect 5626 8916 5632 8928
rect 5684 8956 5690 8968
rect 7101 8959 7159 8965
rect 7101 8956 7113 8959
rect 5684 8928 7113 8956
rect 5684 8916 5690 8928
rect 7101 8925 7113 8928
rect 7147 8925 7159 8959
rect 7101 8919 7159 8925
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 10502 8956 10508 8968
rect 10367 8928 10508 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 10502 8916 10508 8928
rect 10560 8916 10566 8968
rect 2314 8848 2320 8900
rect 2372 8888 2378 8900
rect 2501 8891 2559 8897
rect 2501 8888 2513 8891
rect 2372 8860 2513 8888
rect 2372 8848 2378 8860
rect 2501 8857 2513 8860
rect 2547 8857 2559 8891
rect 2501 8851 2559 8857
rect 2866 8848 2872 8900
rect 2924 8888 2930 8900
rect 5718 8888 5724 8900
rect 2924 8860 5724 8888
rect 2924 8848 2930 8860
rect 5718 8848 5724 8860
rect 5776 8848 5782 8900
rect 5902 8848 5908 8900
rect 5960 8888 5966 8900
rect 6181 8891 6239 8897
rect 6181 8888 6193 8891
rect 5960 8860 6193 8888
rect 5960 8848 5966 8860
rect 6181 8857 6193 8860
rect 6227 8857 6239 8891
rect 11256 8888 11284 8996
rect 11885 8993 11897 9027
rect 11931 9024 11943 9027
rect 11974 9024 11980 9036
rect 11931 8996 11980 9024
rect 11931 8993 11943 8996
rect 11885 8987 11943 8993
rect 11974 8984 11980 8996
rect 12032 8984 12038 9036
rect 20968 9027 21026 9033
rect 20968 8993 20980 9027
rect 21014 9024 21026 9027
rect 21450 9024 21456 9036
rect 21014 8996 21456 9024
rect 21014 8993 21026 8996
rect 20968 8987 21026 8993
rect 21450 8984 21456 8996
rect 21508 8984 21514 9036
rect 13262 8956 13268 8968
rect 13223 8928 13268 8956
rect 13262 8916 13268 8928
rect 13320 8956 13326 8968
rect 14550 8956 14556 8968
rect 13320 8928 14556 8956
rect 13320 8916 13326 8928
rect 14550 8916 14556 8928
rect 14608 8916 14614 8968
rect 15838 8956 15844 8968
rect 15799 8928 15844 8956
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 16206 8956 16212 8968
rect 16167 8928 16212 8956
rect 16206 8916 16212 8928
rect 16264 8916 16270 8968
rect 13538 8888 13544 8900
rect 11256 8860 13544 8888
rect 6181 8851 6239 8857
rect 13538 8848 13544 8860
rect 13596 8848 13602 8900
rect 13814 8848 13820 8900
rect 13872 8888 13878 8900
rect 13872 8860 13917 8888
rect 13872 8848 13878 8860
rect 17218 8848 17224 8900
rect 17276 8888 17282 8900
rect 21039 8891 21097 8897
rect 21039 8888 21051 8891
rect 17276 8860 21051 8888
rect 17276 8848 17282 8860
rect 21039 8857 21051 8860
rect 21085 8857 21097 8891
rect 21039 8851 21097 8857
rect 1394 8780 1400 8832
rect 1452 8820 1458 8832
rect 1673 8823 1731 8829
rect 1673 8820 1685 8823
rect 1452 8792 1685 8820
rect 1452 8780 1458 8792
rect 1673 8789 1685 8792
rect 1719 8820 1731 8823
rect 6638 8820 6644 8832
rect 1719 8792 6644 8820
rect 1719 8789 1731 8792
rect 1673 8783 1731 8789
rect 6638 8780 6644 8792
rect 6696 8780 6702 8832
rect 7834 8820 7840 8832
rect 7795 8792 7840 8820
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 1104 8730 22816 8752
rect 1104 8678 4982 8730
rect 5034 8678 5046 8730
rect 5098 8678 5110 8730
rect 5162 8678 5174 8730
rect 5226 8678 12982 8730
rect 13034 8678 13046 8730
rect 13098 8678 13110 8730
rect 13162 8678 13174 8730
rect 13226 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 22816 8730
rect 1104 8656 22816 8678
rect 2409 8619 2467 8625
rect 2409 8585 2421 8619
rect 2455 8616 2467 8619
rect 2866 8616 2872 8628
rect 2455 8588 2872 8616
rect 2455 8585 2467 8588
rect 2409 8579 2467 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 4157 8619 4215 8625
rect 4157 8616 4169 8619
rect 2976 8588 4169 8616
rect 2038 8548 2044 8560
rect 1951 8520 2044 8548
rect 2038 8508 2044 8520
rect 2096 8548 2102 8560
rect 2976 8548 3004 8588
rect 4157 8585 4169 8588
rect 4203 8585 4215 8619
rect 4157 8579 4215 8585
rect 5077 8619 5135 8625
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 5626 8616 5632 8628
rect 5123 8588 5632 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 10594 8616 10600 8628
rect 10555 8588 10600 8616
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 14550 8616 14556 8628
rect 14511 8588 14556 8616
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 15378 8616 15384 8628
rect 15339 8588 15384 8616
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 16574 8616 16580 8628
rect 16535 8588 16580 8616
rect 16574 8576 16580 8588
rect 16632 8576 16638 8628
rect 21450 8616 21456 8628
rect 21411 8588 21456 8616
rect 21450 8576 21456 8588
rect 21508 8576 21514 8628
rect 21821 8619 21879 8625
rect 21821 8585 21833 8619
rect 21867 8616 21879 8619
rect 22186 8616 22192 8628
rect 21867 8588 22192 8616
rect 21867 8585 21879 8588
rect 21821 8579 21879 8585
rect 2096 8520 3004 8548
rect 2096 8508 2102 8520
rect 3142 8508 3148 8560
rect 3200 8548 3206 8560
rect 4617 8551 4675 8557
rect 4617 8548 4629 8551
rect 3200 8520 4629 8548
rect 3200 8508 3206 8520
rect 4617 8517 4629 8520
rect 4663 8548 4675 8551
rect 4663 8520 5304 8548
rect 4663 8517 4675 8520
rect 4617 8511 4675 8517
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8480 3295 8483
rect 3602 8480 3608 8492
rect 3283 8452 3608 8480
rect 3283 8449 3295 8452
rect 3237 8443 3295 8449
rect 3602 8440 3608 8452
rect 3660 8440 3666 8492
rect 5276 8489 5304 8520
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 9398 8548 9404 8560
rect 8352 8520 9404 8548
rect 8352 8508 8358 8520
rect 9398 8508 9404 8520
rect 9456 8548 9462 8560
rect 10137 8551 10195 8557
rect 10137 8548 10149 8551
rect 9456 8520 10149 8548
rect 9456 8508 9462 8520
rect 10137 8517 10149 8520
rect 10183 8517 10195 8551
rect 11974 8548 11980 8560
rect 11887 8520 11980 8548
rect 10137 8511 10195 8517
rect 11974 8508 11980 8520
rect 12032 8548 12038 8560
rect 13814 8548 13820 8560
rect 12032 8520 13820 8548
rect 12032 8508 12038 8520
rect 13786 8508 13820 8520
rect 13872 8508 13878 8560
rect 16206 8548 16212 8560
rect 16167 8520 16212 8548
rect 16206 8508 16212 8520
rect 16264 8508 16270 8560
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8449 5319 8483
rect 5261 8443 5319 8449
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8480 9091 8483
rect 9585 8483 9643 8489
rect 9585 8480 9597 8483
rect 9079 8452 9597 8480
rect 9079 8449 9091 8452
rect 9033 8443 9091 8449
rect 9585 8449 9597 8452
rect 9631 8480 9643 8483
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 9631 8452 11069 8480
rect 9631 8449 9643 8452
rect 9585 8443 9643 8449
rect 11057 8449 11069 8452
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8480 12587 8483
rect 13262 8480 13268 8492
rect 12575 8452 13268 8480
rect 12575 8449 12587 8452
rect 12529 8443 12587 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 13446 8440 13452 8492
rect 13504 8480 13510 8492
rect 13633 8483 13691 8489
rect 13633 8480 13645 8483
rect 13504 8452 13645 8480
rect 13504 8440 13510 8452
rect 13633 8449 13645 8452
rect 13679 8449 13691 8483
rect 13786 8480 13814 8508
rect 13909 8483 13967 8489
rect 13909 8480 13921 8483
rect 13786 8452 13921 8480
rect 13633 8443 13691 8449
rect 13909 8449 13921 8452
rect 13955 8449 13967 8483
rect 15654 8480 15660 8492
rect 15615 8452 15660 8480
rect 13909 8443 13967 8449
rect 15654 8440 15660 8452
rect 15712 8440 15718 8492
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8412 7803 8415
rect 7834 8412 7840 8424
rect 7791 8384 7840 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 7834 8372 7840 8384
rect 7892 8372 7898 8424
rect 20968 8415 21026 8421
rect 20968 8381 20980 8415
rect 21014 8412 21026 8415
rect 21836 8412 21864 8579
rect 22186 8576 22192 8588
rect 22244 8576 22250 8628
rect 21014 8384 21864 8412
rect 21014 8381 21026 8384
rect 20968 8375 21026 8381
rect 3558 8347 3616 8353
rect 3558 8313 3570 8347
rect 3604 8344 3616 8347
rect 4430 8344 4436 8356
rect 3604 8316 4436 8344
rect 3604 8313 3616 8316
rect 3558 8307 3616 8313
rect 106 8236 112 8288
rect 164 8276 170 8288
rect 1581 8279 1639 8285
rect 1581 8276 1593 8279
rect 164 8248 1593 8276
rect 164 8236 170 8248
rect 1581 8245 1593 8248
rect 1627 8245 1639 8279
rect 3050 8276 3056 8288
rect 3011 8248 3056 8276
rect 1581 8239 1639 8245
rect 3050 8236 3056 8248
rect 3108 8276 3114 8288
rect 3573 8276 3601 8307
rect 4430 8304 4436 8316
rect 4488 8304 4494 8356
rect 5350 8344 5356 8356
rect 5311 8316 5356 8344
rect 5350 8304 5356 8316
rect 5408 8304 5414 8356
rect 5902 8344 5908 8356
rect 5863 8316 5908 8344
rect 5902 8304 5908 8316
rect 5960 8304 5966 8356
rect 7561 8347 7619 8353
rect 7561 8344 7573 8347
rect 6058 8316 7573 8344
rect 3108 8248 3601 8276
rect 4448 8276 4476 8304
rect 6058 8276 6086 8316
rect 7561 8313 7573 8316
rect 7607 8344 7619 8347
rect 8018 8344 8024 8356
rect 7607 8316 8024 8344
rect 7607 8313 7619 8316
rect 7561 8307 7619 8313
rect 8018 8304 8024 8316
rect 8076 8353 8082 8356
rect 8076 8347 8124 8353
rect 8076 8313 8078 8347
rect 8112 8313 8124 8347
rect 8076 8307 8124 8313
rect 8076 8304 8082 8307
rect 9674 8304 9680 8356
rect 9732 8344 9738 8356
rect 9732 8316 9777 8344
rect 9732 8304 9738 8316
rect 13722 8304 13728 8356
rect 13780 8344 13786 8356
rect 15749 8347 15807 8353
rect 13780 8316 13825 8344
rect 13780 8304 13786 8316
rect 15749 8313 15761 8347
rect 15795 8313 15807 8347
rect 15749 8307 15807 8313
rect 6178 8276 6184 8288
rect 4448 8248 6086 8276
rect 6139 8248 6184 8276
rect 3108 8236 3114 8248
rect 6178 8236 6184 8248
rect 6236 8236 6242 8288
rect 8662 8276 8668 8288
rect 8623 8248 8668 8276
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 9401 8279 9459 8285
rect 9401 8245 9413 8279
rect 9447 8276 9459 8279
rect 9692 8276 9720 8304
rect 9447 8248 9720 8276
rect 13265 8279 13323 8285
rect 9447 8245 9459 8248
rect 9401 8239 9459 8245
rect 13265 8245 13277 8279
rect 13311 8276 13323 8279
rect 13354 8276 13360 8288
rect 13311 8248 13360 8276
rect 13311 8245 13323 8248
rect 13265 8239 13323 8245
rect 13354 8236 13360 8248
rect 13412 8236 13418 8288
rect 15010 8276 15016 8288
rect 14971 8248 15016 8276
rect 15010 8236 15016 8248
rect 15068 8236 15074 8288
rect 15378 8236 15384 8288
rect 15436 8276 15442 8288
rect 15764 8276 15792 8307
rect 15436 8248 15792 8276
rect 15436 8236 15442 8248
rect 16298 8236 16304 8288
rect 16356 8276 16362 8288
rect 21039 8279 21097 8285
rect 21039 8276 21051 8279
rect 16356 8248 21051 8276
rect 16356 8236 16362 8248
rect 21039 8245 21051 8248
rect 21085 8245 21097 8279
rect 21039 8239 21097 8245
rect 1104 8186 22816 8208
rect 1104 8134 8982 8186
rect 9034 8134 9046 8186
rect 9098 8134 9110 8186
rect 9162 8134 9174 8186
rect 9226 8134 16982 8186
rect 17034 8134 17046 8186
rect 17098 8134 17110 8186
rect 17162 8134 17174 8186
rect 17226 8134 22816 8186
rect 1104 8112 22816 8134
rect 3878 8072 3884 8084
rect 3839 8044 3884 8072
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 7834 8072 7840 8084
rect 7795 8044 7840 8072
rect 7834 8032 7840 8044
rect 7892 8032 7898 8084
rect 13446 8032 13452 8084
rect 13504 8072 13510 8084
rect 15010 8072 15016 8084
rect 13504 8044 15016 8072
rect 13504 8032 13510 8044
rect 15010 8032 15016 8044
rect 15068 8032 15074 8084
rect 15838 8072 15844 8084
rect 15799 8044 15844 8072
rect 15838 8032 15844 8044
rect 15896 8032 15902 8084
rect 17402 8032 17408 8084
rect 17460 8072 17466 8084
rect 21039 8075 21097 8081
rect 21039 8072 21051 8075
rect 17460 8044 21051 8072
rect 17460 8032 17466 8044
rect 21039 8041 21051 8044
rect 21085 8041 21097 8075
rect 21039 8035 21097 8041
rect 2317 8007 2375 8013
rect 2317 7973 2329 8007
rect 2363 8004 2375 8007
rect 2406 8004 2412 8016
rect 2363 7976 2412 8004
rect 2363 7973 2375 7976
rect 2317 7967 2375 7973
rect 2406 7964 2412 7976
rect 2464 7964 2470 8016
rect 5905 8007 5963 8013
rect 5905 7973 5917 8007
rect 5951 8004 5963 8007
rect 6178 8004 6184 8016
rect 5951 7976 6184 8004
rect 5951 7973 5963 7976
rect 5905 7967 5963 7973
rect 6178 7964 6184 7976
rect 6236 7964 6242 8016
rect 9674 8004 9680 8016
rect 9635 7976 9680 8004
rect 9674 7964 9680 7976
rect 9732 7964 9738 8016
rect 12618 7964 12624 8016
rect 12676 8004 12682 8016
rect 12850 8007 12908 8013
rect 12850 8004 12862 8007
rect 12676 7976 12862 8004
rect 12676 7964 12682 7976
rect 12850 7973 12862 7976
rect 12896 7973 12908 8007
rect 12850 7967 12908 7973
rect 4111 7939 4169 7945
rect 4111 7905 4123 7939
rect 4157 7905 4169 7939
rect 4111 7899 4169 7905
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7936 5135 7939
rect 5350 7936 5356 7948
rect 5123 7908 5356 7936
rect 5123 7905 5135 7908
rect 5077 7899 5135 7905
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7868 2283 7871
rect 2314 7868 2320 7880
rect 2271 7840 2320 7868
rect 2271 7837 2283 7840
rect 2225 7831 2283 7837
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 2498 7868 2504 7880
rect 2459 7840 2504 7868
rect 2498 7828 2504 7840
rect 2556 7868 2562 7880
rect 4126 7868 4154 7899
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 7193 7939 7251 7945
rect 7193 7905 7205 7939
rect 7239 7905 7251 7939
rect 7193 7899 7251 7905
rect 4525 7871 4583 7877
rect 4525 7868 4537 7871
rect 2556 7840 4537 7868
rect 2556 7828 2562 7840
rect 4525 7837 4537 7840
rect 4571 7837 4583 7871
rect 7208 7868 7236 7899
rect 7282 7896 7288 7948
rect 7340 7936 7346 7948
rect 7377 7939 7435 7945
rect 7377 7936 7389 7939
rect 7340 7908 7389 7936
rect 7340 7896 7346 7908
rect 7377 7905 7389 7908
rect 7423 7905 7435 7939
rect 7377 7899 7435 7905
rect 7558 7896 7564 7948
rect 7616 7936 7622 7948
rect 7745 7939 7803 7945
rect 7745 7936 7757 7939
rect 7616 7908 7757 7936
rect 7616 7896 7622 7908
rect 7745 7905 7757 7908
rect 7791 7905 7803 7939
rect 9766 7936 9772 7948
rect 9727 7908 9772 7936
rect 7745 7899 7803 7905
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 15378 7945 15384 7948
rect 15356 7939 15384 7945
rect 15356 7936 15368 7939
rect 15291 7908 15368 7936
rect 15356 7905 15368 7908
rect 15436 7936 15442 7948
rect 16206 7936 16212 7948
rect 15436 7908 16212 7936
rect 15356 7899 15384 7905
rect 15378 7896 15384 7899
rect 15436 7896 15442 7908
rect 16206 7896 16212 7908
rect 16264 7896 16270 7948
rect 20968 7939 21026 7945
rect 20968 7905 20980 7939
rect 21014 7936 21026 7939
rect 21358 7936 21364 7948
rect 21014 7908 21364 7936
rect 21014 7905 21026 7908
rect 20968 7899 21026 7905
rect 21358 7896 21364 7908
rect 21416 7896 21422 7948
rect 7466 7868 7472 7880
rect 7208 7840 7472 7868
rect 4525 7831 4583 7837
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 12529 7871 12587 7877
rect 12529 7837 12541 7871
rect 12575 7868 12587 7871
rect 12802 7868 12808 7880
rect 12575 7840 12808 7868
rect 12575 7837 12587 7840
rect 12529 7831 12587 7837
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 14369 7803 14427 7809
rect 14369 7800 14381 7803
rect 13924 7772 14381 7800
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 1946 7732 1952 7744
rect 1907 7704 1952 7732
rect 1946 7692 1952 7704
rect 2004 7692 2010 7744
rect 3329 7735 3387 7741
rect 3329 7701 3341 7735
rect 3375 7732 3387 7735
rect 3602 7732 3608 7744
rect 3375 7704 3608 7732
rect 3375 7701 3387 7704
rect 3329 7695 3387 7701
rect 3602 7692 3608 7704
rect 3660 7692 3666 7744
rect 3694 7692 3700 7744
rect 3752 7732 3758 7744
rect 4203 7735 4261 7741
rect 4203 7732 4215 7735
rect 3752 7704 4215 7732
rect 3752 7692 3758 7704
rect 4203 7701 4215 7704
rect 4249 7701 4261 7735
rect 8846 7732 8852 7744
rect 8807 7704 8852 7732
rect 4203 7695 4261 7701
rect 8846 7692 8852 7704
rect 8904 7692 8910 7744
rect 10778 7732 10784 7744
rect 10739 7704 10784 7732
rect 10778 7692 10784 7704
rect 10836 7692 10842 7744
rect 13449 7735 13507 7741
rect 13449 7701 13461 7735
rect 13495 7732 13507 7735
rect 13630 7732 13636 7744
rect 13495 7704 13636 7732
rect 13495 7701 13507 7704
rect 13449 7695 13507 7701
rect 13630 7692 13636 7704
rect 13688 7732 13694 7744
rect 13924 7732 13952 7772
rect 14369 7769 14381 7772
rect 14415 7769 14427 7803
rect 14369 7763 14427 7769
rect 14090 7732 14096 7744
rect 13688 7704 13952 7732
rect 14051 7704 14096 7732
rect 13688 7692 13694 7704
rect 14090 7692 14096 7704
rect 14148 7692 14154 7744
rect 15427 7735 15485 7741
rect 15427 7701 15439 7735
rect 15473 7732 15485 7735
rect 15562 7732 15568 7744
rect 15473 7704 15568 7732
rect 15473 7701 15485 7704
rect 15427 7695 15485 7701
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 1104 7642 22816 7664
rect 1104 7590 4982 7642
rect 5034 7590 5046 7642
rect 5098 7590 5110 7642
rect 5162 7590 5174 7642
rect 5226 7590 12982 7642
rect 13034 7590 13046 7642
rect 13098 7590 13110 7642
rect 13162 7590 13174 7642
rect 13226 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 22816 7642
rect 1104 7568 22816 7590
rect 2406 7488 2412 7540
rect 2464 7528 2470 7540
rect 2685 7531 2743 7537
rect 2685 7528 2697 7531
rect 2464 7500 2697 7528
rect 2464 7488 2470 7500
rect 2685 7497 2697 7500
rect 2731 7528 2743 7531
rect 4065 7531 4123 7537
rect 4065 7528 4077 7531
rect 2731 7500 4077 7528
rect 2731 7497 2743 7500
rect 2685 7491 2743 7497
rect 4065 7497 4077 7500
rect 4111 7497 4123 7531
rect 4065 7491 4123 7497
rect 5334 7531 5392 7537
rect 5334 7497 5346 7531
rect 5380 7528 5392 7531
rect 5718 7528 5724 7540
rect 5380 7500 5724 7528
rect 5380 7497 5392 7500
rect 5334 7491 5392 7497
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 8021 7531 8079 7537
rect 8021 7528 8033 7531
rect 7340 7500 8033 7528
rect 7340 7488 7346 7500
rect 8021 7497 8033 7500
rect 8067 7497 8079 7531
rect 8662 7528 8668 7540
rect 8575 7500 8668 7528
rect 8021 7491 8079 7497
rect 8662 7488 8668 7500
rect 8720 7528 8726 7540
rect 8938 7528 8944 7540
rect 8720 7500 8944 7528
rect 8720 7488 8726 7500
rect 8938 7488 8944 7500
rect 8996 7528 9002 7540
rect 9766 7528 9772 7540
rect 8996 7500 9772 7528
rect 8996 7488 9002 7500
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 10962 7488 10968 7540
rect 11020 7528 11026 7540
rect 15378 7528 15384 7540
rect 11020 7500 11192 7528
rect 15339 7500 15384 7528
rect 11020 7488 11026 7500
rect 5442 7460 5448 7472
rect 5403 7432 5448 7460
rect 5442 7420 5448 7432
rect 5500 7420 5506 7472
rect 5997 7463 6055 7469
rect 5997 7429 6009 7463
rect 6043 7460 6055 7463
rect 7742 7460 7748 7472
rect 6043 7432 7748 7460
rect 6043 7429 6055 7432
rect 5997 7423 6055 7429
rect 7742 7420 7748 7432
rect 7800 7420 7806 7472
rect 9398 7460 9404 7472
rect 9359 7432 9404 7460
rect 9398 7420 9404 7432
rect 9456 7420 9462 7472
rect 10594 7420 10600 7472
rect 10652 7460 10658 7472
rect 11057 7463 11115 7469
rect 11057 7460 11069 7463
rect 10652 7432 11069 7460
rect 10652 7420 10658 7432
rect 11057 7429 11069 7432
rect 11103 7429 11115 7463
rect 11057 7423 11115 7429
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7392 2375 7395
rect 2498 7392 2504 7404
rect 2363 7364 2504 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7392 4951 7395
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 4939 7364 5549 7392
rect 4939 7361 4951 7364
rect 4893 7355 4951 7361
rect 5537 7361 5549 7364
rect 5583 7392 5595 7395
rect 6270 7392 6276 7404
rect 5583 7364 6276 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 6270 7352 6276 7364
rect 6328 7352 6334 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 7558 7392 7564 7404
rect 7423 7364 7564 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 8662 7352 8668 7404
rect 8720 7392 8726 7404
rect 10778 7392 10784 7404
rect 8720 7364 10784 7392
rect 8720 7352 8726 7364
rect 10778 7352 10784 7364
rect 10836 7392 10842 7404
rect 11164 7401 11192 7500
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 21177 7531 21235 7537
rect 21177 7497 21189 7531
rect 21223 7528 21235 7531
rect 21358 7528 21364 7540
rect 21223 7500 21364 7528
rect 21223 7497 21235 7500
rect 21177 7491 21235 7497
rect 21358 7488 21364 7500
rect 21416 7488 21422 7540
rect 10928 7395 10986 7401
rect 10928 7392 10940 7395
rect 10836 7364 10940 7392
rect 10836 7352 10842 7364
rect 10928 7361 10940 7364
rect 10974 7361 10986 7395
rect 10928 7355 10986 7361
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7361 11207 7395
rect 11149 7355 11207 7361
rect 11517 7395 11575 7401
rect 11517 7361 11529 7395
rect 11563 7392 11575 7395
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11563 7364 11897 7392
rect 11563 7361 11575 7364
rect 11517 7355 11575 7361
rect 11885 7361 11897 7364
rect 11931 7392 11943 7395
rect 17954 7392 17960 7404
rect 11931 7364 17960 7392
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 3142 7324 3148 7336
rect 3103 7296 3148 7324
rect 3142 7284 3148 7296
rect 3200 7284 3206 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 3252 7296 6837 7324
rect 1670 7256 1676 7268
rect 1583 7228 1676 7256
rect 1670 7216 1676 7228
rect 1728 7216 1734 7268
rect 1762 7216 1768 7268
rect 1820 7256 1826 7268
rect 3252 7256 3280 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 12434 7324 12440 7336
rect 12395 7296 12440 7324
rect 6825 7287 6883 7293
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 13004 7333 13032 7364
rect 17954 7352 17960 7364
rect 18012 7392 18018 7404
rect 18012 7364 18552 7392
rect 18012 7352 18018 7364
rect 12989 7327 13047 7333
rect 12989 7293 13001 7327
rect 13035 7293 13047 7327
rect 12989 7287 13047 7293
rect 14001 7327 14059 7333
rect 14001 7293 14013 7327
rect 14047 7293 14059 7327
rect 14001 7287 14059 7293
rect 1820 7228 1865 7256
rect 1964 7228 3280 7256
rect 3466 7259 3524 7265
rect 1820 7216 1826 7228
rect 1688 7188 1716 7216
rect 1964 7188 1992 7228
rect 3466 7225 3478 7259
rect 3512 7225 3524 7259
rect 3466 7219 3524 7225
rect 4617 7259 4675 7265
rect 4617 7225 4629 7259
rect 4663 7256 4675 7259
rect 5169 7259 5227 7265
rect 5169 7256 5181 7259
rect 4663 7228 5181 7256
rect 4663 7225 4675 7228
rect 4617 7219 4675 7225
rect 5169 7225 5181 7228
rect 5215 7256 5227 7259
rect 5997 7259 6055 7265
rect 5997 7256 6009 7259
rect 5215 7228 6009 7256
rect 5215 7225 5227 7228
rect 5169 7219 5227 7225
rect 5997 7225 6009 7228
rect 6043 7225 6055 7259
rect 5997 7219 6055 7225
rect 6273 7259 6331 7265
rect 6273 7225 6285 7259
rect 6319 7256 6331 7259
rect 8846 7256 8852 7268
rect 6319 7228 7512 7256
rect 8807 7228 8852 7256
rect 6319 7225 6331 7228
rect 6273 7219 6331 7225
rect 3050 7188 3056 7200
rect 1688 7160 1992 7188
rect 3011 7160 3056 7188
rect 3050 7148 3056 7160
rect 3108 7188 3114 7200
rect 3481 7188 3509 7219
rect 7484 7200 7512 7228
rect 8846 7216 8852 7228
rect 8904 7216 8910 7268
rect 8938 7216 8944 7268
rect 8996 7256 9002 7268
rect 10321 7259 10379 7265
rect 8996 7228 9041 7256
rect 8996 7216 9002 7228
rect 10321 7225 10333 7259
rect 10367 7256 10379 7259
rect 10781 7259 10839 7265
rect 10781 7256 10793 7259
rect 10367 7228 10793 7256
rect 10367 7225 10379 7228
rect 10321 7219 10379 7225
rect 10781 7225 10793 7228
rect 10827 7256 10839 7259
rect 11238 7256 11244 7268
rect 10827 7228 11244 7256
rect 10827 7225 10839 7228
rect 10781 7219 10839 7225
rect 3108 7160 3509 7188
rect 3108 7148 3114 7160
rect 4706 7148 4712 7200
rect 4764 7188 4770 7200
rect 4893 7191 4951 7197
rect 4893 7188 4905 7191
rect 4764 7160 4905 7188
rect 4764 7148 4770 7160
rect 4893 7157 4905 7160
rect 4939 7188 4951 7191
rect 4985 7191 5043 7197
rect 4985 7188 4997 7191
rect 4939 7160 4997 7188
rect 4939 7157 4951 7160
rect 4893 7151 4951 7157
rect 4985 7157 4997 7160
rect 5031 7157 5043 7191
rect 4985 7151 5043 7157
rect 5074 7148 5080 7200
rect 5132 7188 5138 7200
rect 5813 7191 5871 7197
rect 5813 7188 5825 7191
rect 5132 7160 5825 7188
rect 5132 7148 5138 7160
rect 5813 7157 5825 7160
rect 5859 7157 5871 7191
rect 6638 7188 6644 7200
rect 6599 7160 6644 7188
rect 5813 7151 5871 7157
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 7466 7148 7472 7200
rect 7524 7188 7530 7200
rect 7745 7191 7803 7197
rect 7745 7188 7757 7191
rect 7524 7160 7757 7188
rect 7524 7148 7530 7160
rect 7745 7157 7757 7160
rect 7791 7188 7803 7191
rect 10336 7188 10364 7219
rect 11238 7216 11244 7228
rect 11296 7216 11302 7268
rect 13538 7216 13544 7268
rect 13596 7256 13602 7268
rect 14016 7256 14044 7287
rect 14090 7284 14096 7336
rect 14148 7324 14154 7336
rect 18524 7333 18552 7364
rect 14461 7327 14519 7333
rect 14461 7324 14473 7327
rect 14148 7296 14473 7324
rect 14148 7284 14154 7296
rect 14461 7293 14473 7296
rect 14507 7293 14519 7327
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 14461 7287 14519 7293
rect 17788 7296 18061 7324
rect 14734 7256 14740 7268
rect 13596 7228 14044 7256
rect 14695 7228 14740 7256
rect 13596 7216 13602 7228
rect 10594 7188 10600 7200
rect 7791 7160 10364 7188
rect 10555 7160 10600 7188
rect 7791 7157 7803 7160
rect 7745 7151 7803 7157
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 12253 7191 12311 7197
rect 12253 7157 12265 7191
rect 12299 7188 12311 7191
rect 12618 7188 12624 7200
rect 12299 7160 12624 7188
rect 12299 7157 12311 7160
rect 12253 7151 12311 7157
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 12713 7191 12771 7197
rect 12713 7157 12725 7191
rect 12759 7188 12771 7191
rect 12802 7188 12808 7200
rect 12759 7160 12808 7188
rect 12759 7157 12771 7160
rect 12713 7151 12771 7157
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 13909 7191 13967 7197
rect 13909 7157 13921 7191
rect 13955 7188 13967 7191
rect 14016 7188 14044 7228
rect 14734 7216 14740 7228
rect 14792 7216 14798 7268
rect 17494 7188 17500 7200
rect 13955 7160 17500 7188
rect 13955 7157 13967 7160
rect 13909 7151 13967 7157
rect 17494 7148 17500 7160
rect 17552 7188 17558 7200
rect 17788 7197 17816 7296
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 18509 7327 18567 7333
rect 18509 7293 18521 7327
rect 18555 7293 18567 7327
rect 18509 7287 18567 7293
rect 19334 7284 19340 7336
rect 19392 7324 19398 7336
rect 19981 7327 20039 7333
rect 19981 7324 19993 7327
rect 19392 7296 19993 7324
rect 19392 7284 19398 7296
rect 19981 7293 19993 7296
rect 20027 7324 20039 7327
rect 20717 7327 20775 7333
rect 20717 7324 20729 7327
rect 20027 7296 20729 7324
rect 20027 7293 20039 7296
rect 19981 7287 20039 7293
rect 20717 7293 20729 7296
rect 20763 7324 20775 7327
rect 21266 7324 21272 7336
rect 20763 7296 21272 7324
rect 20763 7293 20775 7296
rect 20717 7287 20775 7293
rect 21266 7284 21272 7296
rect 21324 7284 21330 7336
rect 17773 7191 17831 7197
rect 17773 7188 17785 7191
rect 17552 7160 17785 7188
rect 17552 7148 17558 7160
rect 17773 7157 17785 7160
rect 17819 7157 17831 7191
rect 18322 7188 18328 7200
rect 18283 7160 18328 7188
rect 17773 7151 17831 7157
rect 18322 7148 18328 7160
rect 18380 7148 18386 7200
rect 20346 7188 20352 7200
rect 20307 7160 20352 7188
rect 20346 7148 20352 7160
rect 20404 7148 20410 7200
rect 1104 7098 22816 7120
rect 1104 7046 8982 7098
rect 9034 7046 9046 7098
rect 9098 7046 9110 7098
rect 9162 7046 9174 7098
rect 9226 7046 16982 7098
rect 17034 7046 17046 7098
rect 17098 7046 17110 7098
rect 17162 7046 17174 7098
rect 17226 7046 22816 7098
rect 1104 7024 22816 7046
rect 2314 6944 2320 6996
rect 2372 6984 2378 6996
rect 2777 6987 2835 6993
rect 2777 6984 2789 6987
rect 2372 6956 2789 6984
rect 2372 6944 2378 6956
rect 2777 6953 2789 6956
rect 2823 6953 2835 6987
rect 2777 6947 2835 6953
rect 3142 6944 3148 6996
rect 3200 6984 3206 6996
rect 3237 6987 3295 6993
rect 3237 6984 3249 6987
rect 3200 6956 3249 6984
rect 3200 6944 3206 6956
rect 3237 6953 3249 6956
rect 3283 6984 3295 6987
rect 4157 6987 4215 6993
rect 4157 6984 4169 6987
rect 3283 6956 4169 6984
rect 3283 6953 3295 6956
rect 3237 6947 3295 6953
rect 4157 6953 4169 6956
rect 4203 6953 4215 6987
rect 4157 6947 4215 6953
rect 5261 6987 5319 6993
rect 5261 6953 5273 6987
rect 5307 6984 5319 6987
rect 5442 6984 5448 6996
rect 5307 6956 5448 6984
rect 5307 6953 5319 6956
rect 5261 6947 5319 6953
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 7282 6984 7288 6996
rect 7243 6956 7288 6984
rect 7282 6944 7288 6956
rect 7340 6944 7346 6996
rect 7650 6944 7656 6996
rect 7708 6984 7714 6996
rect 7837 6987 7895 6993
rect 7837 6984 7849 6987
rect 7708 6956 7849 6984
rect 7708 6944 7714 6956
rect 7837 6953 7849 6956
rect 7883 6953 7895 6987
rect 7837 6947 7895 6953
rect 10873 6987 10931 6993
rect 10873 6953 10885 6987
rect 10919 6984 10931 6987
rect 10962 6984 10968 6996
rect 10919 6956 10968 6984
rect 10919 6953 10931 6956
rect 10873 6947 10931 6953
rect 5629 6919 5687 6925
rect 5629 6885 5641 6919
rect 5675 6916 5687 6919
rect 7009 6919 7067 6925
rect 7009 6916 7021 6919
rect 5675 6888 7021 6916
rect 5675 6885 5687 6888
rect 5629 6879 5687 6885
rect 7009 6885 7021 6888
rect 7055 6916 7067 6919
rect 7466 6916 7472 6928
rect 7055 6888 7472 6916
rect 7055 6885 7067 6888
rect 7009 6879 7067 6885
rect 7466 6876 7472 6888
rect 7524 6876 7530 6928
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 1762 6848 1768 6860
rect 1719 6820 1768 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 2406 6848 2412 6860
rect 2367 6820 2412 6848
rect 2406 6808 2412 6820
rect 2464 6808 2470 6860
rect 4338 6848 4344 6860
rect 4299 6820 4344 6848
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6848 4675 6851
rect 5074 6848 5080 6860
rect 4663 6820 5080 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 3789 6783 3847 6789
rect 3789 6749 3801 6783
rect 3835 6780 3847 6783
rect 4246 6780 4252 6792
rect 3835 6752 4252 6780
rect 3835 6749 3847 6752
rect 3789 6743 3847 6749
rect 4246 6740 4252 6752
rect 4304 6780 4310 6792
rect 4632 6780 4660 6811
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 5718 6808 5724 6860
rect 5776 6857 5782 6860
rect 5776 6851 5834 6857
rect 5776 6817 5788 6851
rect 5822 6848 5834 6851
rect 6638 6848 6644 6860
rect 5822 6820 6644 6848
rect 5822 6817 5834 6820
rect 5776 6811 5834 6817
rect 5776 6808 5782 6811
rect 6638 6808 6644 6820
rect 6696 6808 6702 6860
rect 4304 6752 4660 6780
rect 4304 6740 4310 6752
rect 4706 6740 4712 6792
rect 4764 6780 4770 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 4764 6752 6009 6780
rect 4764 6740 4770 6752
rect 5997 6749 6009 6752
rect 6043 6780 6055 6783
rect 7852 6780 7880 6947
rect 10962 6944 10968 6956
rect 11020 6984 11026 6996
rect 11606 6984 11612 6996
rect 11020 6956 11612 6984
rect 11020 6944 11026 6956
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 12802 6984 12808 6996
rect 12763 6956 12808 6984
rect 12802 6944 12808 6956
rect 12860 6944 12866 6996
rect 13354 6984 13360 6996
rect 13315 6956 13360 6984
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 17954 6944 17960 6996
rect 18012 6984 18018 6996
rect 18049 6987 18107 6993
rect 18049 6984 18061 6987
rect 18012 6956 18061 6984
rect 18012 6944 18018 6956
rect 18049 6953 18061 6956
rect 18095 6953 18107 6987
rect 18782 6984 18788 6996
rect 18743 6956 18788 6984
rect 18049 6947 18107 6953
rect 18782 6944 18788 6956
rect 18840 6944 18846 6996
rect 19334 6984 19340 6996
rect 19295 6956 19340 6984
rect 19334 6944 19340 6956
rect 19392 6944 19398 6996
rect 8202 6916 8208 6928
rect 8163 6888 8208 6916
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 11422 6876 11428 6928
rect 11480 6916 11486 6928
rect 11977 6919 12035 6925
rect 11977 6916 11989 6919
rect 11480 6888 11989 6916
rect 11480 6876 11486 6888
rect 11977 6885 11989 6888
rect 12023 6916 12035 6919
rect 14090 6916 14096 6928
rect 12023 6888 14096 6916
rect 12023 6885 12035 6888
rect 11977 6879 12035 6885
rect 14090 6876 14096 6888
rect 14148 6876 14154 6928
rect 16390 6916 16396 6928
rect 16351 6888 16396 6916
rect 16390 6876 16396 6888
rect 16448 6876 16454 6928
rect 21085 6919 21143 6925
rect 21085 6885 21097 6919
rect 21131 6916 21143 6919
rect 21266 6916 21272 6928
rect 21131 6888 21272 6916
rect 21131 6885 21143 6888
rect 21085 6879 21143 6885
rect 21266 6876 21272 6888
rect 21324 6876 21330 6928
rect 9950 6848 9956 6860
rect 9911 6820 9956 6848
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 11238 6848 11244 6860
rect 11199 6820 11244 6848
rect 11238 6808 11244 6820
rect 11296 6808 11302 6860
rect 12158 6848 12164 6860
rect 11421 6820 12164 6848
rect 8113 6783 8171 6789
rect 8113 6780 8125 6783
rect 6043 6752 7788 6780
rect 7852 6752 8125 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 4614 6672 4620 6724
rect 4672 6712 4678 6724
rect 6089 6715 6147 6721
rect 6089 6712 6101 6715
rect 4672 6684 6101 6712
rect 4672 6672 4678 6684
rect 6089 6681 6101 6684
rect 6135 6681 6147 6715
rect 7760 6712 7788 6752
rect 8113 6749 8125 6752
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 8757 6783 8815 6789
rect 8757 6749 8769 6783
rect 8803 6780 8815 6783
rect 8846 6780 8852 6792
rect 8803 6752 8852 6780
rect 8803 6749 8815 6752
rect 8757 6743 8815 6749
rect 8846 6740 8852 6752
rect 8904 6740 8910 6792
rect 9122 6740 9128 6792
rect 9180 6780 9186 6792
rect 11421 6789 11449 6820
rect 12158 6808 12164 6820
rect 12216 6848 12222 6860
rect 12710 6848 12716 6860
rect 12216 6820 12716 6848
rect 12216 6808 12222 6820
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 13630 6848 13636 6860
rect 13591 6820 13636 6848
rect 13630 6808 13636 6820
rect 13688 6808 13694 6860
rect 18322 6808 18328 6860
rect 18380 6848 18386 6860
rect 18417 6851 18475 6857
rect 18417 6848 18429 6851
rect 18380 6820 18429 6848
rect 18380 6808 18386 6820
rect 18417 6817 18429 6820
rect 18463 6817 18475 6851
rect 18417 6811 18475 6817
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9180 6752 9689 6780
rect 9180 6740 9186 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 11388 6783 11449 6789
rect 11388 6749 11400 6783
rect 11434 6752 11449 6783
rect 11606 6780 11612 6792
rect 11567 6752 11612 6780
rect 11434 6749 11446 6752
rect 11388 6743 11446 6749
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 16298 6780 16304 6792
rect 16259 6752 16304 6780
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 20993 6783 21051 6789
rect 20993 6749 21005 6783
rect 21039 6780 21051 6783
rect 21450 6780 21456 6792
rect 21039 6752 21456 6780
rect 21039 6749 21051 6752
rect 20993 6743 21051 6749
rect 21450 6740 21456 6752
rect 21508 6740 21514 6792
rect 8478 6712 8484 6724
rect 7760 6684 8484 6712
rect 6089 6675 6147 6681
rect 8478 6672 8484 6684
rect 8536 6672 8542 6724
rect 11054 6672 11060 6724
rect 11112 6712 11118 6724
rect 11517 6715 11575 6721
rect 11517 6712 11529 6715
rect 11112 6684 11529 6712
rect 11112 6672 11118 6684
rect 11517 6681 11529 6684
rect 11563 6712 11575 6715
rect 11882 6712 11888 6724
rect 11563 6684 11888 6712
rect 11563 6681 11575 6684
rect 11517 6675 11575 6681
rect 11882 6672 11888 6684
rect 11940 6672 11946 6724
rect 16850 6712 16856 6724
rect 16811 6684 16856 6712
rect 16850 6672 16856 6684
rect 16908 6672 16914 6724
rect 21545 6715 21603 6721
rect 21545 6681 21557 6715
rect 21591 6681 21603 6715
rect 21545 6675 21603 6681
rect 4798 6604 4804 6656
rect 4856 6644 4862 6656
rect 5905 6647 5963 6653
rect 5905 6644 5917 6647
rect 4856 6616 5917 6644
rect 4856 6604 4862 6616
rect 5905 6613 5917 6616
rect 5951 6644 5963 6647
rect 6178 6644 6184 6656
rect 5951 6616 6184 6644
rect 5951 6613 5963 6616
rect 5905 6607 5963 6613
rect 6178 6604 6184 6616
rect 6236 6604 6242 6656
rect 8754 6604 8760 6656
rect 8812 6644 8818 6656
rect 9033 6647 9091 6653
rect 9033 6644 9045 6647
rect 8812 6616 9045 6644
rect 8812 6604 8818 6616
rect 9033 6613 9045 6616
rect 9079 6613 9091 6647
rect 9033 6607 9091 6613
rect 10870 6604 10876 6656
rect 10928 6644 10934 6656
rect 12434 6644 12440 6656
rect 10928 6616 12440 6644
rect 10928 6604 10934 6616
rect 12434 6604 12440 6616
rect 12492 6604 12498 6656
rect 15010 6604 15016 6656
rect 15068 6644 15074 6656
rect 21358 6644 21364 6656
rect 15068 6616 21364 6644
rect 15068 6604 15074 6616
rect 21358 6604 21364 6616
rect 21416 6644 21422 6656
rect 21560 6644 21588 6675
rect 21416 6616 21588 6644
rect 21416 6604 21422 6616
rect 1104 6554 22816 6576
rect 1104 6502 4982 6554
rect 5034 6502 5046 6554
rect 5098 6502 5110 6554
rect 5162 6502 5174 6554
rect 5226 6502 12982 6554
rect 13034 6502 13046 6554
rect 13098 6502 13110 6554
rect 13162 6502 13174 6554
rect 13226 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 22816 6554
rect 1104 6480 22816 6502
rect 2409 6443 2467 6449
rect 2409 6409 2421 6443
rect 2455 6440 2467 6443
rect 3694 6440 3700 6452
rect 2455 6412 3700 6440
rect 2455 6409 2467 6412
rect 2409 6403 2467 6409
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6304 2099 6307
rect 2406 6304 2412 6316
rect 2087 6276 2412 6304
rect 2087 6273 2099 6276
rect 2041 6267 2099 6273
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 1394 6236 1400 6248
rect 1307 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6236 1458 6248
rect 1946 6236 1952 6248
rect 1452 6208 1952 6236
rect 1452 6196 1458 6208
rect 1946 6196 1952 6208
rect 2004 6196 2010 6248
rect 2516 6245 2544 6412
rect 3694 6400 3700 6412
rect 3752 6400 3758 6452
rect 4706 6400 4712 6452
rect 4764 6440 4770 6452
rect 4801 6443 4859 6449
rect 4801 6440 4813 6443
rect 4764 6412 4813 6440
rect 4764 6400 4770 6412
rect 4801 6409 4813 6412
rect 4847 6409 4859 6443
rect 6178 6440 6184 6452
rect 6139 6412 6184 6440
rect 4801 6403 4859 6409
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 8202 6400 8208 6452
rect 8260 6440 8266 6452
rect 8389 6443 8447 6449
rect 8389 6440 8401 6443
rect 8260 6412 8401 6440
rect 8260 6400 8266 6412
rect 8389 6409 8401 6412
rect 8435 6440 8447 6443
rect 8570 6440 8576 6452
rect 8435 6412 8576 6440
rect 8435 6409 8447 6412
rect 8389 6403 8447 6409
rect 8570 6400 8576 6412
rect 8628 6440 8634 6452
rect 9950 6440 9956 6452
rect 8628 6412 9956 6440
rect 8628 6400 8634 6412
rect 9950 6400 9956 6412
rect 10008 6400 10014 6452
rect 10413 6443 10471 6449
rect 10413 6409 10425 6443
rect 10459 6440 10471 6443
rect 10962 6440 10968 6452
rect 10459 6412 10968 6440
rect 10459 6409 10471 6412
rect 10413 6403 10471 6409
rect 3237 6375 3295 6381
rect 3237 6341 3249 6375
rect 3283 6372 3295 6375
rect 4338 6372 4344 6384
rect 3283 6344 4344 6372
rect 3283 6341 3295 6344
rect 3237 6335 3295 6341
rect 4338 6332 4344 6344
rect 4396 6332 4402 6384
rect 8110 6332 8116 6384
rect 8168 6372 8174 6384
rect 10428 6372 10456 6403
rect 10962 6400 10968 6412
rect 11020 6440 11026 6452
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 11020 6412 11529 6440
rect 11020 6400 11026 6412
rect 11517 6409 11529 6412
rect 11563 6409 11575 6443
rect 11882 6440 11888 6452
rect 11843 6412 11888 6440
rect 11517 6403 11575 6409
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12710 6440 12716 6452
rect 12671 6412 12716 6440
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 14826 6440 14832 6452
rect 14787 6412 14832 6440
rect 14826 6400 14832 6412
rect 14884 6400 14890 6452
rect 15838 6440 15844 6452
rect 15751 6412 15844 6440
rect 15838 6400 15844 6412
rect 15896 6440 15902 6452
rect 16301 6443 16359 6449
rect 16301 6440 16313 6443
rect 15896 6412 16313 6440
rect 15896 6400 15902 6412
rect 16301 6409 16313 6412
rect 16347 6440 16359 6443
rect 16390 6440 16396 6452
rect 16347 6412 16396 6440
rect 16347 6409 16359 6412
rect 16301 6403 16359 6409
rect 16390 6400 16396 6412
rect 16448 6400 16454 6452
rect 18322 6400 18328 6452
rect 18380 6440 18386 6452
rect 18785 6443 18843 6449
rect 18785 6440 18797 6443
rect 18380 6412 18797 6440
rect 18380 6400 18386 6412
rect 18785 6409 18797 6412
rect 18831 6409 18843 6443
rect 20346 6440 20352 6452
rect 20307 6412 20352 6440
rect 18785 6403 18843 6409
rect 20346 6400 20352 6412
rect 20404 6400 20410 6452
rect 21266 6400 21272 6452
rect 21324 6440 21330 6452
rect 21545 6443 21603 6449
rect 21545 6440 21557 6443
rect 21324 6412 21557 6440
rect 21324 6400 21330 6412
rect 21545 6409 21557 6412
rect 21591 6409 21603 6443
rect 21545 6403 21603 6409
rect 8168 6344 10456 6372
rect 21177 6375 21235 6381
rect 8168 6332 8174 6344
rect 21177 6341 21189 6375
rect 21223 6372 21235 6375
rect 21358 6372 21364 6384
rect 21223 6344 21364 6372
rect 21223 6341 21235 6344
rect 21177 6335 21235 6341
rect 21358 6332 21364 6344
rect 21416 6332 21422 6384
rect 7466 6304 7472 6316
rect 3988 6276 4154 6304
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6205 2559 6239
rect 2501 6199 2559 6205
rect 3605 6239 3663 6245
rect 3605 6205 3617 6239
rect 3651 6236 3663 6239
rect 3786 6236 3792 6248
rect 3651 6208 3792 6236
rect 3651 6205 3663 6208
rect 3605 6199 3663 6205
rect 3786 6196 3792 6208
rect 3844 6236 3850 6248
rect 3988 6245 4016 6276
rect 3973 6239 4031 6245
rect 3973 6236 3985 6239
rect 3844 6208 3985 6236
rect 3844 6196 3850 6208
rect 3973 6205 3985 6208
rect 4019 6205 4031 6239
rect 3973 6199 4031 6205
rect 198 6128 204 6180
rect 256 6168 262 6180
rect 256 6140 2728 6168
rect 256 6128 262 6140
rect 106 6060 112 6112
rect 164 6100 170 6112
rect 2700 6109 2728 6140
rect 1581 6103 1639 6109
rect 1581 6100 1593 6103
rect 164 6072 1593 6100
rect 164 6060 170 6072
rect 1581 6069 1593 6072
rect 1627 6069 1639 6103
rect 1581 6063 1639 6069
rect 2685 6103 2743 6109
rect 2685 6069 2697 6103
rect 2731 6069 2743 6103
rect 2685 6063 2743 6069
rect 3602 6060 3608 6112
rect 3660 6100 3666 6112
rect 3789 6103 3847 6109
rect 3789 6100 3801 6103
rect 3660 6072 3801 6100
rect 3660 6060 3666 6072
rect 3789 6069 3801 6072
rect 3835 6069 3847 6103
rect 4126 6100 4154 6276
rect 7208 6276 7472 6304
rect 7208 6248 7236 6276
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 8846 6264 8852 6316
rect 8904 6304 8910 6316
rect 9309 6307 9367 6313
rect 9309 6304 9321 6307
rect 8904 6276 9321 6304
rect 8904 6264 8910 6276
rect 9309 6273 9321 6276
rect 9355 6273 9367 6307
rect 9309 6267 9367 6273
rect 14734 6264 14740 6316
rect 14792 6304 14798 6316
rect 14921 6307 14979 6313
rect 14921 6304 14933 6307
rect 14792 6276 14933 6304
rect 14792 6264 14798 6276
rect 14921 6273 14933 6276
rect 14967 6273 14979 6307
rect 14921 6267 14979 6273
rect 16298 6264 16304 6316
rect 16356 6304 16362 6316
rect 16577 6307 16635 6313
rect 16577 6304 16589 6307
rect 16356 6276 16589 6304
rect 16356 6264 16362 6276
rect 16577 6273 16589 6276
rect 16623 6273 16635 6307
rect 16577 6267 16635 6273
rect 18509 6307 18567 6313
rect 18509 6273 18521 6307
rect 18555 6304 18567 6307
rect 18782 6304 18788 6316
rect 18555 6276 18788 6304
rect 18555 6273 18567 6276
rect 18509 6267 18567 6273
rect 18782 6264 18788 6276
rect 18840 6264 18846 6316
rect 20073 6307 20131 6313
rect 20073 6273 20085 6307
rect 20119 6304 20131 6307
rect 21450 6304 21456 6316
rect 20119 6276 21456 6304
rect 20119 6273 20131 6276
rect 20073 6267 20131 6273
rect 21450 6264 21456 6276
rect 21508 6264 21514 6316
rect 4246 6236 4252 6248
rect 4207 6208 4252 6236
rect 4246 6196 4252 6208
rect 4304 6196 4310 6248
rect 4798 6196 4804 6248
rect 4856 6236 4862 6248
rect 5169 6239 5227 6245
rect 5169 6236 5181 6239
rect 4856 6208 5181 6236
rect 4856 6196 4862 6208
rect 5169 6205 5181 6208
rect 5215 6236 5227 6239
rect 5537 6239 5595 6245
rect 5537 6236 5549 6239
rect 5215 6208 5549 6236
rect 5215 6205 5227 6208
rect 5169 6199 5227 6205
rect 5537 6205 5549 6208
rect 5583 6205 5595 6239
rect 7190 6236 7196 6248
rect 7103 6208 7196 6236
rect 5537 6199 5595 6205
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 7282 6196 7288 6248
rect 7340 6236 7346 6248
rect 7377 6239 7435 6245
rect 7377 6236 7389 6239
rect 7340 6208 7389 6236
rect 7340 6196 7346 6208
rect 7377 6205 7389 6208
rect 7423 6205 7435 6239
rect 7377 6199 7435 6205
rect 7558 6196 7564 6248
rect 7616 6236 7622 6248
rect 7745 6239 7803 6245
rect 7745 6236 7757 6239
rect 7616 6208 7757 6236
rect 7616 6196 7622 6208
rect 7745 6205 7757 6208
rect 7791 6236 7803 6239
rect 7926 6236 7932 6248
rect 7791 6208 7932 6236
rect 7791 6205 7803 6208
rect 7745 6199 7803 6205
rect 7926 6196 7932 6208
rect 7984 6196 7990 6248
rect 10962 6236 10968 6248
rect 10923 6208 10968 6236
rect 10962 6196 10968 6208
rect 11020 6196 11026 6248
rect 13354 6196 13360 6248
rect 13412 6236 13418 6248
rect 13633 6239 13691 6245
rect 13633 6236 13645 6239
rect 13412 6208 13645 6236
rect 13412 6196 13418 6208
rect 13633 6205 13645 6208
rect 13679 6236 13691 6239
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13679 6208 14013 6236
rect 13679 6205 13691 6208
rect 13633 6199 13691 6205
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14001 6199 14059 6205
rect 16828 6239 16886 6245
rect 16828 6205 16840 6239
rect 16874 6236 16886 6239
rect 16874 6208 17356 6236
rect 16874 6205 16886 6208
rect 16828 6199 16886 6205
rect 5350 6168 5356 6180
rect 5311 6140 5356 6168
rect 5350 6128 5356 6140
rect 5408 6128 5414 6180
rect 5905 6171 5963 6177
rect 5905 6137 5917 6171
rect 5951 6168 5963 6171
rect 6362 6168 6368 6180
rect 5951 6140 6368 6168
rect 5951 6137 5963 6140
rect 5905 6131 5963 6137
rect 6362 6128 6368 6140
rect 6420 6168 6426 6180
rect 8662 6168 8668 6180
rect 6420 6140 8668 6168
rect 6420 6128 6426 6140
rect 8662 6128 8668 6140
rect 8720 6128 8726 6180
rect 8754 6128 8760 6180
rect 8812 6168 8818 6180
rect 9033 6171 9091 6177
rect 9033 6168 9045 6171
rect 8812 6140 9045 6168
rect 8812 6128 8818 6140
rect 9033 6137 9045 6140
rect 9079 6137 9091 6171
rect 9033 6131 9091 6137
rect 9122 6128 9128 6180
rect 9180 6168 9186 6180
rect 10502 6168 10508 6180
rect 9180 6140 9225 6168
rect 10463 6140 10508 6168
rect 9180 6128 9186 6140
rect 10502 6128 10508 6140
rect 10560 6128 10566 6180
rect 12710 6128 12716 6180
rect 12768 6168 12774 6180
rect 14826 6168 14832 6180
rect 12768 6140 14832 6168
rect 12768 6128 12774 6140
rect 14826 6128 14832 6140
rect 14884 6168 14890 6180
rect 15242 6171 15300 6177
rect 15242 6168 15254 6171
rect 14884 6140 15254 6168
rect 14884 6128 14890 6140
rect 15242 6137 15254 6140
rect 15288 6137 15300 6171
rect 15242 6131 15300 6137
rect 6641 6103 6699 6109
rect 6641 6100 6653 6103
rect 4126 6072 6653 6100
rect 3789 6063 3847 6069
rect 6641 6069 6653 6072
rect 6687 6100 6699 6103
rect 7558 6100 7564 6112
rect 6687 6072 7564 6100
rect 6687 6069 6699 6072
rect 6641 6063 6699 6069
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 7834 6100 7840 6112
rect 7795 6072 7840 6100
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8849 6103 8907 6109
rect 8849 6069 8861 6103
rect 8895 6100 8907 6103
rect 9140 6100 9168 6128
rect 13262 6100 13268 6112
rect 8895 6072 9168 6100
rect 13223 6072 13268 6100
rect 8895 6069 8907 6072
rect 8849 6063 8907 6069
rect 13262 6060 13268 6072
rect 13320 6060 13326 6112
rect 16666 6060 16672 6112
rect 16724 6100 16730 6112
rect 17328 6109 17356 6208
rect 20622 6168 20628 6180
rect 20583 6140 20628 6168
rect 20622 6128 20628 6140
rect 20680 6128 20686 6180
rect 20717 6171 20775 6177
rect 20717 6137 20729 6171
rect 20763 6137 20775 6171
rect 20717 6131 20775 6137
rect 16899 6103 16957 6109
rect 16899 6100 16911 6103
rect 16724 6072 16911 6100
rect 16724 6060 16730 6072
rect 16899 6069 16911 6072
rect 16945 6069 16957 6103
rect 16899 6063 16957 6069
rect 17313 6103 17371 6109
rect 17313 6069 17325 6103
rect 17359 6100 17371 6103
rect 18046 6100 18052 6112
rect 17359 6072 18052 6100
rect 17359 6069 17371 6072
rect 17313 6063 17371 6069
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 20346 6060 20352 6112
rect 20404 6100 20410 6112
rect 20732 6100 20760 6131
rect 20404 6072 20760 6100
rect 20404 6060 20410 6072
rect 1104 6010 22816 6032
rect 1104 5958 8982 6010
rect 9034 5958 9046 6010
rect 9098 5958 9110 6010
rect 9162 5958 9174 6010
rect 9226 5958 16982 6010
rect 17034 5958 17046 6010
rect 17098 5958 17110 6010
rect 17162 5958 17174 6010
rect 17226 5958 22816 6010
rect 1104 5936 22816 5958
rect 2038 5856 2044 5908
rect 2096 5896 2102 5908
rect 2869 5899 2927 5905
rect 2869 5896 2881 5899
rect 2096 5868 2881 5896
rect 2096 5856 2102 5868
rect 2869 5865 2881 5868
rect 2915 5896 2927 5899
rect 4157 5899 4215 5905
rect 4157 5896 4169 5899
rect 2915 5868 4169 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 4157 5865 4169 5868
rect 4203 5865 4215 5899
rect 8018 5896 8024 5908
rect 7979 5868 8024 5896
rect 4157 5859 4215 5865
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 8570 5896 8576 5908
rect 8531 5868 8576 5896
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 8662 5856 8668 5908
rect 8720 5896 8726 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 8720 5868 9045 5896
rect 8720 5856 8726 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 11238 5856 11244 5908
rect 11296 5896 11302 5908
rect 11885 5899 11943 5905
rect 11885 5896 11897 5899
rect 11296 5868 11897 5896
rect 11296 5856 11302 5868
rect 11885 5865 11897 5868
rect 11931 5865 11943 5899
rect 13354 5896 13360 5908
rect 13315 5868 13360 5896
rect 11885 5859 11943 5865
rect 13354 5856 13360 5868
rect 13412 5856 13418 5908
rect 13630 5896 13636 5908
rect 13591 5868 13636 5896
rect 13630 5856 13636 5868
rect 13688 5856 13694 5908
rect 14734 5856 14740 5908
rect 14792 5896 14798 5908
rect 14921 5899 14979 5905
rect 14921 5896 14933 5899
rect 14792 5868 14933 5896
rect 14792 5856 14798 5868
rect 14921 5865 14933 5868
rect 14967 5865 14979 5899
rect 14921 5859 14979 5865
rect 18417 5899 18475 5905
rect 18417 5865 18429 5899
rect 18463 5896 18475 5899
rect 18782 5896 18788 5908
rect 18463 5868 18788 5896
rect 18463 5865 18475 5868
rect 18417 5859 18475 5865
rect 18782 5856 18788 5868
rect 18840 5856 18846 5908
rect 20162 5896 20168 5908
rect 20075 5868 20168 5896
rect 20162 5856 20168 5868
rect 20220 5896 20226 5908
rect 20438 5896 20444 5908
rect 20220 5868 20444 5896
rect 20220 5856 20226 5868
rect 20438 5856 20444 5868
rect 20496 5856 20502 5908
rect 20622 5896 20628 5908
rect 20583 5868 20628 5896
rect 20622 5856 20628 5868
rect 20680 5896 20686 5908
rect 21039 5899 21097 5905
rect 21039 5896 21051 5899
rect 20680 5868 21051 5896
rect 20680 5856 20686 5868
rect 21039 5865 21051 5868
rect 21085 5865 21097 5899
rect 21039 5859 21097 5865
rect 3513 5831 3571 5837
rect 3513 5797 3525 5831
rect 3559 5828 3571 5831
rect 4246 5828 4252 5840
rect 3559 5800 4252 5828
rect 3559 5797 3571 5800
rect 3513 5791 3571 5797
rect 4246 5788 4252 5800
rect 4304 5788 4310 5840
rect 12618 5788 12624 5840
rect 12676 5828 12682 5840
rect 12758 5831 12816 5837
rect 12758 5828 12770 5831
rect 12676 5800 12770 5828
rect 12676 5788 12682 5800
rect 12758 5797 12770 5800
rect 12804 5797 12816 5831
rect 16574 5828 16580 5840
rect 16535 5800 16580 5828
rect 12758 5791 12816 5797
rect 16574 5788 16580 5800
rect 16632 5788 16638 5840
rect 21266 5828 21272 5840
rect 20983 5800 21272 5828
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5760 1731 5763
rect 1857 5763 1915 5769
rect 1857 5760 1869 5763
rect 1719 5732 1869 5760
rect 1719 5729 1731 5732
rect 1673 5723 1731 5729
rect 1857 5729 1869 5732
rect 1903 5760 1915 5763
rect 2958 5760 2964 5772
rect 1903 5732 2964 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 2958 5720 2964 5732
rect 3016 5720 3022 5772
rect 4338 5760 4344 5772
rect 4299 5732 4344 5760
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 4614 5760 4620 5772
rect 4575 5732 4620 5760
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 5994 5760 6000 5772
rect 5955 5732 6000 5760
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 6270 5760 6276 5772
rect 6231 5732 6276 5760
rect 6270 5720 6276 5732
rect 6328 5760 6334 5772
rect 6825 5763 6883 5769
rect 6825 5760 6837 5763
rect 6328 5732 6837 5760
rect 6328 5720 6334 5732
rect 6825 5729 6837 5732
rect 6871 5729 6883 5763
rect 6825 5723 6883 5729
rect 7653 5763 7711 5769
rect 7653 5729 7665 5763
rect 7699 5760 7711 5763
rect 7834 5760 7840 5772
rect 7699 5732 7840 5760
rect 7699 5729 7711 5732
rect 7653 5723 7711 5729
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 10870 5760 10876 5772
rect 10831 5732 10876 5760
rect 10870 5720 10876 5732
rect 10928 5720 10934 5772
rect 11422 5760 11428 5772
rect 11383 5732 11428 5760
rect 11422 5720 11428 5732
rect 11480 5720 11486 5772
rect 20983 5769 21011 5800
rect 21266 5788 21272 5800
rect 21324 5828 21330 5840
rect 21726 5828 21732 5840
rect 21324 5800 21732 5828
rect 21324 5788 21330 5800
rect 21726 5788 21732 5800
rect 21784 5788 21790 5840
rect 20968 5763 21026 5769
rect 20968 5729 20980 5763
rect 21014 5729 21026 5763
rect 20968 5723 21026 5729
rect 1762 5692 1768 5704
rect 1723 5664 1768 5692
rect 1762 5652 1768 5664
rect 1820 5652 1826 5704
rect 3881 5695 3939 5701
rect 3881 5661 3893 5695
rect 3927 5692 3939 5695
rect 4632 5692 4660 5720
rect 3927 5664 4660 5692
rect 3927 5661 3939 5664
rect 3881 5655 3939 5661
rect 5350 5652 5356 5704
rect 5408 5692 5414 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 5408 5664 5457 5692
rect 5408 5652 5414 5664
rect 5445 5661 5457 5664
rect 5491 5692 5503 5695
rect 5810 5692 5816 5704
rect 5491 5664 5816 5692
rect 5491 5661 5503 5664
rect 5445 5655 5503 5661
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 11609 5695 11667 5701
rect 11609 5661 11621 5695
rect 11655 5692 11667 5695
rect 12434 5692 12440 5704
rect 11655 5664 12440 5692
rect 11655 5661 11667 5664
rect 11609 5655 11667 5661
rect 12434 5652 12440 5664
rect 12492 5652 12498 5704
rect 16485 5695 16543 5701
rect 16485 5661 16497 5695
rect 16531 5692 16543 5695
rect 16666 5692 16672 5704
rect 16531 5664 16672 5692
rect 16531 5661 16543 5664
rect 16485 5655 16543 5661
rect 16666 5652 16672 5664
rect 16724 5652 16730 5704
rect 16850 5692 16856 5704
rect 16811 5664 16856 5692
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 5813 5559 5871 5565
rect 5813 5525 5825 5559
rect 5859 5556 5871 5559
rect 6638 5556 6644 5568
rect 5859 5528 6644 5556
rect 5859 5525 5871 5528
rect 5813 5519 5871 5525
rect 6638 5516 6644 5528
rect 6696 5556 6702 5568
rect 7285 5559 7343 5565
rect 7285 5556 7297 5559
rect 6696 5528 7297 5556
rect 6696 5516 6702 5528
rect 7285 5525 7297 5528
rect 7331 5556 7343 5559
rect 9398 5556 9404 5568
rect 7331 5528 9404 5556
rect 7331 5525 7343 5528
rect 7285 5519 7343 5525
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 1104 5466 22816 5488
rect 1104 5414 4982 5466
rect 5034 5414 5046 5466
rect 5098 5414 5110 5466
rect 5162 5414 5174 5466
rect 5226 5414 12982 5466
rect 13034 5414 13046 5466
rect 13098 5414 13110 5466
rect 13162 5414 13174 5466
rect 13226 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 22816 5466
rect 1104 5392 22816 5414
rect 2958 5352 2964 5364
rect 2919 5324 2964 5352
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 3786 5352 3792 5364
rect 3747 5324 3792 5352
rect 3786 5312 3792 5324
rect 3844 5312 3850 5364
rect 6178 5312 6184 5364
rect 6236 5352 6242 5364
rect 6549 5355 6607 5361
rect 6549 5352 6561 5355
rect 6236 5324 6561 5352
rect 6236 5312 6242 5324
rect 6549 5321 6561 5324
rect 6595 5352 6607 5355
rect 7101 5355 7159 5361
rect 7101 5352 7113 5355
rect 6595 5324 7113 5352
rect 6595 5321 6607 5324
rect 6549 5315 6607 5321
rect 7101 5321 7113 5324
rect 7147 5321 7159 5355
rect 7282 5352 7288 5364
rect 7243 5324 7288 5352
rect 7101 5315 7159 5321
rect 14 5244 20 5296
rect 72 5284 78 5296
rect 5261 5287 5319 5293
rect 5261 5284 5273 5287
rect 72 5256 5273 5284
rect 72 5244 78 5256
rect 5261 5253 5273 5256
rect 5307 5253 5319 5287
rect 7116 5284 7144 5315
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 7929 5355 7987 5361
rect 7929 5321 7941 5355
rect 7975 5352 7987 5355
rect 8018 5352 8024 5364
rect 7975 5324 8024 5352
rect 7975 5321 7987 5324
rect 7929 5315 7987 5321
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 8662 5312 8668 5364
rect 8720 5352 8726 5364
rect 9171 5355 9229 5361
rect 9171 5352 9183 5355
rect 8720 5324 9183 5352
rect 8720 5312 8726 5324
rect 9171 5321 9183 5324
rect 9217 5321 9229 5355
rect 9171 5315 9229 5321
rect 9398 5312 9404 5364
rect 9456 5352 9462 5364
rect 10946 5355 11004 5361
rect 10946 5352 10958 5355
rect 9456 5324 10958 5352
rect 9456 5312 9462 5324
rect 10946 5321 10958 5324
rect 10992 5352 11004 5355
rect 12158 5352 12164 5364
rect 10992 5324 12164 5352
rect 10992 5321 11004 5324
rect 10946 5315 11004 5321
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 13265 5355 13323 5361
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 13354 5352 13360 5364
rect 13311 5324 13360 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 15838 5352 15844 5364
rect 15799 5324 15844 5352
rect 15838 5312 15844 5324
rect 15896 5312 15902 5364
rect 21177 5355 21235 5361
rect 21177 5321 21189 5355
rect 21223 5352 21235 5355
rect 21266 5352 21272 5364
rect 21223 5324 21272 5352
rect 21223 5321 21235 5324
rect 21177 5315 21235 5321
rect 21266 5312 21272 5324
rect 21324 5312 21330 5364
rect 8849 5287 8907 5293
rect 8849 5284 8861 5287
rect 7116 5256 8861 5284
rect 5261 5247 5319 5253
rect 8849 5253 8861 5256
rect 8895 5284 8907 5287
rect 9309 5287 9367 5293
rect 9309 5284 9321 5287
rect 8895 5256 9321 5284
rect 8895 5253 8907 5256
rect 8849 5247 8907 5253
rect 9309 5253 9321 5256
rect 9355 5284 9367 5287
rect 10594 5284 10600 5296
rect 9355 5256 10600 5284
rect 9355 5253 9367 5256
rect 9309 5247 9367 5253
rect 2038 5216 2044 5228
rect 1999 5188 2044 5216
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 3421 5219 3479 5225
rect 3421 5185 3433 5219
rect 3467 5216 3479 5219
rect 4338 5216 4344 5228
rect 3467 5188 4344 5216
rect 3467 5185 3479 5188
rect 3421 5179 3479 5185
rect 4338 5176 4344 5188
rect 4396 5176 4402 5228
rect 3786 5108 3792 5160
rect 3844 5148 3850 5160
rect 3881 5151 3939 5157
rect 3881 5148 3893 5151
rect 3844 5120 3893 5148
rect 3844 5108 3850 5120
rect 3881 5117 3893 5120
rect 3927 5117 3939 5151
rect 3881 5111 3939 5117
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5148 4491 5151
rect 4614 5148 4620 5160
rect 4479 5120 4620 5148
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 5276 5148 5304 5247
rect 10594 5244 10600 5256
rect 10652 5284 10658 5296
rect 11057 5287 11115 5293
rect 11057 5284 11069 5287
rect 10652 5256 11069 5284
rect 10652 5244 10658 5256
rect 11057 5253 11069 5256
rect 11103 5284 11115 5287
rect 11790 5284 11796 5296
rect 11103 5256 11796 5284
rect 11103 5253 11115 5256
rect 11057 5247 11115 5253
rect 11790 5244 11796 5256
rect 11848 5244 11854 5296
rect 14461 5287 14519 5293
rect 14461 5284 14473 5287
rect 13556 5256 14473 5284
rect 6822 5176 6828 5228
rect 6880 5216 6886 5228
rect 7193 5219 7251 5225
rect 7193 5216 7205 5219
rect 6880 5188 7205 5216
rect 6880 5176 6886 5188
rect 7193 5185 7205 5188
rect 7239 5216 7251 5219
rect 8110 5216 8116 5228
rect 7239 5188 8116 5216
rect 7239 5185 7251 5188
rect 7193 5179 7251 5185
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 8478 5176 8484 5228
rect 8536 5216 8542 5228
rect 9401 5219 9459 5225
rect 9401 5216 9413 5219
rect 8536 5188 9413 5216
rect 8536 5176 8542 5188
rect 9401 5185 9413 5188
rect 9447 5216 9459 5219
rect 10502 5216 10508 5228
rect 9447 5188 10508 5216
rect 9447 5185 9459 5188
rect 9401 5179 9459 5185
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 10962 5176 10968 5228
rect 11020 5216 11026 5228
rect 11149 5219 11207 5225
rect 11149 5216 11161 5219
rect 11020 5188 11161 5216
rect 11020 5176 11026 5188
rect 11149 5185 11161 5188
rect 11195 5185 11207 5219
rect 11149 5179 11207 5185
rect 13449 5219 13507 5225
rect 13449 5185 13461 5219
rect 13495 5216 13507 5219
rect 13556 5216 13584 5256
rect 14461 5253 14473 5256
rect 14507 5284 14519 5287
rect 16850 5284 16856 5296
rect 14507 5256 16856 5284
rect 14507 5253 14519 5256
rect 14461 5247 14519 5253
rect 16850 5244 16856 5256
rect 16908 5244 16914 5296
rect 13495 5188 13584 5216
rect 13495 5185 13507 5188
rect 13449 5179 13507 5185
rect 13814 5176 13820 5228
rect 13872 5216 13878 5228
rect 13872 5188 13917 5216
rect 13872 5176 13878 5188
rect 16574 5176 16580 5228
rect 16632 5216 16638 5228
rect 16669 5219 16727 5225
rect 16669 5216 16681 5219
rect 16632 5188 16681 5216
rect 16632 5176 16638 5188
rect 16669 5185 16681 5188
rect 16715 5216 16727 5219
rect 16945 5219 17003 5225
rect 16945 5216 16957 5219
rect 16715 5188 16957 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 16945 5185 16957 5188
rect 16991 5185 17003 5219
rect 20162 5216 20168 5228
rect 20123 5188 20168 5216
rect 16945 5179 17003 5185
rect 20162 5176 20168 5188
rect 20220 5176 20226 5228
rect 20438 5216 20444 5228
rect 20399 5188 20444 5216
rect 20438 5176 20444 5188
rect 20496 5176 20502 5228
rect 5480 5151 5538 5157
rect 5480 5148 5492 5151
rect 5276 5120 5492 5148
rect 5480 5117 5492 5120
rect 5526 5117 5538 5151
rect 6270 5148 6276 5160
rect 5480 5111 5538 5117
rect 5920 5120 6276 5148
rect 4154 5040 4160 5092
rect 4212 5080 4218 5092
rect 4798 5080 4804 5092
rect 4212 5052 4804 5080
rect 4212 5040 4218 5052
rect 4798 5040 4804 5052
rect 4856 5080 4862 5092
rect 5920 5089 5948 5120
rect 6270 5108 6276 5120
rect 6328 5148 6334 5160
rect 6972 5151 7030 5157
rect 6972 5148 6984 5151
rect 6328 5120 6984 5148
rect 6328 5108 6334 5120
rect 6972 5117 6984 5120
rect 7018 5117 7030 5151
rect 6972 5111 7030 5117
rect 7742 5108 7748 5160
rect 7800 5148 7806 5160
rect 8573 5151 8631 5157
rect 8573 5148 8585 5151
rect 7800 5120 8585 5148
rect 7800 5108 7806 5120
rect 8128 5092 8156 5120
rect 8573 5117 8585 5120
rect 8619 5148 8631 5151
rect 9033 5151 9091 5157
rect 9033 5148 9045 5151
rect 8619 5120 9045 5148
rect 8619 5117 8631 5120
rect 8573 5111 8631 5117
rect 9033 5117 9045 5120
rect 9079 5148 9091 5151
rect 10781 5151 10839 5157
rect 10781 5148 10793 5151
rect 9079 5120 10793 5148
rect 9079 5117 9091 5120
rect 9033 5111 9091 5117
rect 10781 5117 10793 5120
rect 10827 5148 10839 5151
rect 11793 5151 11851 5157
rect 11793 5148 11805 5151
rect 10827 5120 11805 5148
rect 10827 5117 10839 5120
rect 10781 5111 10839 5117
rect 11793 5117 11805 5120
rect 11839 5117 11851 5151
rect 11793 5111 11851 5117
rect 15838 5108 15844 5160
rect 15896 5148 15902 5160
rect 16025 5151 16083 5157
rect 16025 5148 16037 5151
rect 15896 5120 16037 5148
rect 15896 5108 15902 5120
rect 16025 5117 16037 5120
rect 16071 5117 16083 5151
rect 16025 5111 16083 5117
rect 17865 5151 17923 5157
rect 17865 5117 17877 5151
rect 17911 5148 17923 5151
rect 18138 5148 18144 5160
rect 17911 5120 18144 5148
rect 17911 5117 17923 5120
rect 17865 5111 17923 5117
rect 18138 5108 18144 5120
rect 18196 5148 18202 5160
rect 18325 5151 18383 5157
rect 18325 5148 18337 5151
rect 18196 5120 18337 5148
rect 18196 5108 18202 5120
rect 18325 5117 18337 5120
rect 18371 5117 18383 5151
rect 18325 5111 18383 5117
rect 5905 5083 5963 5089
rect 5905 5080 5917 5083
rect 4856 5052 5917 5080
rect 4856 5040 4862 5052
rect 5905 5049 5917 5052
rect 5951 5049 5963 5083
rect 5905 5043 5963 5049
rect 5994 5040 6000 5092
rect 6052 5080 6058 5092
rect 6825 5083 6883 5089
rect 6825 5080 6837 5083
rect 6052 5052 6837 5080
rect 6052 5040 6058 5052
rect 6825 5049 6837 5052
rect 6871 5049 6883 5083
rect 6825 5043 6883 5049
rect 8110 5040 8116 5092
rect 8168 5040 8174 5092
rect 11514 5080 11520 5092
rect 11475 5052 11520 5080
rect 11514 5040 11520 5052
rect 11572 5040 11578 5092
rect 13446 5040 13452 5092
rect 13504 5080 13510 5092
rect 13541 5083 13599 5089
rect 13541 5080 13553 5083
rect 13504 5052 13553 5080
rect 13504 5040 13510 5052
rect 13541 5049 13553 5052
rect 13587 5049 13599 5083
rect 13541 5043 13599 5049
rect 18687 5083 18745 5089
rect 18687 5049 18699 5083
rect 18733 5080 18745 5083
rect 18782 5080 18788 5092
rect 18733 5052 18788 5080
rect 18733 5049 18745 5052
rect 18687 5043 18745 5049
rect 18782 5040 18788 5052
rect 18840 5040 18846 5092
rect 20257 5083 20315 5089
rect 20257 5049 20269 5083
rect 20303 5049 20315 5083
rect 20257 5043 20315 5049
rect 1949 5015 2007 5021
rect 1949 4981 1961 5015
rect 1995 5012 2007 5015
rect 2406 5012 2412 5024
rect 1995 4984 2412 5012
rect 1995 4981 2007 4984
rect 1949 4975 2007 4981
rect 2406 4972 2412 4984
rect 2464 4972 2470 5024
rect 3970 5012 3976 5024
rect 3931 4984 3976 5012
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 4982 5012 4988 5024
rect 4943 4984 4988 5012
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 5350 4972 5356 5024
rect 5408 5012 5414 5024
rect 5583 5015 5641 5021
rect 5583 5012 5595 5015
rect 5408 4984 5595 5012
rect 5408 4972 5414 4984
rect 5583 4981 5595 4984
rect 5629 4981 5641 5015
rect 5583 4975 5641 4981
rect 9490 4972 9496 5024
rect 9548 5012 9554 5024
rect 9677 5015 9735 5021
rect 9677 5012 9689 5015
rect 9548 4984 9689 5012
rect 9548 4972 9554 4984
rect 9677 4981 9689 4984
rect 9723 4981 9735 5015
rect 9677 4975 9735 4981
rect 9766 4972 9772 5024
rect 9824 5012 9830 5024
rect 10229 5015 10287 5021
rect 10229 5012 10241 5015
rect 9824 4984 10241 5012
rect 9824 4972 9830 4984
rect 10229 4981 10241 4984
rect 10275 5012 10287 5015
rect 10870 5012 10876 5024
rect 10275 4984 10876 5012
rect 10275 4981 10287 4984
rect 10229 4975 10287 4981
rect 10870 4972 10876 4984
rect 10928 4972 10934 5024
rect 12618 5012 12624 5024
rect 12579 4984 12624 5012
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 19245 5015 19303 5021
rect 19245 5012 19257 5015
rect 19155 4984 19257 5012
rect 19245 4981 19257 4984
rect 19291 5012 19303 5015
rect 19886 5012 19892 5024
rect 19291 4984 19892 5012
rect 19291 4981 19303 4984
rect 19245 4975 19303 4981
rect 19886 4972 19892 4984
rect 19944 5012 19950 5024
rect 20272 5012 20300 5043
rect 19944 4984 20300 5012
rect 19944 4972 19950 4984
rect 1104 4922 22816 4944
rect 1104 4870 8982 4922
rect 9034 4870 9046 4922
rect 9098 4870 9110 4922
rect 9162 4870 9174 4922
rect 9226 4870 16982 4922
rect 17034 4870 17046 4922
rect 17098 4870 17110 4922
rect 17162 4870 17174 4922
rect 17226 4870 22816 4922
rect 1104 4848 22816 4870
rect 2498 4768 2504 4820
rect 2556 4808 2562 4820
rect 3050 4808 3056 4820
rect 2556 4780 3056 4808
rect 2556 4768 2562 4780
rect 3050 4768 3056 4780
rect 3108 4808 3114 4820
rect 3881 4811 3939 4817
rect 3108 4780 3601 4808
rect 3108 4768 3114 4780
rect 2409 4743 2467 4749
rect 2409 4709 2421 4743
rect 2455 4740 2467 4743
rect 2958 4740 2964 4752
rect 2455 4712 2964 4740
rect 2455 4709 2467 4712
rect 2409 4703 2467 4709
rect 2958 4700 2964 4712
rect 3016 4700 3022 4752
rect 3573 4740 3601 4780
rect 3881 4777 3893 4811
rect 3927 4808 3939 4811
rect 4614 4808 4620 4820
rect 3927 4780 4620 4808
rect 3927 4777 3939 4780
rect 3881 4771 3939 4777
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 4982 4768 4988 4820
rect 5040 4808 5046 4820
rect 5994 4808 6000 4820
rect 5040 4780 6000 4808
rect 5040 4768 5046 4780
rect 5994 4768 6000 4780
rect 6052 4808 6058 4820
rect 6089 4811 6147 4817
rect 6089 4808 6101 4811
rect 6052 4780 6101 4808
rect 6052 4768 6058 4780
rect 6089 4777 6101 4780
rect 6135 4808 6147 4811
rect 7193 4811 7251 4817
rect 7193 4808 7205 4811
rect 6135 4780 7205 4808
rect 6135 4777 6147 4780
rect 6089 4771 6147 4777
rect 7193 4777 7205 4780
rect 7239 4777 7251 4811
rect 7193 4771 7251 4777
rect 7745 4811 7803 4817
rect 7745 4777 7757 4811
rect 7791 4808 7803 4811
rect 7834 4808 7840 4820
rect 7791 4780 7840 4808
rect 7791 4777 7803 4780
rect 7745 4771 7803 4777
rect 7834 4768 7840 4780
rect 7892 4768 7898 4820
rect 8478 4768 8484 4820
rect 8536 4808 8542 4820
rect 9033 4811 9091 4817
rect 9033 4808 9045 4811
rect 8536 4780 9045 4808
rect 8536 4768 8542 4780
rect 9033 4777 9045 4780
rect 9079 4777 9091 4811
rect 9033 4771 9091 4777
rect 10873 4811 10931 4817
rect 10873 4777 10885 4811
rect 10919 4808 10931 4811
rect 10962 4808 10968 4820
rect 10919 4780 10968 4808
rect 10919 4777 10931 4780
rect 10873 4771 10931 4777
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 11514 4768 11520 4820
rect 11572 4808 11578 4820
rect 14001 4811 14059 4817
rect 14001 4808 14013 4811
rect 11572 4780 14013 4808
rect 11572 4768 11578 4780
rect 14001 4777 14013 4780
rect 14047 4777 14059 4811
rect 14001 4771 14059 4777
rect 15470 4768 15476 4820
rect 15528 4808 15534 4820
rect 15657 4811 15715 4817
rect 15657 4808 15669 4811
rect 15528 4780 15669 4808
rect 15528 4768 15534 4780
rect 15657 4777 15669 4780
rect 15703 4777 15715 4811
rect 15657 4771 15715 4777
rect 16577 4811 16635 4817
rect 16577 4777 16589 4811
rect 16623 4808 16635 4811
rect 16666 4808 16672 4820
rect 16623 4780 16672 4808
rect 16623 4777 16635 4780
rect 16577 4771 16635 4777
rect 16666 4768 16672 4780
rect 16724 4768 16730 4820
rect 4246 4740 4252 4752
rect 3573 4712 4252 4740
rect 4246 4700 4252 4712
rect 4304 4740 4310 4752
rect 4386 4743 4444 4749
rect 4386 4740 4398 4743
rect 4304 4712 4398 4740
rect 4304 4700 4310 4712
rect 4386 4709 4398 4712
rect 4432 4709 4444 4743
rect 6822 4740 6828 4752
rect 6783 4712 6828 4740
rect 4386 4703 4444 4709
rect 6822 4700 6828 4712
rect 6880 4700 6886 4752
rect 11422 4700 11428 4752
rect 11480 4740 11486 4752
rect 11701 4743 11759 4749
rect 11701 4740 11713 4743
rect 11480 4712 11713 4740
rect 11480 4700 11486 4712
rect 11701 4709 11713 4712
rect 11747 4709 11759 4743
rect 12434 4740 12440 4752
rect 12395 4712 12440 4740
rect 11701 4703 11759 4709
rect 12434 4700 12440 4712
rect 12492 4700 12498 4752
rect 13262 4740 13268 4752
rect 13223 4712 13268 4740
rect 13262 4700 13268 4712
rect 13320 4700 13326 4752
rect 13814 4700 13820 4752
rect 13872 4740 13878 4752
rect 18138 4740 18144 4752
rect 13872 4712 13917 4740
rect 18099 4712 18144 4740
rect 13872 4700 13878 4712
rect 18138 4700 18144 4712
rect 18196 4700 18202 4752
rect 20806 4700 20812 4752
rect 20864 4740 20870 4752
rect 21085 4743 21143 4749
rect 21085 4740 21097 4743
rect 20864 4712 21097 4740
rect 20864 4700 20870 4712
rect 21085 4709 21097 4712
rect 21131 4709 21143 4743
rect 21085 4703 21143 4709
rect 5810 4632 5816 4684
rect 5868 4672 5874 4684
rect 5905 4675 5963 4681
rect 5905 4672 5917 4675
rect 5868 4644 5917 4672
rect 5868 4632 5874 4644
rect 5905 4641 5917 4644
rect 5951 4641 5963 4675
rect 5905 4635 5963 4641
rect 7650 4632 7656 4684
rect 7708 4672 7714 4684
rect 9674 4672 9680 4684
rect 7708 4644 9680 4672
rect 7708 4632 7714 4644
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 10137 4675 10195 4681
rect 10137 4672 10149 4675
rect 9784 4644 10149 4672
rect 2314 4604 2320 4616
rect 2275 4576 2320 4604
rect 2314 4564 2320 4576
rect 2372 4564 2378 4616
rect 2498 4564 2504 4616
rect 2556 4604 2562 4616
rect 2593 4607 2651 4613
rect 2593 4604 2605 4607
rect 2556 4576 2605 4604
rect 2556 4564 2562 4576
rect 2593 4573 2605 4576
rect 2639 4573 2651 4607
rect 2593 4567 2651 4573
rect 3970 4564 3976 4616
rect 4028 4604 4034 4616
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 4028 4576 4077 4604
rect 4028 4564 4034 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 8665 4607 8723 4613
rect 8665 4573 8677 4607
rect 8711 4604 8723 4607
rect 9490 4604 9496 4616
rect 8711 4576 9496 4604
rect 8711 4573 8723 4576
rect 8665 4567 8723 4573
rect 9490 4564 9496 4576
rect 9548 4604 9554 4616
rect 9784 4604 9812 4644
rect 10137 4641 10149 4644
rect 10183 4672 10195 4675
rect 11330 4672 11336 4684
rect 10183 4644 11336 4672
rect 10183 4641 10195 4644
rect 10137 4635 10195 4641
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 17494 4672 17500 4684
rect 17455 4644 17500 4672
rect 17494 4632 17500 4644
rect 17552 4632 17558 4684
rect 17862 4672 17868 4684
rect 17823 4644 17868 4672
rect 17862 4632 17868 4644
rect 17920 4632 17926 4684
rect 19848 4675 19906 4681
rect 19848 4641 19860 4675
rect 19894 4672 19906 4675
rect 20070 4672 20076 4684
rect 19894 4644 20076 4672
rect 19894 4641 19906 4644
rect 19848 4635 19906 4641
rect 20070 4632 20076 4644
rect 20128 4632 20134 4684
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 9548 4576 9812 4604
rect 10152 4576 10241 4604
rect 9548 4564 9554 4576
rect 10152 4548 10180 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 11238 4604 11244 4616
rect 11199 4576 11244 4604
rect 10229 4567 10287 4573
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 12802 4564 12808 4616
rect 12860 4604 12866 4616
rect 13173 4607 13231 4613
rect 13173 4604 13185 4607
rect 12860 4576 13185 4604
rect 12860 4564 12866 4576
rect 13173 4573 13185 4576
rect 13219 4573 13231 4607
rect 15286 4604 15292 4616
rect 15247 4576 15292 4604
rect 13173 4567 13231 4573
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 19935 4607 19993 4613
rect 19935 4573 19947 4607
rect 19981 4604 19993 4607
rect 20993 4607 21051 4613
rect 20993 4604 21005 4607
rect 19981 4576 21005 4604
rect 19981 4573 19993 4576
rect 19935 4567 19993 4573
rect 20993 4573 21005 4576
rect 21039 4604 21051 4607
rect 21266 4604 21272 4616
rect 21039 4576 21272 4604
rect 21039 4573 21051 4576
rect 20993 4567 21051 4573
rect 21266 4564 21272 4576
rect 21324 4564 21330 4616
rect 10134 4496 10140 4548
rect 10192 4496 10198 4548
rect 20438 4496 20444 4548
rect 20496 4536 20502 4548
rect 21545 4539 21603 4545
rect 21545 4536 21557 4539
rect 20496 4508 21557 4536
rect 20496 4496 20502 4508
rect 21545 4505 21557 4508
rect 21591 4505 21603 4539
rect 21545 4499 21603 4505
rect 1854 4468 1860 4480
rect 1815 4440 1860 4468
rect 1854 4428 1860 4440
rect 1912 4428 1918 4480
rect 3786 4428 3792 4480
rect 3844 4468 3850 4480
rect 4985 4471 5043 4477
rect 4985 4468 4997 4471
rect 3844 4440 4997 4468
rect 3844 4428 3850 4440
rect 4985 4437 4997 4440
rect 5031 4437 5043 4471
rect 4985 4431 5043 4437
rect 14001 4471 14059 4477
rect 14001 4437 14013 4471
rect 14047 4468 14059 4471
rect 14185 4471 14243 4477
rect 14185 4468 14197 4471
rect 14047 4440 14197 4468
rect 14047 4437 14059 4440
rect 14001 4431 14059 4437
rect 14185 4437 14197 4440
rect 14231 4468 14243 4471
rect 14458 4468 14464 4480
rect 14231 4440 14464 4468
rect 14231 4437 14243 4440
rect 14185 4431 14243 4437
rect 14458 4428 14464 4440
rect 14516 4428 14522 4480
rect 16206 4468 16212 4480
rect 16167 4440 16212 4468
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 1104 4378 22816 4400
rect 1104 4326 4982 4378
rect 5034 4326 5046 4378
rect 5098 4326 5110 4378
rect 5162 4326 5174 4378
rect 5226 4326 12982 4378
rect 13034 4326 13046 4378
rect 13098 4326 13110 4378
rect 13162 4326 13174 4378
rect 13226 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 22816 4378
rect 1104 4304 22816 4326
rect 1673 4267 1731 4273
rect 1673 4233 1685 4267
rect 1719 4264 1731 4267
rect 1762 4264 1768 4276
rect 1719 4236 1768 4264
rect 1719 4233 1731 4236
rect 1673 4227 1731 4233
rect 1688 3924 1716 4227
rect 1762 4224 1768 4236
rect 1820 4224 1826 4276
rect 2314 4224 2320 4276
rect 2372 4264 2378 4276
rect 2372 4236 4154 4264
rect 2372 4224 2378 4236
rect 2869 4199 2927 4205
rect 2869 4165 2881 4199
rect 2915 4196 2927 4199
rect 2958 4196 2964 4208
rect 2915 4168 2964 4196
rect 2915 4165 2927 4168
rect 2869 4159 2927 4165
rect 2958 4156 2964 4168
rect 3016 4156 3022 4208
rect 4126 4196 4154 4236
rect 4246 4224 4252 4276
rect 4304 4264 4310 4276
rect 4985 4267 5043 4273
rect 4985 4264 4997 4267
rect 4304 4236 4997 4264
rect 4304 4224 4310 4236
rect 4985 4233 4997 4236
rect 5031 4264 5043 4267
rect 8018 4264 8024 4276
rect 5031 4236 8024 4264
rect 5031 4233 5043 4236
rect 4985 4227 5043 4233
rect 8018 4224 8024 4236
rect 8076 4224 8082 4276
rect 9674 4264 9680 4276
rect 9635 4236 9680 4264
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 11330 4264 11336 4276
rect 11291 4236 11336 4264
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 12802 4264 12808 4276
rect 12763 4236 12808 4264
rect 12802 4224 12808 4236
rect 12860 4264 12866 4276
rect 15286 4264 15292 4276
rect 12860 4236 12940 4264
rect 15199 4236 15292 4264
rect 12860 4224 12866 4236
rect 4525 4199 4583 4205
rect 4525 4196 4537 4199
rect 4126 4168 4537 4196
rect 4525 4165 4537 4168
rect 4571 4196 4583 4199
rect 4798 4196 4804 4208
rect 4571 4168 4804 4196
rect 4571 4165 4583 4168
rect 4525 4159 4583 4165
rect 4798 4156 4804 4168
rect 4856 4156 4862 4208
rect 7926 4156 7932 4208
rect 7984 4196 7990 4208
rect 8389 4199 8447 4205
rect 8389 4196 8401 4199
rect 7984 4168 8401 4196
rect 7984 4156 7990 4168
rect 8389 4165 8401 4168
rect 8435 4165 8447 4199
rect 8389 4159 8447 4165
rect 2498 4128 2504 4140
rect 2459 4100 2504 4128
rect 2498 4088 2504 4100
rect 2556 4088 2562 4140
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4128 3479 4131
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3467 4100 3985 4128
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 3973 4097 3985 4100
rect 4019 4128 4031 4131
rect 5350 4128 5356 4140
rect 4019 4100 5356 4128
rect 4019 4097 4031 4100
rect 3973 4091 4031 4097
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5902 4020 5908 4072
rect 5960 4060 5966 4072
rect 6860 4063 6918 4069
rect 6860 4060 6872 4063
rect 5960 4032 6872 4060
rect 5960 4020 5966 4032
rect 6860 4029 6872 4032
rect 6906 4060 6918 4063
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 6906 4032 7297 4060
rect 6906 4029 6918 4032
rect 6860 4023 6918 4029
rect 7285 4029 7297 4032
rect 7331 4029 7343 4063
rect 8404 4060 8432 4159
rect 12912 4137 12940 4236
rect 15286 4224 15292 4236
rect 15344 4264 15350 4276
rect 17037 4267 17095 4273
rect 17037 4264 17049 4267
rect 15344 4236 17049 4264
rect 15344 4224 15350 4236
rect 17037 4233 17049 4236
rect 17083 4233 17095 4267
rect 17037 4227 17095 4233
rect 19705 4267 19763 4273
rect 19705 4233 19717 4267
rect 19751 4264 19763 4267
rect 20070 4264 20076 4276
rect 19751 4236 20076 4264
rect 19751 4233 19763 4236
rect 19705 4227 19763 4233
rect 20070 4224 20076 4236
rect 20128 4224 20134 4276
rect 21266 4264 21272 4276
rect 21227 4236 21272 4264
rect 21266 4224 21272 4236
rect 21324 4224 21330 4276
rect 13262 4156 13268 4208
rect 13320 4196 13326 4208
rect 13357 4199 13415 4205
rect 13357 4196 13369 4199
rect 13320 4168 13369 4196
rect 13320 4156 13326 4168
rect 13357 4165 13369 4168
rect 13403 4165 13415 4199
rect 13357 4159 13415 4165
rect 12897 4131 12955 4137
rect 12897 4097 12909 4131
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 14737 4131 14795 4137
rect 14737 4097 14749 4131
rect 14783 4128 14795 4131
rect 15304 4128 15332 4224
rect 17773 4199 17831 4205
rect 17773 4196 17785 4199
rect 14783 4100 15332 4128
rect 15396 4168 17785 4196
rect 14783 4097 14795 4100
rect 14737 4091 14795 4097
rect 8573 4063 8631 4069
rect 8573 4060 8585 4063
rect 8404 4032 8585 4060
rect 7285 4023 7343 4029
rect 8573 4029 8585 4032
rect 8619 4029 8631 4063
rect 8573 4023 8631 4029
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4060 9183 4063
rect 9490 4060 9496 4072
rect 9171 4032 9496 4060
rect 9171 4029 9183 4032
rect 9125 4023 9183 4029
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 10134 4060 10140 4072
rect 10095 4032 10140 4060
rect 10134 4020 10140 4032
rect 10192 4020 10198 4072
rect 12526 4020 12532 4072
rect 12584 4060 12590 4072
rect 13909 4063 13967 4069
rect 13909 4060 13921 4063
rect 12584 4032 13921 4060
rect 12584 4020 12590 4032
rect 13909 4029 13921 4032
rect 13955 4060 13967 4063
rect 14001 4063 14059 4069
rect 14001 4060 14013 4063
rect 13955 4032 14013 4060
rect 13955 4029 13967 4032
rect 13909 4023 13967 4029
rect 14001 4029 14013 4032
rect 14047 4029 14059 4063
rect 14458 4060 14464 4072
rect 14419 4032 14464 4060
rect 14001 4023 14059 4029
rect 14458 4020 14464 4032
rect 14516 4060 14522 4072
rect 15396 4060 15424 4168
rect 17773 4165 17785 4168
rect 17819 4196 17831 4199
rect 17862 4196 17868 4208
rect 17819 4168 17868 4196
rect 17819 4165 17831 4168
rect 17773 4159 17831 4165
rect 17862 4156 17868 4168
rect 17920 4156 17926 4208
rect 16482 4128 16488 4140
rect 16443 4100 16488 4128
rect 16482 4088 16488 4100
rect 16540 4088 16546 4140
rect 19886 4060 19892 4072
rect 14516 4032 15424 4060
rect 19847 4032 19892 4060
rect 14516 4020 14522 4032
rect 19886 4020 19892 4032
rect 19944 4020 19950 4072
rect 1854 3992 1860 4004
rect 1815 3964 1860 3992
rect 1854 3952 1860 3964
rect 1912 3952 1918 4004
rect 1949 3995 2007 4001
rect 1949 3961 1961 3995
rect 1995 3961 2007 3995
rect 3786 3992 3792 4004
rect 3747 3964 3792 3992
rect 1949 3955 2007 3961
rect 1964 3924 1992 3955
rect 3786 3952 3792 3964
rect 3844 3952 3850 4004
rect 4074 3995 4132 4001
rect 4074 3961 4086 3995
rect 4120 3992 4132 3995
rect 9306 3992 9312 4004
rect 4120 3961 4154 3992
rect 9267 3964 9312 3992
rect 4074 3955 4154 3961
rect 1688 3896 1992 3924
rect 3804 3924 3832 3952
rect 4126 3924 4154 3955
rect 9306 3952 9312 3964
rect 9364 3952 9370 4004
rect 10042 3992 10048 4004
rect 9955 3964 10048 3992
rect 10042 3952 10048 3964
rect 10100 3992 10106 4004
rect 10499 3995 10557 4001
rect 10499 3992 10511 3995
rect 10100 3964 10511 3992
rect 10100 3952 10106 3964
rect 10499 3961 10511 3964
rect 10545 3992 10557 3995
rect 12618 3992 12624 4004
rect 10545 3964 12624 3992
rect 10545 3961 10557 3964
rect 10499 3955 10557 3961
rect 12618 3952 12624 3964
rect 12676 3992 12682 4004
rect 15289 3995 15347 4001
rect 15289 3992 15301 3995
rect 12676 3964 15301 3992
rect 12676 3952 12682 3964
rect 15289 3961 15301 3964
rect 15335 3992 15347 3995
rect 15470 3992 15476 4004
rect 15335 3964 15476 3992
rect 15335 3961 15347 3964
rect 15289 3955 15347 3961
rect 15470 3952 15476 3964
rect 15528 3952 15534 4004
rect 16114 3992 16120 4004
rect 16075 3964 16120 3992
rect 16114 3952 16120 3964
rect 16172 3952 16178 4004
rect 16206 3952 16212 4004
rect 16264 3992 16270 4004
rect 20533 3995 20591 4001
rect 16264 3964 16309 3992
rect 16264 3952 16270 3964
rect 20533 3961 20545 3995
rect 20579 3992 20591 3995
rect 20806 3992 20812 4004
rect 20579 3964 20812 3992
rect 20579 3961 20591 3964
rect 20533 3955 20591 3961
rect 20806 3952 20812 3964
rect 20864 3992 20870 4004
rect 20901 3995 20959 4001
rect 20901 3992 20913 3995
rect 20864 3964 20913 3992
rect 20864 3952 20870 3964
rect 20901 3961 20913 3964
rect 20947 3961 20959 3995
rect 20901 3955 20959 3961
rect 5810 3924 5816 3936
rect 3804 3896 4154 3924
rect 5771 3896 5816 3924
rect 5810 3884 5816 3896
rect 5868 3884 5874 3936
rect 6963 3927 7021 3933
rect 6963 3893 6975 3927
rect 7009 3924 7021 3927
rect 8294 3924 8300 3936
rect 7009 3896 8300 3924
rect 7009 3893 7021 3896
rect 6963 3887 7021 3893
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 11057 3927 11115 3933
rect 11057 3893 11069 3927
rect 11103 3924 11115 3927
rect 11606 3924 11612 3936
rect 11103 3896 11612 3924
rect 11103 3893 11115 3896
rect 11057 3887 11115 3893
rect 11606 3884 11612 3896
rect 11664 3884 11670 3936
rect 15933 3927 15991 3933
rect 15933 3893 15945 3927
rect 15979 3924 15991 3927
rect 16224 3924 16252 3952
rect 17494 3924 17500 3936
rect 15979 3896 16252 3924
rect 17455 3896 17500 3924
rect 15979 3893 15991 3896
rect 15933 3887 15991 3893
rect 17494 3884 17500 3896
rect 17552 3884 17558 3936
rect 1104 3834 22816 3856
rect 1104 3782 8982 3834
rect 9034 3782 9046 3834
rect 9098 3782 9110 3834
rect 9162 3782 9174 3834
rect 9226 3782 16982 3834
rect 17034 3782 17046 3834
rect 17098 3782 17110 3834
rect 17162 3782 17174 3834
rect 17226 3782 22816 3834
rect 1104 3760 22816 3782
rect 106 3680 112 3732
rect 164 3720 170 3732
rect 1581 3723 1639 3729
rect 1581 3720 1593 3723
rect 164 3692 1593 3720
rect 164 3680 170 3692
rect 1581 3689 1593 3692
rect 1627 3689 1639 3723
rect 2314 3720 2320 3732
rect 2275 3692 2320 3720
rect 1581 3683 1639 3689
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 4249 3723 4307 3729
rect 4249 3720 4261 3723
rect 4028 3692 4261 3720
rect 4028 3680 4034 3692
rect 4249 3689 4261 3692
rect 4295 3689 4307 3723
rect 8386 3720 8392 3732
rect 8347 3692 8392 3720
rect 4249 3683 4307 3689
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 9306 3680 9312 3732
rect 9364 3720 9370 3732
rect 9401 3723 9459 3729
rect 9401 3720 9413 3723
rect 9364 3692 9413 3720
rect 9364 3680 9370 3692
rect 9401 3689 9413 3692
rect 9447 3689 9459 3723
rect 10042 3720 10048 3732
rect 10003 3692 10048 3720
rect 9401 3683 9459 3689
rect 1854 3612 1860 3664
rect 1912 3652 1918 3664
rect 2501 3655 2559 3661
rect 2501 3652 2513 3655
rect 1912 3624 2513 3652
rect 1912 3612 1918 3624
rect 2501 3621 2513 3624
rect 2547 3621 2559 3655
rect 4614 3652 4620 3664
rect 4575 3624 4620 3652
rect 2501 3615 2559 3621
rect 4614 3612 4620 3624
rect 4672 3612 4678 3664
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3584 1455 3587
rect 2314 3584 2320 3596
rect 1443 3556 2320 3584
rect 1443 3553 1455 3556
rect 1397 3547 1455 3553
rect 2314 3544 2320 3556
rect 2372 3544 2378 3596
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 7044 3587 7102 3593
rect 7044 3584 7056 3587
rect 6972 3556 7056 3584
rect 6972 3544 6978 3556
rect 7044 3553 7056 3556
rect 7090 3553 7102 3587
rect 7044 3547 7102 3553
rect 8272 3587 8330 3593
rect 8272 3553 8284 3587
rect 8318 3584 8330 3587
rect 8478 3584 8484 3596
rect 8318 3556 8484 3584
rect 8318 3553 8330 3556
rect 8272 3547 8330 3553
rect 8478 3544 8484 3556
rect 8536 3544 8542 3596
rect 9416 3584 9444 3683
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 10134 3680 10140 3732
rect 10192 3720 10198 3732
rect 10873 3723 10931 3729
rect 10873 3720 10885 3723
rect 10192 3692 10885 3720
rect 10192 3680 10198 3692
rect 10873 3689 10885 3692
rect 10919 3689 10931 3723
rect 10873 3683 10931 3689
rect 11238 3680 11244 3732
rect 11296 3720 11302 3732
rect 12437 3723 12495 3729
rect 12437 3720 12449 3723
rect 11296 3692 12449 3720
rect 11296 3680 11302 3692
rect 12437 3689 12449 3692
rect 12483 3720 12495 3723
rect 12526 3720 12532 3732
rect 12483 3692 12532 3720
rect 12483 3689 12495 3692
rect 12437 3683 12495 3689
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 15657 3723 15715 3729
rect 15657 3689 15669 3723
rect 15703 3720 15715 3723
rect 16206 3720 16212 3732
rect 15703 3692 16212 3720
rect 15703 3689 15715 3692
rect 15657 3683 15715 3689
rect 16206 3680 16212 3692
rect 16264 3680 16270 3732
rect 19886 3720 19892 3732
rect 19847 3692 19892 3720
rect 19886 3680 19892 3692
rect 19944 3680 19950 3732
rect 11606 3652 11612 3664
rect 11567 3624 11612 3652
rect 11606 3612 11612 3624
rect 11664 3612 11670 3664
rect 11698 3612 11704 3664
rect 11756 3652 11762 3664
rect 15930 3652 15936 3664
rect 11756 3624 13032 3652
rect 15891 3624 15936 3652
rect 11756 3612 11762 3624
rect 13004 3593 13032 3624
rect 15930 3612 15936 3624
rect 15988 3612 15994 3664
rect 16114 3612 16120 3664
rect 16172 3652 16178 3664
rect 16853 3655 16911 3661
rect 16853 3652 16865 3655
rect 16172 3624 16865 3652
rect 16172 3612 16178 3624
rect 16853 3621 16865 3624
rect 16899 3652 16911 3655
rect 20438 3652 20444 3664
rect 16899 3624 20444 3652
rect 16899 3621 16911 3624
rect 16853 3615 16911 3621
rect 20438 3612 20444 3624
rect 20496 3612 20502 3664
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 9416 3556 9689 3584
rect 9677 3553 9689 3556
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 12989 3587 13047 3593
rect 12989 3553 13001 3587
rect 13035 3584 13047 3587
rect 13446 3584 13452 3596
rect 13035 3556 13452 3584
rect 13035 3553 13047 3556
rect 12989 3547 13047 3553
rect 13446 3544 13452 3556
rect 13504 3544 13510 3596
rect 13814 3544 13820 3596
rect 13872 3584 13878 3596
rect 14128 3587 14186 3593
rect 14128 3584 14140 3587
rect 13872 3556 14140 3584
rect 13872 3544 13878 3556
rect 14128 3553 14140 3556
rect 14174 3553 14186 3587
rect 14128 3547 14186 3553
rect 16482 3544 16488 3596
rect 16540 3584 16546 3596
rect 16540 3556 16585 3584
rect 16540 3544 16546 3556
rect 4522 3516 4528 3528
rect 4483 3488 4528 3516
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 4798 3516 4804 3528
rect 4759 3488 4804 3516
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 10962 3476 10968 3528
rect 11020 3516 11026 3528
rect 11517 3519 11575 3525
rect 11517 3516 11529 3519
rect 11020 3488 11529 3516
rect 11020 3476 11026 3488
rect 11517 3485 11529 3488
rect 11563 3485 11575 3519
rect 11517 3479 11575 3485
rect 12161 3519 12219 3525
rect 12161 3485 12173 3519
rect 12207 3516 12219 3519
rect 12802 3516 12808 3528
rect 12207 3488 12808 3516
rect 12207 3485 12219 3488
rect 12161 3479 12219 3485
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 15470 3476 15476 3528
rect 15528 3516 15534 3528
rect 15841 3519 15899 3525
rect 15841 3516 15853 3519
rect 15528 3488 15853 3516
rect 15528 3476 15534 3488
rect 15841 3485 15853 3488
rect 15887 3516 15899 3519
rect 17313 3519 17371 3525
rect 17313 3516 17325 3519
rect 15887 3488 17325 3516
rect 15887 3485 15899 3488
rect 15841 3479 15899 3485
rect 17313 3485 17325 3488
rect 17359 3485 17371 3519
rect 17313 3479 17371 3485
rect 6822 3380 6828 3392
rect 6783 3352 6828 3380
rect 6822 3340 6828 3352
rect 6880 3340 6886 3392
rect 7147 3383 7205 3389
rect 7147 3349 7159 3383
rect 7193 3380 7205 3383
rect 9858 3380 9864 3392
rect 7193 3352 9864 3380
rect 7193 3349 7205 3352
rect 7147 3343 7205 3349
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 10410 3340 10416 3392
rect 10468 3380 10474 3392
rect 10597 3383 10655 3389
rect 10597 3380 10609 3383
rect 10468 3352 10609 3380
rect 10468 3340 10474 3352
rect 10597 3349 10609 3352
rect 10643 3349 10655 3383
rect 10597 3343 10655 3349
rect 11790 3340 11796 3392
rect 11848 3380 11854 3392
rect 13173 3383 13231 3389
rect 13173 3380 13185 3383
rect 11848 3352 13185 3380
rect 11848 3340 11854 3352
rect 13173 3349 13185 3352
rect 13219 3349 13231 3383
rect 13173 3343 13231 3349
rect 13354 3340 13360 3392
rect 13412 3380 13418 3392
rect 14231 3383 14289 3389
rect 14231 3380 14243 3383
rect 13412 3352 14243 3380
rect 13412 3340 13418 3352
rect 14231 3349 14243 3352
rect 14277 3349 14289 3383
rect 14231 3343 14289 3349
rect 1104 3290 22816 3312
rect 1104 3238 4982 3290
rect 5034 3238 5046 3290
rect 5098 3238 5110 3290
rect 5162 3238 5174 3290
rect 5226 3238 12982 3290
rect 13034 3238 13046 3290
rect 13098 3238 13110 3290
rect 13162 3238 13174 3290
rect 13226 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 22816 3290
rect 1104 3216 22816 3238
rect 1394 3136 1400 3188
rect 1452 3176 1458 3188
rect 2547 3179 2605 3185
rect 2547 3176 2559 3179
rect 1452 3148 2559 3176
rect 1452 3136 1458 3148
rect 2547 3145 2559 3148
rect 2593 3145 2605 3179
rect 2547 3139 2605 3145
rect 3786 3136 3792 3188
rect 3844 3176 3850 3188
rect 4065 3179 4123 3185
rect 4065 3176 4077 3179
rect 3844 3148 4077 3176
rect 3844 3136 3850 3148
rect 4065 3145 4077 3148
rect 4111 3145 4123 3179
rect 10042 3176 10048 3188
rect 10003 3148 10048 3176
rect 4065 3139 4123 3145
rect 106 3000 112 3052
rect 164 3040 170 3052
rect 2314 3040 2320 3052
rect 164 3012 1507 3040
rect 2275 3012 2320 3040
rect 164 3000 170 3012
rect 1479 2981 1507 3012
rect 2314 3000 2320 3012
rect 2372 3000 2378 3052
rect 2498 2981 2504 2984
rect 1464 2975 1522 2981
rect 1464 2941 1476 2975
rect 1510 2972 1522 2975
rect 1857 2975 1915 2981
rect 1857 2972 1869 2975
rect 1510 2944 1869 2972
rect 1510 2941 1522 2944
rect 1464 2935 1522 2941
rect 1857 2941 1869 2944
rect 1903 2941 1915 2975
rect 2476 2975 2504 2981
rect 2476 2972 2488 2975
rect 2411 2944 2488 2972
rect 1857 2935 1915 2941
rect 2476 2941 2488 2944
rect 2556 2972 2562 2984
rect 2869 2975 2927 2981
rect 2869 2972 2881 2975
rect 2556 2944 2881 2972
rect 2476 2935 2504 2941
rect 2498 2932 2504 2935
rect 2556 2932 2562 2944
rect 2869 2941 2881 2944
rect 2915 2941 2927 2975
rect 4080 2972 4108 3139
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 10410 3176 10416 3188
rect 10371 3148 10416 3176
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 13446 3176 13452 3188
rect 13407 3148 13452 3176
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 14093 3179 14151 3185
rect 14093 3176 14105 3179
rect 13872 3148 14105 3176
rect 13872 3136 13878 3148
rect 14093 3145 14105 3148
rect 14139 3145 14151 3179
rect 15470 3176 15476 3188
rect 15431 3148 15476 3176
rect 14093 3139 14151 3145
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 11146 3108 11152 3120
rect 5368 3080 11152 3108
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4672 3012 4997 3040
rect 4672 3000 4678 3012
rect 4985 3009 4997 3012
rect 5031 3040 5043 3043
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 5031 3012 5273 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5261 3009 5273 3012
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 4341 2975 4399 2981
rect 4341 2972 4353 2975
rect 4080 2944 4353 2972
rect 2869 2935 2927 2941
rect 4341 2941 4353 2944
rect 4387 2941 4399 2975
rect 4341 2935 4399 2941
rect 1673 2907 1731 2913
rect 1673 2873 1685 2907
rect 1719 2904 1731 2907
rect 5368 2904 5396 3080
rect 11146 3068 11152 3080
rect 11204 3068 11210 3120
rect 15105 3111 15163 3117
rect 15105 3077 15117 3111
rect 15151 3108 15163 3111
rect 16482 3108 16488 3120
rect 15151 3080 16488 3108
rect 15151 3077 15163 3080
rect 15105 3071 15163 3077
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3040 7435 3043
rect 8110 3040 8116 3052
rect 7423 3012 8116 3040
rect 7423 3009 7435 3012
rect 7377 3003 7435 3009
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 10226 3000 10232 3052
rect 10284 3040 10290 3052
rect 10597 3043 10655 3049
rect 10597 3040 10609 3043
rect 10284 3012 10609 3040
rect 10284 3000 10290 3012
rect 10597 3009 10609 3012
rect 10643 3040 10655 3043
rect 10686 3040 10692 3052
rect 10643 3012 10692 3040
rect 10643 3009 10655 3012
rect 10597 3003 10655 3009
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 10962 3040 10968 3052
rect 10923 3012 10968 3040
rect 10962 3000 10968 3012
rect 11020 3000 11026 3052
rect 12526 3040 12532 3052
rect 12487 3012 12532 3040
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 12802 3040 12808 3052
rect 12763 3012 12808 3040
rect 12802 3000 12808 3012
rect 12860 3000 12866 3052
rect 7009 2975 7067 2981
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 8849 2975 8907 2981
rect 7055 2944 7788 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 1719 2876 5396 2904
rect 1719 2873 1731 2876
rect 1673 2867 1731 2873
rect 5994 2864 6000 2916
rect 6052 2904 6058 2916
rect 6822 2904 6828 2916
rect 6052 2876 6828 2904
rect 6052 2864 6058 2876
rect 6822 2864 6828 2876
rect 6880 2864 6886 2916
rect 7760 2848 7788 2944
rect 8849 2941 8861 2975
rect 8895 2972 8907 2975
rect 9585 2975 9643 2981
rect 9585 2972 9597 2975
rect 8895 2944 9597 2972
rect 8895 2941 8907 2944
rect 8849 2935 8907 2941
rect 9585 2941 9597 2944
rect 9631 2941 9643 2975
rect 9585 2935 9643 2941
rect 14604 2975 14662 2981
rect 14604 2941 14616 2975
rect 14650 2972 14662 2975
rect 15120 2972 15148 3071
rect 16482 3068 16488 3080
rect 16540 3068 16546 3120
rect 15930 3000 15936 3052
rect 15988 3040 15994 3052
rect 16301 3043 16359 3049
rect 16301 3040 16313 3043
rect 15988 3012 16313 3040
rect 15988 3000 15994 3012
rect 16301 3009 16313 3012
rect 16347 3040 16359 3043
rect 16577 3043 16635 3049
rect 16577 3040 16589 3043
rect 16347 3012 16589 3040
rect 16347 3009 16359 3012
rect 16301 3003 16359 3009
rect 16577 3009 16589 3012
rect 16623 3009 16635 3043
rect 16577 3003 16635 3009
rect 16206 2972 16212 2984
rect 14650 2944 15148 2972
rect 16167 2944 16212 2972
rect 14650 2941 14662 2944
rect 14604 2935 14662 2941
rect 9600 2904 9628 2935
rect 16206 2932 16212 2944
rect 16264 2932 16270 2984
rect 18392 2975 18450 2981
rect 18392 2941 18404 2975
rect 18438 2972 18450 2975
rect 18438 2944 18920 2972
rect 18438 2941 18450 2944
rect 18392 2935 18450 2941
rect 10410 2904 10416 2916
rect 9600 2876 10416 2904
rect 10410 2864 10416 2876
rect 10468 2904 10474 2916
rect 10689 2907 10747 2913
rect 10689 2904 10701 2907
rect 10468 2876 10701 2904
rect 10468 2864 10474 2876
rect 10689 2873 10701 2876
rect 10735 2873 10747 2907
rect 10689 2867 10747 2873
rect 12618 2864 12624 2916
rect 12676 2904 12682 2916
rect 14691 2907 14749 2913
rect 12676 2876 12721 2904
rect 12676 2864 12682 2876
rect 14691 2873 14703 2907
rect 14737 2904 14749 2907
rect 16574 2904 16580 2916
rect 14737 2876 16580 2904
rect 14737 2873 14749 2876
rect 14691 2867 14749 2873
rect 16574 2864 16580 2876
rect 16632 2864 16638 2916
rect 6641 2839 6699 2845
rect 6641 2805 6653 2839
rect 6687 2836 6699 2839
rect 6914 2836 6920 2848
rect 6687 2808 6920 2836
rect 6687 2805 6699 2808
rect 6641 2799 6699 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7742 2836 7748 2848
rect 7703 2808 7748 2836
rect 7742 2796 7748 2808
rect 7800 2796 7806 2848
rect 8297 2839 8355 2845
rect 8297 2805 8309 2839
rect 8343 2836 8355 2839
rect 8478 2836 8484 2848
rect 8343 2808 8484 2836
rect 8343 2805 8355 2808
rect 8297 2799 8355 2805
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 9398 2836 9404 2848
rect 9359 2808 9404 2836
rect 9398 2796 9404 2808
rect 9456 2796 9462 2848
rect 11606 2836 11612 2848
rect 11567 2808 11612 2836
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 12253 2839 12311 2845
rect 12253 2805 12265 2839
rect 12299 2836 12311 2839
rect 12636 2836 12664 2864
rect 12299 2808 12664 2836
rect 12299 2805 12311 2808
rect 12253 2799 12311 2805
rect 16022 2796 16028 2848
rect 16080 2836 16086 2848
rect 18892 2845 18920 2944
rect 18463 2839 18521 2845
rect 18463 2836 18475 2839
rect 16080 2808 18475 2836
rect 16080 2796 16086 2808
rect 18463 2805 18475 2808
rect 18509 2805 18521 2839
rect 18463 2799 18521 2805
rect 18877 2839 18935 2845
rect 18877 2805 18889 2839
rect 18923 2836 18935 2839
rect 19518 2836 19524 2848
rect 18923 2808 19524 2836
rect 18923 2805 18935 2808
rect 18877 2799 18935 2805
rect 19518 2796 19524 2808
rect 19576 2796 19582 2848
rect 1104 2746 22816 2768
rect 1104 2694 8982 2746
rect 9034 2694 9046 2746
rect 9098 2694 9110 2746
rect 9162 2694 9174 2746
rect 9226 2694 16982 2746
rect 17034 2694 17046 2746
rect 17098 2694 17110 2746
rect 17162 2694 17174 2746
rect 17226 2694 22816 2746
rect 1104 2672 22816 2694
rect 1535 2635 1593 2641
rect 1535 2601 1547 2635
rect 1581 2632 1593 2635
rect 2222 2632 2228 2644
rect 1581 2604 2228 2632
rect 1581 2601 1593 2604
rect 1535 2595 1593 2601
rect 2222 2592 2228 2604
rect 2280 2592 2286 2644
rect 9398 2592 9404 2644
rect 9456 2632 9462 2644
rect 9493 2635 9551 2641
rect 9493 2632 9505 2635
rect 9456 2604 9505 2632
rect 9456 2592 9462 2604
rect 9493 2601 9505 2604
rect 9539 2632 9551 2635
rect 9539 2604 9996 2632
rect 9539 2601 9551 2604
rect 9493 2595 9551 2601
rect 5994 2564 6000 2576
rect 5955 2536 6000 2564
rect 5994 2524 6000 2536
rect 6052 2524 6058 2576
rect 9858 2564 9864 2576
rect 9819 2536 9864 2564
rect 9858 2524 9864 2536
rect 9916 2524 9922 2576
rect 9968 2573 9996 2604
rect 10686 2592 10692 2644
rect 10744 2632 10750 2644
rect 10781 2635 10839 2641
rect 10781 2632 10793 2635
rect 10744 2604 10793 2632
rect 10744 2592 10750 2604
rect 10781 2601 10793 2604
rect 10827 2601 10839 2635
rect 10781 2595 10839 2601
rect 21315 2635 21373 2641
rect 21315 2601 21327 2635
rect 21361 2632 21373 2635
rect 21450 2632 21456 2644
rect 21361 2604 21456 2632
rect 21361 2601 21373 2604
rect 21315 2595 21373 2601
rect 21450 2592 21456 2604
rect 21508 2592 21514 2644
rect 9953 2567 10011 2573
rect 9953 2533 9965 2567
rect 9999 2533 10011 2567
rect 9953 2527 10011 2533
rect 10505 2567 10563 2573
rect 10505 2533 10517 2567
rect 10551 2564 10563 2567
rect 10962 2564 10968 2576
rect 10551 2536 10968 2564
rect 10551 2533 10563 2536
rect 10505 2527 10563 2533
rect 10962 2524 10968 2536
rect 11020 2564 11026 2576
rect 11977 2567 12035 2573
rect 11977 2564 11989 2567
rect 11020 2536 11989 2564
rect 11020 2524 11026 2536
rect 11977 2533 11989 2536
rect 12023 2533 12035 2567
rect 12618 2564 12624 2576
rect 12579 2536 12624 2564
rect 11977 2527 12035 2533
rect 12618 2524 12624 2536
rect 12676 2524 12682 2576
rect 1464 2499 1522 2505
rect 1464 2465 1476 2499
rect 1510 2496 1522 2499
rect 1854 2496 1860 2508
rect 1510 2468 1860 2496
rect 1510 2465 1522 2468
rect 1464 2459 1522 2465
rect 1854 2456 1860 2468
rect 1912 2456 1918 2508
rect 4522 2496 4528 2508
rect 4483 2468 4528 2496
rect 4522 2456 4528 2468
rect 4580 2456 4586 2508
rect 5169 2499 5227 2505
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5905 2499 5963 2505
rect 5905 2496 5917 2499
rect 5215 2468 5917 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5905 2465 5917 2468
rect 5951 2496 5963 2499
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 5951 2468 6377 2496
rect 5951 2465 5963 2468
rect 5905 2459 5963 2465
rect 6365 2465 6377 2468
rect 6411 2496 6423 2499
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6411 2468 6929 2496
rect 6411 2465 6423 2468
rect 6365 2459 6423 2465
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 1026 2320 1032 2372
rect 1084 2360 1090 2372
rect 5184 2360 5212 2459
rect 7190 2456 7196 2508
rect 7248 2496 7254 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 7248 2468 7297 2496
rect 7248 2456 7254 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 7653 2499 7711 2505
rect 7653 2465 7665 2499
rect 7699 2465 7711 2499
rect 7653 2459 7711 2465
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 7668 2428 7696 2459
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 8352 2468 8493 2496
rect 8352 2456 8358 2468
rect 8481 2465 8493 2468
rect 8527 2496 8539 2499
rect 9033 2499 9091 2505
rect 9033 2496 9045 2499
rect 8527 2468 9045 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 9033 2465 9045 2468
rect 9079 2465 9091 2499
rect 9033 2459 9091 2465
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2465 11483 2499
rect 11425 2459 11483 2465
rect 7742 2428 7748 2440
rect 6779 2400 7748 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 9858 2388 9864 2440
rect 9916 2428 9922 2440
rect 11149 2431 11207 2437
rect 11149 2428 11161 2431
rect 9916 2400 11161 2428
rect 9916 2388 9922 2400
rect 11149 2397 11161 2400
rect 11195 2397 11207 2431
rect 11440 2428 11468 2459
rect 11606 2456 11612 2508
rect 11664 2496 11670 2508
rect 12437 2499 12495 2505
rect 12437 2496 12449 2499
rect 11664 2468 12449 2496
rect 11664 2456 11670 2468
rect 12437 2465 12449 2468
rect 12483 2496 12495 2499
rect 12713 2499 12771 2505
rect 12713 2496 12725 2499
rect 12483 2468 12725 2496
rect 12483 2465 12495 2468
rect 12437 2459 12495 2465
rect 12713 2465 12725 2468
rect 12759 2465 12771 2499
rect 12713 2459 12771 2465
rect 12802 2456 12808 2508
rect 12860 2496 12866 2508
rect 14236 2499 14294 2505
rect 14236 2496 14248 2499
rect 12860 2468 14248 2496
rect 12860 2456 12866 2468
rect 14236 2465 14248 2468
rect 14282 2496 14294 2499
rect 14645 2499 14703 2505
rect 14645 2496 14657 2499
rect 14282 2468 14657 2496
rect 14282 2465 14294 2468
rect 14236 2459 14294 2465
rect 14645 2465 14657 2468
rect 14691 2465 14703 2499
rect 14645 2459 14703 2465
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2496 15531 2499
rect 15562 2496 15568 2508
rect 15519 2468 15568 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 15562 2456 15568 2468
rect 15620 2496 15626 2508
rect 16025 2499 16083 2505
rect 16025 2496 16037 2499
rect 15620 2468 16037 2496
rect 15620 2456 15626 2468
rect 16025 2465 16037 2468
rect 16071 2465 16083 2499
rect 16574 2496 16580 2508
rect 16535 2468 16580 2496
rect 16025 2459 16083 2465
rect 16574 2456 16580 2468
rect 16632 2496 16638 2508
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 16632 2468 17141 2496
rect 16632 2456 16638 2468
rect 17129 2465 17141 2468
rect 17175 2465 17187 2499
rect 17129 2459 17187 2465
rect 20048 2499 20106 2505
rect 20048 2465 20060 2499
rect 20094 2496 20106 2499
rect 21244 2499 21302 2505
rect 20094 2468 20576 2496
rect 20094 2465 20106 2468
rect 20048 2459 20106 2465
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 11440 2400 13645 2428
rect 11149 2391 11207 2397
rect 13633 2397 13645 2400
rect 13679 2428 13691 2431
rect 14323 2431 14381 2437
rect 14323 2428 14335 2431
rect 13679 2400 14335 2428
rect 13679 2397 13691 2400
rect 13633 2391 13691 2397
rect 14323 2397 14335 2400
rect 14369 2397 14381 2431
rect 14323 2391 14381 2397
rect 1084 2332 5212 2360
rect 8665 2363 8723 2369
rect 1084 2320 1090 2332
rect 8665 2329 8677 2363
rect 8711 2360 8723 2363
rect 9950 2360 9956 2372
rect 8711 2332 9956 2360
rect 8711 2329 8723 2332
rect 8665 2323 8723 2329
rect 9950 2320 9956 2332
rect 10008 2320 10014 2372
rect 11609 2363 11667 2369
rect 11609 2329 11621 2363
rect 11655 2360 11667 2363
rect 13262 2360 13268 2372
rect 11655 2332 13268 2360
rect 11655 2329 11667 2332
rect 11609 2323 11667 2329
rect 13262 2320 13268 2332
rect 13320 2320 13326 2372
rect 15378 2252 15384 2304
rect 15436 2292 15442 2304
rect 15657 2295 15715 2301
rect 15657 2292 15669 2295
rect 15436 2264 15669 2292
rect 15436 2252 15442 2264
rect 15657 2261 15669 2264
rect 15703 2261 15715 2295
rect 15657 2255 15715 2261
rect 16761 2295 16819 2301
rect 16761 2261 16773 2295
rect 16807 2292 16819 2295
rect 16850 2292 16856 2304
rect 16807 2264 16856 2292
rect 16807 2261 16819 2264
rect 16761 2255 16819 2261
rect 16850 2252 16856 2264
rect 16908 2252 16914 2304
rect 17218 2252 17224 2304
rect 17276 2292 17282 2304
rect 20548 2301 20576 2468
rect 21244 2465 21256 2499
rect 21290 2496 21302 2499
rect 21290 2468 21772 2496
rect 21290 2465 21302 2468
rect 21244 2459 21302 2465
rect 20119 2295 20177 2301
rect 20119 2292 20131 2295
rect 17276 2264 20131 2292
rect 17276 2252 17282 2264
rect 20119 2261 20131 2264
rect 20165 2261 20177 2295
rect 20119 2255 20177 2261
rect 20533 2295 20591 2301
rect 20533 2261 20545 2295
rect 20579 2292 20591 2295
rect 21266 2292 21272 2304
rect 20579 2264 21272 2292
rect 20579 2261 20591 2264
rect 20533 2255 20591 2261
rect 21266 2252 21272 2264
rect 21324 2252 21330 2304
rect 21744 2301 21772 2468
rect 21729 2295 21787 2301
rect 21729 2261 21741 2295
rect 21775 2292 21787 2295
rect 22830 2292 22836 2304
rect 21775 2264 22836 2292
rect 21775 2261 21787 2264
rect 21729 2255 21787 2261
rect 22830 2252 22836 2264
rect 22888 2252 22894 2304
rect 1104 2202 22816 2224
rect 1104 2150 4982 2202
rect 5034 2150 5046 2202
rect 5098 2150 5110 2202
rect 5162 2150 5174 2202
rect 5226 2150 12982 2202
rect 13034 2150 13046 2202
rect 13098 2150 13110 2202
rect 13162 2150 13174 2202
rect 13226 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 22816 2202
rect 1104 2128 22816 2150
<< via1 >>
rect 4982 21734 5034 21786
rect 5046 21734 5098 21786
rect 5110 21734 5162 21786
rect 5174 21734 5226 21786
rect 12982 21734 13034 21786
rect 13046 21734 13098 21786
rect 13110 21734 13162 21786
rect 13174 21734 13226 21786
rect 20982 21734 21034 21786
rect 21046 21734 21098 21786
rect 21110 21734 21162 21786
rect 21174 21734 21226 21786
rect 11152 21360 11204 21412
rect 23572 21360 23624 21412
rect 8982 21190 9034 21242
rect 9046 21190 9098 21242
rect 9110 21190 9162 21242
rect 9174 21190 9226 21242
rect 16982 21190 17034 21242
rect 17046 21190 17098 21242
rect 17110 21190 17162 21242
rect 17174 21190 17226 21242
rect 11152 20952 11204 21004
rect 9956 20748 10008 20800
rect 4982 20646 5034 20698
rect 5046 20646 5098 20698
rect 5110 20646 5162 20698
rect 5174 20646 5226 20698
rect 12982 20646 13034 20698
rect 13046 20646 13098 20698
rect 13110 20646 13162 20698
rect 13174 20646 13226 20698
rect 20982 20646 21034 20698
rect 21046 20646 21098 20698
rect 21110 20646 21162 20698
rect 21174 20646 21226 20698
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 3424 20587 3476 20596
rect 3424 20553 3433 20587
rect 3433 20553 3467 20587
rect 3467 20553 3476 20587
rect 3424 20544 3476 20553
rect 10692 20587 10744 20596
rect 10692 20553 10701 20587
rect 10701 20553 10735 20587
rect 10735 20553 10744 20587
rect 10692 20544 10744 20553
rect 11152 20587 11204 20596
rect 11152 20553 11161 20587
rect 11161 20553 11195 20587
rect 11195 20553 11204 20587
rect 11152 20544 11204 20553
rect 12808 20544 12860 20596
rect 5816 20383 5868 20392
rect 5816 20349 5825 20383
rect 5825 20349 5859 20383
rect 5859 20349 5868 20383
rect 5816 20340 5868 20349
rect 12440 20383 12492 20392
rect 2044 20247 2096 20256
rect 2044 20213 2053 20247
rect 2053 20213 2087 20247
rect 2087 20213 2096 20247
rect 2044 20204 2096 20213
rect 3884 20247 3936 20256
rect 3884 20213 3893 20247
rect 3893 20213 3927 20247
rect 3927 20213 3936 20247
rect 3884 20204 3936 20213
rect 5816 20204 5868 20256
rect 12440 20349 12449 20383
rect 12449 20349 12483 20383
rect 12483 20349 12492 20383
rect 12440 20340 12492 20349
rect 17684 20544 17736 20596
rect 21640 20544 21692 20596
rect 22468 20544 22520 20596
rect 10692 20204 10744 20256
rect 16488 20204 16540 20256
rect 20536 20204 20588 20256
rect 21824 20204 21876 20256
rect 8982 20102 9034 20154
rect 9046 20102 9098 20154
rect 9110 20102 9162 20154
rect 9174 20102 9226 20154
rect 16982 20102 17034 20154
rect 17046 20102 17098 20154
rect 17110 20102 17162 20154
rect 17174 20102 17226 20154
rect 3884 20000 3936 20052
rect 12440 20000 12492 20052
rect 1216 19932 1268 19984
rect 11704 19864 11756 19916
rect 2872 19660 2924 19712
rect 8300 19660 8352 19712
rect 4982 19558 5034 19610
rect 5046 19558 5098 19610
rect 5110 19558 5162 19610
rect 5174 19558 5226 19610
rect 12982 19558 13034 19610
rect 13046 19558 13098 19610
rect 13110 19558 13162 19610
rect 13174 19558 13226 19610
rect 20982 19558 21034 19610
rect 21046 19558 21098 19610
rect 21110 19558 21162 19610
rect 21174 19558 21226 19610
rect 1216 19456 1268 19508
rect 11704 19499 11756 19508
rect 11704 19465 11713 19499
rect 11713 19465 11747 19499
rect 11747 19465 11756 19499
rect 11704 19456 11756 19465
rect 15660 19456 15712 19508
rect 10968 19295 11020 19304
rect 10968 19261 10977 19295
rect 10977 19261 11011 19295
rect 11011 19261 11020 19295
rect 10968 19252 11020 19261
rect 8300 19159 8352 19168
rect 8300 19125 8309 19159
rect 8309 19125 8343 19159
rect 8343 19125 8352 19159
rect 8300 19116 8352 19125
rect 11152 19159 11204 19168
rect 11152 19125 11161 19159
rect 11161 19125 11195 19159
rect 11195 19125 11204 19159
rect 11152 19116 11204 19125
rect 14832 19159 14884 19168
rect 14832 19125 14841 19159
rect 14841 19125 14875 19159
rect 14875 19125 14884 19159
rect 14832 19116 14884 19125
rect 8982 19014 9034 19066
rect 9046 19014 9098 19066
rect 9110 19014 9162 19066
rect 9174 19014 9226 19066
rect 16982 19014 17034 19066
rect 17046 19014 17098 19066
rect 17110 19014 17162 19066
rect 17174 19014 17226 19066
rect 8484 18912 8536 18964
rect 11152 18844 11204 18896
rect 1308 18776 1360 18828
rect 6920 18819 6972 18828
rect 6920 18785 6929 18819
rect 6929 18785 6963 18819
rect 6963 18785 6972 18819
rect 6920 18776 6972 18785
rect 13636 18819 13688 18828
rect 13636 18785 13645 18819
rect 13645 18785 13679 18819
rect 13679 18785 13688 18819
rect 13636 18776 13688 18785
rect 20812 18776 20864 18828
rect 21272 18776 21324 18828
rect 10600 18708 10652 18760
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 11704 18683 11756 18692
rect 11704 18649 11713 18683
rect 11713 18649 11747 18683
rect 11747 18649 11756 18683
rect 11704 18640 11756 18649
rect 8116 18572 8168 18624
rect 8392 18615 8444 18624
rect 8392 18581 8401 18615
rect 8401 18581 8435 18615
rect 8435 18581 8444 18615
rect 8392 18572 8444 18581
rect 10968 18572 11020 18624
rect 16028 18572 16080 18624
rect 4982 18470 5034 18522
rect 5046 18470 5098 18522
rect 5110 18470 5162 18522
rect 5174 18470 5226 18522
rect 12982 18470 13034 18522
rect 13046 18470 13098 18522
rect 13110 18470 13162 18522
rect 13174 18470 13226 18522
rect 20982 18470 21034 18522
rect 21046 18470 21098 18522
rect 21110 18470 21162 18522
rect 21174 18470 21226 18522
rect 1308 18368 1360 18420
rect 6184 18411 6236 18420
rect 6184 18377 6193 18411
rect 6193 18377 6227 18411
rect 6227 18377 6236 18411
rect 6184 18368 6236 18377
rect 10600 18411 10652 18420
rect 10600 18377 10609 18411
rect 10609 18377 10643 18411
rect 10643 18377 10652 18411
rect 10600 18368 10652 18377
rect 11152 18368 11204 18420
rect 13360 18411 13412 18420
rect 13360 18377 13369 18411
rect 13369 18377 13403 18411
rect 13403 18377 13412 18411
rect 13360 18368 13412 18377
rect 14832 18368 14884 18420
rect 20812 18368 20864 18420
rect 6920 18300 6972 18352
rect 5908 18232 5960 18284
rect 8668 18275 8720 18284
rect 1216 18164 1268 18216
rect 6184 18164 6236 18216
rect 8668 18241 8677 18275
rect 8677 18241 8711 18275
rect 8711 18241 8720 18275
rect 8668 18232 8720 18241
rect 11704 18232 11756 18284
rect 13636 18232 13688 18284
rect 8392 18139 8444 18148
rect 8392 18105 8401 18139
rect 8401 18105 8435 18139
rect 8435 18105 8444 18139
rect 8392 18096 8444 18105
rect 10876 18139 10928 18148
rect 2504 18028 2556 18080
rect 7932 18028 7984 18080
rect 8208 18071 8260 18080
rect 8208 18037 8217 18071
rect 8217 18037 8251 18071
rect 8251 18037 8260 18071
rect 10876 18105 10885 18139
rect 10885 18105 10919 18139
rect 10919 18105 10928 18139
rect 10876 18096 10928 18105
rect 10968 18139 11020 18148
rect 10968 18105 10977 18139
rect 10977 18105 11011 18139
rect 11011 18105 11020 18139
rect 10968 18096 11020 18105
rect 14280 18139 14332 18148
rect 8208 18028 8260 18037
rect 13360 18028 13412 18080
rect 14280 18105 14289 18139
rect 14289 18105 14323 18139
rect 14323 18105 14332 18139
rect 14280 18096 14332 18105
rect 8982 17926 9034 17978
rect 9046 17926 9098 17978
rect 9110 17926 9162 17978
rect 9174 17926 9226 17978
rect 16982 17926 17034 17978
rect 17046 17926 17098 17978
rect 17110 17926 17162 17978
rect 17174 17926 17226 17978
rect 2872 17824 2924 17876
rect 8852 17824 8904 17876
rect 6000 17756 6052 17808
rect 8024 17799 8076 17808
rect 8024 17765 8033 17799
rect 8033 17765 8067 17799
rect 8067 17765 8076 17799
rect 8024 17756 8076 17765
rect 10232 17799 10284 17808
rect 10232 17765 10241 17799
rect 10241 17765 10275 17799
rect 10275 17765 10284 17799
rect 10232 17756 10284 17765
rect 10876 17756 10928 17808
rect 13636 17799 13688 17808
rect 13636 17765 13645 17799
rect 13645 17765 13679 17799
rect 13679 17765 13688 17799
rect 13636 17756 13688 17765
rect 14280 17756 14332 17808
rect 112 17688 164 17740
rect 1860 17688 1912 17740
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 11704 17731 11756 17740
rect 11704 17697 11713 17731
rect 11713 17697 11747 17731
rect 11747 17697 11756 17731
rect 11704 17688 11756 17697
rect 15384 17731 15436 17740
rect 15384 17697 15402 17731
rect 15402 17697 15436 17731
rect 15384 17688 15436 17697
rect 20076 17688 20128 17740
rect 21272 17688 21324 17740
rect 5632 17663 5684 17672
rect 5632 17629 5641 17663
rect 5641 17629 5675 17663
rect 5675 17629 5684 17663
rect 5632 17620 5684 17629
rect 5908 17663 5960 17672
rect 5908 17629 5917 17663
rect 5917 17629 5951 17663
rect 5951 17629 5960 17663
rect 5908 17620 5960 17629
rect 7932 17663 7984 17672
rect 7932 17629 7941 17663
rect 7941 17629 7975 17663
rect 7975 17629 7984 17663
rect 7932 17620 7984 17629
rect 8668 17620 8720 17672
rect 10140 17663 10192 17672
rect 10140 17629 10149 17663
rect 10149 17629 10183 17663
rect 10183 17629 10192 17663
rect 10140 17620 10192 17629
rect 10784 17620 10836 17672
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13544 17620 13596 17629
rect 13268 17595 13320 17604
rect 13268 17561 13277 17595
rect 13277 17561 13311 17595
rect 13311 17561 13320 17595
rect 13268 17552 13320 17561
rect 1676 17484 1728 17536
rect 2688 17527 2740 17536
rect 2688 17493 2697 17527
rect 2697 17493 2731 17527
rect 2731 17493 2740 17527
rect 2688 17484 2740 17493
rect 5356 17484 5408 17536
rect 19340 17484 19392 17536
rect 4982 17382 5034 17434
rect 5046 17382 5098 17434
rect 5110 17382 5162 17434
rect 5174 17382 5226 17434
rect 12982 17382 13034 17434
rect 13046 17382 13098 17434
rect 13110 17382 13162 17434
rect 13174 17382 13226 17434
rect 20982 17382 21034 17434
rect 21046 17382 21098 17434
rect 21110 17382 21162 17434
rect 21174 17382 21226 17434
rect 1860 17323 1912 17332
rect 1860 17289 1869 17323
rect 1869 17289 1903 17323
rect 1903 17289 1912 17323
rect 1860 17280 1912 17289
rect 8208 17323 8260 17332
rect 8208 17289 8217 17323
rect 8217 17289 8251 17323
rect 8251 17289 8260 17323
rect 8208 17280 8260 17289
rect 10232 17280 10284 17332
rect 10508 17280 10560 17332
rect 11704 17323 11756 17332
rect 11704 17289 11713 17323
rect 11713 17289 11747 17323
rect 11747 17289 11756 17323
rect 11704 17280 11756 17289
rect 15384 17323 15436 17332
rect 15384 17289 15393 17323
rect 15393 17289 15427 17323
rect 15427 17289 15436 17323
rect 15384 17280 15436 17289
rect 21272 17280 21324 17332
rect 7932 17212 7984 17264
rect 2504 17144 2556 17196
rect 3148 17187 3200 17196
rect 3148 17153 3157 17187
rect 3157 17153 3191 17187
rect 3191 17153 3200 17187
rect 3148 17144 3200 17153
rect 5908 17187 5960 17196
rect 5908 17153 5917 17187
rect 5917 17153 5951 17187
rect 5951 17153 5960 17187
rect 5908 17144 5960 17153
rect 8116 17144 8168 17196
rect 10140 17144 10192 17196
rect 10876 17187 10928 17196
rect 10876 17153 10885 17187
rect 10885 17153 10919 17187
rect 10919 17153 10928 17187
rect 10876 17144 10928 17153
rect 13268 17187 13320 17196
rect 13268 17153 13277 17187
rect 13277 17153 13311 17187
rect 13311 17153 13320 17187
rect 13268 17144 13320 17153
rect 13544 17187 13596 17196
rect 13544 17153 13553 17187
rect 13553 17153 13587 17187
rect 13587 17153 13596 17187
rect 13544 17144 13596 17153
rect 1467 17119 1519 17128
rect 1467 17085 1476 17119
rect 1476 17085 1510 17119
rect 1510 17085 1519 17119
rect 1467 17076 1519 17085
rect 8024 17076 8076 17128
rect 8392 17119 8444 17128
rect 8392 17085 8401 17119
rect 8401 17085 8435 17119
rect 8435 17085 8444 17119
rect 8392 17076 8444 17085
rect 2780 17051 2832 17060
rect 2780 17017 2789 17051
rect 2789 17017 2823 17051
rect 2823 17017 2832 17051
rect 2780 17008 2832 17017
rect 3792 17008 3844 17060
rect 5356 17051 5408 17060
rect 5356 17017 5365 17051
rect 5365 17017 5399 17051
rect 5399 17017 5408 17051
rect 5356 17008 5408 17017
rect 5632 17008 5684 17060
rect 10324 17008 10376 17060
rect 1860 16940 1912 16992
rect 6000 16940 6052 16992
rect 10784 17008 10836 17060
rect 12808 16940 12860 16992
rect 13452 16940 13504 16992
rect 13636 16940 13688 16992
rect 8982 16838 9034 16890
rect 9046 16838 9098 16890
rect 9110 16838 9162 16890
rect 9174 16838 9226 16890
rect 16982 16838 17034 16890
rect 17046 16838 17098 16890
rect 17110 16838 17162 16890
rect 17174 16838 17226 16890
rect 2504 16736 2556 16788
rect 8392 16779 8444 16788
rect 8392 16745 8401 16779
rect 8401 16745 8435 16779
rect 8435 16745 8444 16779
rect 8392 16736 8444 16745
rect 2688 16668 2740 16720
rect 3148 16711 3200 16720
rect 3148 16677 3157 16711
rect 3157 16677 3191 16711
rect 3191 16677 3200 16711
rect 3148 16668 3200 16677
rect 6000 16711 6052 16720
rect 6000 16677 6009 16711
rect 6009 16677 6043 16711
rect 6043 16677 6052 16711
rect 6000 16668 6052 16677
rect 8024 16668 8076 16720
rect 1952 16600 2004 16652
rect 5356 16643 5408 16652
rect 5356 16609 5365 16643
rect 5365 16609 5399 16643
rect 5399 16609 5408 16643
rect 5356 16600 5408 16609
rect 10416 16668 10468 16720
rect 11888 16668 11940 16720
rect 13544 16736 13596 16788
rect 10140 16643 10192 16652
rect 10140 16609 10149 16643
rect 10149 16609 10183 16643
rect 10183 16609 10192 16643
rect 10140 16600 10192 16609
rect 21272 16600 21324 16652
rect 2228 16532 2280 16584
rect 8392 16532 8444 16584
rect 10232 16575 10284 16584
rect 10232 16541 10241 16575
rect 10241 16541 10275 16575
rect 10275 16541 10284 16575
rect 10232 16532 10284 16541
rect 12716 16575 12768 16584
rect 12716 16541 12725 16575
rect 12725 16541 12759 16575
rect 12759 16541 12768 16575
rect 12716 16532 12768 16541
rect 1768 16396 1820 16448
rect 7104 16439 7156 16448
rect 7104 16405 7113 16439
rect 7113 16405 7147 16439
rect 7147 16405 7156 16439
rect 7104 16396 7156 16405
rect 10324 16396 10376 16448
rect 20444 16396 20496 16448
rect 4982 16294 5034 16346
rect 5046 16294 5098 16346
rect 5110 16294 5162 16346
rect 5174 16294 5226 16346
rect 12982 16294 13034 16346
rect 13046 16294 13098 16346
rect 13110 16294 13162 16346
rect 13174 16294 13226 16346
rect 20982 16294 21034 16346
rect 21046 16294 21098 16346
rect 21110 16294 21162 16346
rect 21174 16294 21226 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 2688 16192 2740 16244
rect 3792 16235 3844 16244
rect 3792 16201 3801 16235
rect 3801 16201 3835 16235
rect 3835 16201 3844 16235
rect 3792 16192 3844 16201
rect 5356 16192 5408 16244
rect 10508 16235 10560 16244
rect 10508 16201 10517 16235
rect 10517 16201 10551 16235
rect 10551 16201 10560 16235
rect 10508 16192 10560 16201
rect 11888 16235 11940 16244
rect 11888 16201 11897 16235
rect 11897 16201 11931 16235
rect 11931 16201 11940 16235
rect 11888 16192 11940 16201
rect 12808 16192 12860 16244
rect 21272 16192 21324 16244
rect 7380 16099 7432 16108
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 13452 16167 13504 16176
rect 13452 16133 13461 16167
rect 13461 16133 13495 16167
rect 13495 16133 13504 16167
rect 13452 16124 13504 16133
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 2872 16031 2924 16040
rect 2872 15997 2881 16031
rect 2881 15997 2915 16031
rect 2915 15997 2924 16031
rect 2872 15988 2924 15997
rect 4712 16031 4764 16040
rect 4712 15997 4721 16031
rect 4721 15997 4755 16031
rect 4755 15997 4764 16031
rect 4712 15988 4764 15997
rect 9772 15988 9824 16040
rect 13268 15988 13320 16040
rect 2780 15963 2832 15972
rect 2780 15929 2789 15963
rect 2789 15929 2823 15963
rect 2823 15929 2832 15963
rect 2780 15920 2832 15929
rect 7104 15963 7156 15972
rect 7104 15929 7113 15963
rect 7113 15929 7147 15963
rect 7147 15929 7156 15963
rect 7104 15920 7156 15929
rect 1952 15895 2004 15904
rect 1952 15861 1961 15895
rect 1961 15861 1995 15895
rect 1995 15861 2004 15895
rect 1952 15852 2004 15861
rect 2228 15852 2280 15904
rect 6552 15895 6604 15904
rect 6552 15861 6561 15895
rect 6561 15861 6595 15895
rect 6595 15861 6604 15895
rect 10048 15920 10100 15972
rect 8024 15895 8076 15904
rect 6552 15852 6604 15861
rect 8024 15861 8033 15895
rect 8033 15861 8067 15895
rect 8067 15861 8076 15895
rect 8024 15852 8076 15861
rect 8392 15895 8444 15904
rect 8392 15861 8401 15895
rect 8401 15861 8435 15895
rect 8435 15861 8444 15895
rect 8392 15852 8444 15861
rect 10416 15852 10468 15904
rect 12256 15895 12308 15904
rect 12256 15861 12265 15895
rect 12265 15861 12299 15895
rect 12299 15861 12308 15895
rect 12256 15852 12308 15861
rect 8982 15750 9034 15802
rect 9046 15750 9098 15802
rect 9110 15750 9162 15802
rect 9174 15750 9226 15802
rect 16982 15750 17034 15802
rect 17046 15750 17098 15802
rect 17110 15750 17162 15802
rect 17174 15750 17226 15802
rect 1400 15648 1452 15700
rect 2872 15648 2924 15700
rect 7104 15648 7156 15700
rect 10140 15648 10192 15700
rect 10968 15691 11020 15700
rect 10968 15657 10977 15691
rect 10977 15657 11011 15691
rect 11011 15657 11020 15691
rect 10968 15648 11020 15657
rect 12808 15648 12860 15700
rect 6552 15580 6604 15632
rect 7196 15623 7248 15632
rect 7196 15589 7205 15623
rect 7205 15589 7239 15623
rect 7239 15589 7248 15623
rect 7196 15580 7248 15589
rect 2688 15555 2740 15564
rect 2688 15521 2697 15555
rect 2697 15521 2731 15555
rect 2731 15521 2740 15555
rect 2688 15512 2740 15521
rect 2964 15555 3016 15564
rect 2964 15521 2973 15555
rect 2973 15521 3007 15555
rect 3007 15521 3016 15555
rect 2964 15512 3016 15521
rect 6092 15555 6144 15564
rect 6092 15521 6101 15555
rect 6101 15521 6135 15555
rect 6135 15521 6144 15555
rect 6092 15512 6144 15521
rect 10232 15512 10284 15564
rect 1584 15444 1636 15496
rect 7104 15487 7156 15496
rect 7104 15453 7113 15487
rect 7113 15453 7147 15487
rect 7147 15453 7156 15487
rect 7104 15444 7156 15453
rect 7380 15487 7432 15496
rect 7380 15453 7389 15487
rect 7389 15453 7423 15487
rect 7423 15453 7432 15487
rect 7380 15444 7432 15453
rect 10048 15376 10100 15428
rect 12256 15580 12308 15632
rect 12164 15487 12216 15496
rect 12164 15453 12173 15487
rect 12173 15453 12207 15487
rect 12207 15453 12216 15487
rect 12164 15444 12216 15453
rect 4712 15351 4764 15360
rect 4712 15317 4721 15351
rect 4721 15317 4755 15351
rect 4755 15317 4764 15351
rect 4712 15308 4764 15317
rect 6828 15351 6880 15360
rect 6828 15317 6837 15351
rect 6837 15317 6871 15351
rect 6871 15317 6880 15351
rect 6828 15308 6880 15317
rect 11152 15308 11204 15360
rect 12716 15308 12768 15360
rect 4982 15206 5034 15258
rect 5046 15206 5098 15258
rect 5110 15206 5162 15258
rect 5174 15206 5226 15258
rect 12982 15206 13034 15258
rect 13046 15206 13098 15258
rect 13110 15206 13162 15258
rect 13174 15206 13226 15258
rect 20982 15206 21034 15258
rect 21046 15206 21098 15258
rect 21110 15206 21162 15258
rect 21174 15206 21226 15258
rect 2964 15104 3016 15156
rect 2136 14900 2188 14952
rect 6092 15104 6144 15156
rect 7196 15104 7248 15156
rect 8944 15104 8996 15156
rect 10232 15036 10284 15088
rect 14556 15079 14608 15088
rect 14556 15045 14565 15079
rect 14565 15045 14599 15079
rect 14599 15045 14608 15079
rect 14556 15036 14608 15045
rect 4712 15011 4764 15020
rect 4712 14977 4721 15011
rect 4721 14977 4755 15011
rect 4755 14977 4764 15011
rect 4712 14968 4764 14977
rect 9772 15011 9824 15020
rect 9772 14977 9781 15011
rect 9781 14977 9815 15011
rect 9815 14977 9824 15011
rect 9772 14968 9824 14977
rect 10048 14968 10100 15020
rect 12256 15011 12308 15020
rect 12256 14977 12265 15011
rect 12265 14977 12299 15011
rect 12299 14977 12308 15011
rect 12256 14968 12308 14977
rect 13268 14968 13320 15020
rect 4436 14943 4488 14952
rect 4436 14909 4445 14943
rect 4445 14909 4479 14943
rect 4479 14909 4488 14943
rect 4436 14900 4488 14909
rect 4620 14943 4672 14952
rect 4620 14909 4629 14943
rect 4629 14909 4663 14943
rect 4663 14909 4672 14943
rect 4620 14900 4672 14909
rect 5632 14900 5684 14952
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 2044 14807 2096 14816
rect 2044 14773 2053 14807
rect 2053 14773 2087 14807
rect 2087 14773 2096 14807
rect 2044 14764 2096 14773
rect 2688 14764 2740 14816
rect 6276 14764 6328 14816
rect 8024 14832 8076 14884
rect 9312 14900 9364 14952
rect 10140 14900 10192 14952
rect 12164 14900 12216 14952
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12440 14900 12492 14909
rect 11980 14832 12032 14884
rect 14372 14943 14424 14952
rect 14372 14909 14381 14943
rect 14381 14909 14415 14943
rect 14415 14909 14424 14943
rect 14372 14900 14424 14909
rect 15660 14900 15712 14952
rect 9404 14764 9456 14816
rect 8982 14662 9034 14714
rect 9046 14662 9098 14714
rect 9110 14662 9162 14714
rect 9174 14662 9226 14714
rect 16982 14662 17034 14714
rect 17046 14662 17098 14714
rect 17110 14662 17162 14714
rect 17174 14662 17226 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 8760 14560 8812 14612
rect 9312 14603 9364 14612
rect 9312 14569 9321 14603
rect 9321 14569 9355 14603
rect 9355 14569 9364 14603
rect 9312 14560 9364 14569
rect 10508 14560 10560 14612
rect 12440 14603 12492 14612
rect 12440 14569 12449 14603
rect 12449 14569 12483 14603
rect 12483 14569 12492 14603
rect 12440 14560 12492 14569
rect 14372 14560 14424 14612
rect 1860 14535 1912 14544
rect 1860 14501 1869 14535
rect 1869 14501 1903 14535
rect 1903 14501 1912 14535
rect 1860 14492 1912 14501
rect 2044 14492 2096 14544
rect 5632 14535 5684 14544
rect 5632 14501 5641 14535
rect 5641 14501 5675 14535
rect 5675 14501 5684 14535
rect 5632 14492 5684 14501
rect 5816 14492 5868 14544
rect 6828 14492 6880 14544
rect 9404 14492 9456 14544
rect 12164 14535 12216 14544
rect 4436 14424 4488 14476
rect 2596 14356 2648 14408
rect 5724 14424 5776 14476
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 12164 14501 12173 14535
rect 12173 14501 12207 14535
rect 12207 14501 12216 14535
rect 12164 14492 12216 14501
rect 15476 14535 15528 14544
rect 15476 14501 15485 14535
rect 15485 14501 15519 14535
rect 15519 14501 15528 14535
rect 15476 14492 15528 14501
rect 11796 14424 11848 14476
rect 11980 14467 12032 14476
rect 11980 14433 11989 14467
rect 11989 14433 12023 14467
rect 12023 14433 12032 14467
rect 11980 14424 12032 14433
rect 13452 14424 13504 14476
rect 5356 14356 5408 14408
rect 10508 14356 10560 14408
rect 14740 14356 14792 14408
rect 15660 14399 15712 14408
rect 15660 14365 15669 14399
rect 15669 14365 15703 14399
rect 15703 14365 15712 14399
rect 15660 14356 15712 14365
rect 7104 14331 7156 14340
rect 7104 14297 7113 14331
rect 7113 14297 7147 14331
rect 7147 14297 7156 14331
rect 7104 14288 7156 14297
rect 3792 14263 3844 14272
rect 3792 14229 3801 14263
rect 3801 14229 3835 14263
rect 3835 14229 3844 14263
rect 3792 14220 3844 14229
rect 8024 14220 8076 14272
rect 9772 14220 9824 14272
rect 14924 14263 14976 14272
rect 14924 14229 14933 14263
rect 14933 14229 14967 14263
rect 14967 14229 14976 14263
rect 14924 14220 14976 14229
rect 4982 14118 5034 14170
rect 5046 14118 5098 14170
rect 5110 14118 5162 14170
rect 5174 14118 5226 14170
rect 12982 14118 13034 14170
rect 13046 14118 13098 14170
rect 13110 14118 13162 14170
rect 13174 14118 13226 14170
rect 20982 14118 21034 14170
rect 21046 14118 21098 14170
rect 21110 14118 21162 14170
rect 21174 14118 21226 14170
rect 2044 14016 2096 14068
rect 2136 14016 2188 14068
rect 1860 13948 1912 14000
rect 5356 14016 5408 14068
rect 5816 14059 5868 14068
rect 5816 14025 5825 14059
rect 5825 14025 5859 14059
rect 5859 14025 5868 14059
rect 5816 14016 5868 14025
rect 10048 14059 10100 14068
rect 10048 14025 10057 14059
rect 10057 14025 10091 14059
rect 10091 14025 10100 14059
rect 10048 14016 10100 14025
rect 11796 14059 11848 14068
rect 11796 14025 11805 14059
rect 11805 14025 11839 14059
rect 11839 14025 11848 14059
rect 11796 14016 11848 14025
rect 14740 14059 14792 14068
rect 14740 14025 14749 14059
rect 14749 14025 14783 14059
rect 14783 14025 14792 14059
rect 14740 14016 14792 14025
rect 15476 14016 15528 14068
rect 1768 13880 1820 13932
rect 3792 13923 3844 13932
rect 3792 13889 3801 13923
rect 3801 13889 3835 13923
rect 3835 13889 3844 13923
rect 3792 13880 3844 13889
rect 8852 13880 8904 13932
rect 14924 13923 14976 13932
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 14924 13880 14976 13889
rect 15660 13880 15712 13932
rect 16488 13923 16540 13932
rect 16488 13889 16497 13923
rect 16497 13889 16531 13923
rect 16531 13889 16540 13923
rect 16488 13880 16540 13889
rect 17316 13880 17368 13932
rect 6828 13812 6880 13864
rect 2136 13744 2188 13796
rect 2596 13787 2648 13796
rect 2596 13753 2605 13787
rect 2605 13753 2639 13787
rect 2639 13753 2648 13787
rect 2596 13744 2648 13753
rect 3148 13744 3200 13796
rect 7564 13787 7616 13796
rect 2780 13676 2832 13728
rect 7564 13753 7573 13787
rect 7573 13753 7607 13787
rect 7607 13753 7616 13787
rect 7564 13744 7616 13753
rect 9312 13744 9364 13796
rect 9864 13744 9916 13796
rect 12532 13787 12584 13796
rect 12532 13753 12541 13787
rect 12541 13753 12575 13787
rect 12575 13753 12584 13787
rect 12532 13744 12584 13753
rect 15016 13787 15068 13796
rect 4436 13676 4488 13728
rect 5724 13676 5776 13728
rect 11612 13676 11664 13728
rect 11704 13676 11756 13728
rect 12164 13719 12216 13728
rect 12164 13685 12173 13719
rect 12173 13685 12207 13719
rect 12207 13685 12216 13719
rect 12164 13676 12216 13685
rect 12440 13676 12492 13728
rect 15016 13753 15025 13787
rect 15025 13753 15059 13787
rect 15059 13753 15068 13787
rect 15016 13744 15068 13753
rect 16580 13787 16632 13796
rect 16580 13753 16589 13787
rect 16589 13753 16623 13787
rect 16623 13753 16632 13787
rect 16580 13744 16632 13753
rect 13452 13719 13504 13728
rect 13452 13685 13461 13719
rect 13461 13685 13495 13719
rect 13495 13685 13504 13719
rect 13452 13676 13504 13685
rect 8982 13574 9034 13626
rect 9046 13574 9098 13626
rect 9110 13574 9162 13626
rect 9174 13574 9226 13626
rect 16982 13574 17034 13626
rect 17046 13574 17098 13626
rect 17110 13574 17162 13626
rect 17174 13574 17226 13626
rect 1768 13472 1820 13524
rect 3792 13472 3844 13524
rect 6276 13515 6328 13524
rect 6276 13481 6285 13515
rect 6285 13481 6319 13515
rect 6319 13481 6328 13515
rect 6276 13472 6328 13481
rect 6828 13515 6880 13524
rect 6828 13481 6837 13515
rect 6837 13481 6871 13515
rect 6871 13481 6880 13515
rect 6828 13472 6880 13481
rect 8852 13472 8904 13524
rect 11520 13472 11572 13524
rect 12532 13472 12584 13524
rect 15476 13472 15528 13524
rect 16488 13515 16540 13524
rect 16488 13481 16497 13515
rect 16497 13481 16531 13515
rect 16531 13481 16540 13515
rect 16488 13472 16540 13481
rect 7564 13404 7616 13456
rect 9772 13404 9824 13456
rect 10232 13404 10284 13456
rect 13268 13404 13320 13456
rect 17040 13447 17092 13456
rect 17040 13413 17049 13447
rect 17049 13413 17083 13447
rect 17083 13413 17092 13447
rect 17040 13404 17092 13413
rect 1768 13379 1820 13388
rect 1768 13345 1777 13379
rect 1777 13345 1811 13379
rect 1811 13345 1820 13379
rect 1768 13336 1820 13345
rect 4068 13379 4120 13388
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 4252 13336 4304 13388
rect 15016 13336 15068 13388
rect 15476 13379 15528 13388
rect 15476 13345 15485 13379
rect 15485 13345 15519 13379
rect 15519 13345 15528 13379
rect 15476 13336 15528 13345
rect 21456 13336 21508 13388
rect 5908 13311 5960 13320
rect 5908 13277 5917 13311
rect 5917 13277 5951 13311
rect 5951 13277 5960 13311
rect 5908 13268 5960 13277
rect 8024 13311 8076 13320
rect 8024 13277 8033 13311
rect 8033 13277 8067 13311
rect 8067 13277 8076 13311
rect 8024 13268 8076 13277
rect 9772 13311 9824 13320
rect 9772 13277 9781 13311
rect 9781 13277 9815 13311
rect 9815 13277 9824 13311
rect 9772 13268 9824 13277
rect 9864 13268 9916 13320
rect 11336 13268 11388 13320
rect 11612 13268 11664 13320
rect 12808 13268 12860 13320
rect 13452 13311 13504 13320
rect 13452 13277 13461 13311
rect 13461 13277 13495 13311
rect 13495 13277 13504 13311
rect 13452 13268 13504 13277
rect 17316 13311 17368 13320
rect 8116 13200 8168 13252
rect 16856 13200 16908 13252
rect 17316 13277 17325 13311
rect 17325 13277 17359 13311
rect 17359 13277 17368 13311
rect 17316 13268 17368 13277
rect 1860 13175 1912 13184
rect 1860 13141 1869 13175
rect 1869 13141 1903 13175
rect 1903 13141 1912 13175
rect 1860 13132 1912 13141
rect 2964 13175 3016 13184
rect 2964 13141 2973 13175
rect 2973 13141 3007 13175
rect 3007 13141 3016 13175
rect 2964 13132 3016 13141
rect 3700 13175 3752 13184
rect 3700 13141 3709 13175
rect 3709 13141 3743 13175
rect 3743 13141 3752 13175
rect 3700 13132 3752 13141
rect 5724 13132 5776 13184
rect 6736 13132 6788 13184
rect 10140 13132 10192 13184
rect 11244 13132 11296 13184
rect 12440 13175 12492 13184
rect 12440 13141 12449 13175
rect 12449 13141 12483 13175
rect 12483 13141 12492 13175
rect 12440 13132 12492 13141
rect 14280 13175 14332 13184
rect 14280 13141 14289 13175
rect 14289 13141 14323 13175
rect 14323 13141 14332 13175
rect 14280 13132 14332 13141
rect 20812 13132 20864 13184
rect 4982 13030 5034 13082
rect 5046 13030 5098 13082
rect 5110 13030 5162 13082
rect 5174 13030 5226 13082
rect 12982 13030 13034 13082
rect 13046 13030 13098 13082
rect 13110 13030 13162 13082
rect 13174 13030 13226 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 2688 12928 2740 12980
rect 1768 12860 1820 12912
rect 3056 12903 3108 12912
rect 3056 12869 3065 12903
rect 3065 12869 3099 12903
rect 3099 12869 3108 12903
rect 3056 12860 3108 12869
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 2964 12792 3016 12844
rect 4068 12928 4120 12980
rect 7564 12928 7616 12980
rect 9312 12928 9364 12980
rect 10048 12928 10100 12980
rect 10232 12971 10284 12980
rect 10232 12937 10241 12971
rect 10241 12937 10275 12971
rect 10275 12937 10284 12971
rect 10232 12928 10284 12937
rect 15476 12971 15528 12980
rect 15476 12937 15485 12971
rect 15485 12937 15519 12971
rect 15519 12937 15528 12971
rect 15476 12928 15528 12937
rect 16580 12928 16632 12980
rect 21456 12971 21508 12980
rect 21456 12937 21465 12971
rect 21465 12937 21499 12971
rect 21499 12937 21508 12971
rect 21456 12928 21508 12937
rect 4436 12860 4488 12912
rect 6276 12860 6328 12912
rect 6368 12860 6420 12912
rect 11428 12860 11480 12912
rect 5908 12835 5960 12844
rect 5908 12801 5917 12835
rect 5917 12801 5951 12835
rect 5951 12801 5960 12835
rect 5908 12792 5960 12801
rect 9312 12792 9364 12844
rect 11336 12835 11388 12844
rect 11336 12801 11345 12835
rect 11345 12801 11379 12835
rect 11379 12801 11388 12835
rect 11336 12792 11388 12801
rect 13268 12792 13320 12844
rect 14280 12835 14332 12844
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 20444 12835 20496 12844
rect 20444 12801 20453 12835
rect 20453 12801 20487 12835
rect 20487 12801 20496 12835
rect 20444 12792 20496 12801
rect 3700 12724 3752 12776
rect 4528 12724 4580 12776
rect 5080 12724 5132 12776
rect 5448 12767 5500 12776
rect 5448 12733 5457 12767
rect 5457 12733 5491 12767
rect 5491 12733 5500 12767
rect 5448 12724 5500 12733
rect 5724 12767 5776 12776
rect 5724 12733 5733 12767
rect 5733 12733 5767 12767
rect 5767 12733 5776 12767
rect 5724 12724 5776 12733
rect 6552 12724 6604 12776
rect 6736 12724 6788 12776
rect 10508 12724 10560 12776
rect 11244 12767 11296 12776
rect 11244 12733 11253 12767
rect 11253 12733 11287 12767
rect 11287 12733 11296 12767
rect 11244 12724 11296 12733
rect 12440 12724 12492 12776
rect 16580 12724 16632 12776
rect 17040 12767 17092 12776
rect 17040 12733 17049 12767
rect 17049 12733 17083 12767
rect 17083 12733 17092 12767
rect 17040 12724 17092 12733
rect 1860 12656 1912 12708
rect 2044 12656 2096 12708
rect 6276 12656 6328 12708
rect 11520 12656 11572 12708
rect 13452 12656 13504 12708
rect 16212 12656 16264 12708
rect 21088 12699 21140 12708
rect 4068 12588 4120 12640
rect 5448 12588 5500 12640
rect 6460 12588 6512 12640
rect 6644 12588 6696 12640
rect 8116 12631 8168 12640
rect 8116 12597 8125 12631
rect 8125 12597 8159 12631
rect 8159 12597 8168 12631
rect 8116 12588 8168 12597
rect 10508 12588 10560 12640
rect 20168 12631 20220 12640
rect 20168 12597 20177 12631
rect 20177 12597 20211 12631
rect 20211 12597 20220 12631
rect 21088 12665 21097 12699
rect 21097 12665 21131 12699
rect 21131 12665 21140 12699
rect 21088 12656 21140 12665
rect 20168 12588 20220 12597
rect 8982 12486 9034 12538
rect 9046 12486 9098 12538
rect 9110 12486 9162 12538
rect 9174 12486 9226 12538
rect 16982 12486 17034 12538
rect 17046 12486 17098 12538
rect 17110 12486 17162 12538
rect 17174 12486 17226 12538
rect 3056 12384 3108 12436
rect 5080 12384 5132 12436
rect 9312 12384 9364 12436
rect 11336 12384 11388 12436
rect 12808 12384 12860 12436
rect 16580 12427 16632 12436
rect 16580 12393 16589 12427
rect 16589 12393 16623 12427
rect 16623 12393 16632 12427
rect 16580 12384 16632 12393
rect 20444 12427 20496 12436
rect 20444 12393 20453 12427
rect 20453 12393 20487 12427
rect 20487 12393 20496 12427
rect 20444 12384 20496 12393
rect 1768 12359 1820 12368
rect 1768 12325 1777 12359
rect 1777 12325 1811 12359
rect 1811 12325 1820 12359
rect 1768 12316 1820 12325
rect 4252 12316 4304 12368
rect 4436 12359 4488 12368
rect 4436 12325 4439 12359
rect 4439 12325 4473 12359
rect 4473 12325 4488 12359
rect 4436 12316 4488 12325
rect 11520 12316 11572 12368
rect 14280 12316 14332 12368
rect 16212 12316 16264 12368
rect 20168 12316 20220 12368
rect 4068 12291 4120 12300
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 4068 12248 4120 12257
rect 5540 12248 5592 12300
rect 7380 12291 7432 12300
rect 1676 12223 1728 12232
rect 1676 12189 1685 12223
rect 1685 12189 1719 12223
rect 1719 12189 1728 12223
rect 1676 12180 1728 12189
rect 2044 12223 2096 12232
rect 2044 12189 2053 12223
rect 2053 12189 2087 12223
rect 2087 12189 2096 12223
rect 2044 12180 2096 12189
rect 5632 12180 5684 12232
rect 6276 12180 6328 12232
rect 6368 12112 6420 12164
rect 7380 12257 7389 12291
rect 7389 12257 7423 12291
rect 7423 12257 7432 12291
rect 7380 12248 7432 12257
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 10048 12248 10100 12300
rect 11428 12291 11480 12300
rect 11428 12257 11434 12291
rect 11434 12257 11480 12291
rect 11428 12248 11480 12257
rect 12716 12248 12768 12300
rect 13360 12248 13412 12300
rect 14188 12291 14240 12300
rect 14188 12257 14197 12291
rect 14197 12257 14231 12291
rect 14231 12257 14240 12291
rect 14188 12248 14240 12257
rect 19616 12248 19668 12300
rect 20812 12316 20864 12368
rect 21732 12316 21784 12368
rect 10968 12180 11020 12232
rect 15660 12223 15712 12232
rect 15660 12189 15669 12223
rect 15669 12189 15703 12223
rect 15703 12189 15712 12223
rect 15660 12180 15712 12189
rect 15752 12180 15804 12232
rect 21088 12180 21140 12232
rect 11244 12112 11296 12164
rect 2780 12087 2832 12096
rect 2780 12053 2789 12087
rect 2789 12053 2823 12087
rect 2823 12053 2832 12087
rect 2780 12044 2832 12053
rect 5356 12087 5408 12096
rect 5356 12053 5365 12087
rect 5365 12053 5399 12087
rect 5399 12053 5408 12087
rect 5356 12044 5408 12053
rect 5724 12087 5776 12096
rect 5724 12053 5733 12087
rect 5733 12053 5767 12087
rect 5767 12053 5776 12087
rect 5724 12044 5776 12053
rect 6092 12087 6144 12096
rect 6092 12053 6101 12087
rect 6101 12053 6135 12087
rect 6135 12053 6144 12087
rect 6092 12044 6144 12053
rect 7288 12087 7340 12096
rect 7288 12053 7297 12087
rect 7297 12053 7331 12087
rect 7331 12053 7340 12087
rect 7288 12044 7340 12053
rect 7656 12044 7708 12096
rect 8484 12044 8536 12096
rect 9772 12044 9824 12096
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 11888 12087 11940 12096
rect 11888 12053 11897 12087
rect 11897 12053 11931 12087
rect 11931 12053 11940 12087
rect 11888 12044 11940 12053
rect 16948 12087 17000 12096
rect 16948 12053 16957 12087
rect 16957 12053 16991 12087
rect 16991 12053 17000 12087
rect 16948 12044 17000 12053
rect 18328 12087 18380 12096
rect 18328 12053 18337 12087
rect 18337 12053 18371 12087
rect 18371 12053 18380 12087
rect 18328 12044 18380 12053
rect 4982 11942 5034 11994
rect 5046 11942 5098 11994
rect 5110 11942 5162 11994
rect 5174 11942 5226 11994
rect 12982 11942 13034 11994
rect 13046 11942 13098 11994
rect 13110 11942 13162 11994
rect 13174 11942 13226 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 4620 11840 4672 11892
rect 8392 11840 8444 11892
rect 10048 11840 10100 11892
rect 11888 11840 11940 11892
rect 19616 11883 19668 11892
rect 19616 11849 19625 11883
rect 19625 11849 19659 11883
rect 19659 11849 19668 11883
rect 19616 11840 19668 11849
rect 20812 11883 20864 11892
rect 20812 11849 20821 11883
rect 20821 11849 20855 11883
rect 20855 11849 20864 11883
rect 20812 11840 20864 11849
rect 21732 11883 21784 11892
rect 21732 11849 21741 11883
rect 21741 11849 21775 11883
rect 21775 11849 21784 11883
rect 21732 11840 21784 11849
rect 4804 11772 4856 11824
rect 1124 11704 1176 11756
rect 4712 11704 4764 11756
rect 10232 11772 10284 11824
rect 14188 11772 14240 11824
rect 10416 11747 10468 11756
rect 10416 11713 10425 11747
rect 10425 11713 10459 11747
rect 10459 11713 10468 11747
rect 10416 11704 10468 11713
rect 2780 11636 2832 11688
rect 4160 11636 4212 11688
rect 5356 11679 5408 11688
rect 5356 11645 5362 11679
rect 5362 11645 5408 11679
rect 5356 11636 5408 11645
rect 6368 11636 6420 11688
rect 7104 11679 7156 11688
rect 7104 11645 7113 11679
rect 7113 11645 7147 11679
rect 7147 11645 7156 11679
rect 7104 11636 7156 11645
rect 7288 11636 7340 11688
rect 7840 11679 7892 11688
rect 7840 11645 7849 11679
rect 7849 11645 7883 11679
rect 7883 11645 7892 11679
rect 7840 11636 7892 11645
rect 9680 11636 9732 11688
rect 10784 11636 10836 11688
rect 11244 11636 11296 11688
rect 14004 11679 14056 11688
rect 14004 11645 14013 11679
rect 14013 11645 14047 11679
rect 14047 11645 14056 11679
rect 14004 11636 14056 11645
rect 16948 11772 17000 11824
rect 21456 11815 21508 11824
rect 21456 11781 21465 11815
rect 21465 11781 21499 11815
rect 21499 11781 21508 11815
rect 21456 11772 21508 11781
rect 15660 11704 15712 11756
rect 1676 11500 1728 11552
rect 3608 11543 3660 11552
rect 3608 11509 3617 11543
rect 3617 11509 3651 11543
rect 3651 11509 3660 11543
rect 3608 11500 3660 11509
rect 5724 11568 5776 11620
rect 10048 11611 10100 11620
rect 4436 11500 4488 11552
rect 4712 11543 4764 11552
rect 4712 11509 4721 11543
rect 4721 11509 4755 11543
rect 4755 11509 4764 11543
rect 4712 11500 4764 11509
rect 6276 11543 6328 11552
rect 6276 11509 6285 11543
rect 6285 11509 6319 11543
rect 6319 11509 6328 11543
rect 6276 11500 6328 11509
rect 6460 11500 6512 11552
rect 7840 11500 7892 11552
rect 9680 11543 9732 11552
rect 9680 11509 9689 11543
rect 9689 11509 9723 11543
rect 9723 11509 9732 11543
rect 9680 11500 9732 11509
rect 10048 11577 10057 11611
rect 10057 11577 10091 11611
rect 10091 11577 10100 11611
rect 10048 11568 10100 11577
rect 13544 11568 13596 11620
rect 10416 11500 10468 11552
rect 10968 11500 11020 11552
rect 11520 11500 11572 11552
rect 12716 11543 12768 11552
rect 12716 11509 12725 11543
rect 12725 11509 12759 11543
rect 12759 11509 12768 11543
rect 12716 11500 12768 11509
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 17868 11636 17920 11688
rect 18328 11679 18380 11688
rect 18328 11645 18337 11679
rect 18337 11645 18371 11679
rect 18371 11645 18380 11679
rect 18328 11636 18380 11645
rect 16212 11611 16264 11620
rect 16212 11577 16221 11611
rect 16221 11577 16255 11611
rect 16255 11577 16264 11611
rect 16212 11568 16264 11577
rect 18420 11568 18472 11620
rect 8982 11398 9034 11450
rect 9046 11398 9098 11450
rect 9110 11398 9162 11450
rect 9174 11398 9226 11450
rect 16982 11398 17034 11450
rect 17046 11398 17098 11450
rect 17110 11398 17162 11450
rect 17174 11398 17226 11450
rect 1676 11296 1728 11348
rect 4160 11339 4212 11348
rect 4160 11305 4169 11339
rect 4169 11305 4203 11339
rect 4203 11305 4212 11339
rect 4160 11296 4212 11305
rect 4712 11296 4764 11348
rect 5356 11296 5408 11348
rect 6552 11339 6604 11348
rect 6552 11305 6561 11339
rect 6561 11305 6595 11339
rect 6595 11305 6604 11339
rect 6552 11296 6604 11305
rect 7380 11339 7432 11348
rect 7380 11305 7389 11339
rect 7389 11305 7423 11339
rect 7423 11305 7432 11339
rect 7380 11296 7432 11305
rect 10232 11339 10284 11348
rect 10232 11305 10241 11339
rect 10241 11305 10275 11339
rect 10275 11305 10284 11339
rect 10232 11296 10284 11305
rect 1860 11228 1912 11280
rect 4068 11228 4120 11280
rect 5724 11228 5776 11280
rect 7104 11228 7156 11280
rect 8760 11271 8812 11280
rect 8760 11237 8769 11271
rect 8769 11237 8803 11271
rect 8803 11237 8812 11271
rect 8760 11228 8812 11237
rect 4344 11203 4396 11212
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 4528 11203 4580 11212
rect 4528 11169 4537 11203
rect 4537 11169 4571 11203
rect 4571 11169 4580 11203
rect 4528 11160 4580 11169
rect 6368 11160 6420 11212
rect 7840 11160 7892 11212
rect 11520 11228 11572 11280
rect 11704 11271 11756 11280
rect 11704 11237 11713 11271
rect 11713 11237 11747 11271
rect 11747 11237 11756 11271
rect 11704 11228 11756 11237
rect 9404 11160 9456 11212
rect 10048 11160 10100 11212
rect 10692 11160 10744 11212
rect 1952 11092 2004 11144
rect 6276 11135 6328 11144
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6276 11092 6328 11101
rect 7932 11092 7984 11144
rect 1768 11024 1820 11076
rect 2596 11024 2648 11076
rect 6736 11024 6788 11076
rect 6920 11024 6972 11076
rect 12532 11160 12584 11212
rect 18420 11339 18472 11348
rect 18420 11305 18429 11339
rect 18429 11305 18463 11339
rect 18463 11305 18472 11339
rect 18420 11296 18472 11305
rect 13452 11228 13504 11280
rect 17868 11271 17920 11280
rect 17868 11237 17877 11271
rect 17877 11237 17911 11271
rect 17911 11237 17920 11271
rect 17868 11228 17920 11237
rect 14004 11203 14056 11212
rect 14004 11169 14013 11203
rect 14013 11169 14047 11203
rect 14047 11169 14056 11203
rect 14004 11160 14056 11169
rect 15384 11203 15436 11212
rect 15384 11169 15393 11203
rect 15393 11169 15427 11203
rect 15427 11169 15436 11203
rect 15384 11160 15436 11169
rect 15844 11203 15896 11212
rect 15844 11169 15853 11203
rect 15853 11169 15887 11203
rect 15887 11169 15896 11203
rect 15844 11160 15896 11169
rect 17592 11203 17644 11212
rect 11060 11092 11112 11144
rect 17592 11169 17601 11203
rect 17601 11169 17635 11203
rect 17635 11169 17644 11203
rect 17592 11160 17644 11169
rect 17500 11092 17552 11144
rect 5448 10956 5500 11008
rect 6092 10956 6144 11008
rect 6552 10956 6604 11008
rect 7104 10999 7156 11008
rect 7104 10965 7113 10999
rect 7113 10965 7147 10999
rect 7147 10965 7156 10999
rect 7104 10956 7156 10965
rect 8024 10956 8076 11008
rect 8208 10999 8260 11008
rect 8208 10965 8232 10999
rect 8232 10965 8260 10999
rect 8208 10956 8260 10965
rect 8484 10956 8536 11008
rect 9404 10999 9456 11008
rect 9404 10965 9413 10999
rect 9413 10965 9447 10999
rect 9447 10965 9456 10999
rect 9404 10956 9456 10965
rect 10784 10956 10836 11008
rect 11244 10999 11296 11008
rect 11244 10965 11253 10999
rect 11253 10965 11287 10999
rect 11287 10965 11296 10999
rect 11244 10956 11296 10965
rect 11336 10956 11388 11008
rect 4982 10854 5034 10906
rect 5046 10854 5098 10906
rect 5110 10854 5162 10906
rect 5174 10854 5226 10906
rect 12982 10854 13034 10906
rect 13046 10854 13098 10906
rect 13110 10854 13162 10906
rect 13174 10854 13226 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 4528 10752 4580 10804
rect 4804 10752 4856 10804
rect 2596 10727 2648 10736
rect 2596 10693 2605 10727
rect 2605 10693 2639 10727
rect 2639 10693 2648 10727
rect 2596 10684 2648 10693
rect 5632 10752 5684 10804
rect 6552 10795 6604 10804
rect 6552 10761 6561 10795
rect 6561 10761 6595 10795
rect 6595 10761 6604 10795
rect 6552 10752 6604 10761
rect 8484 10752 8536 10804
rect 13452 10795 13504 10804
rect 13452 10761 13461 10795
rect 13461 10761 13495 10795
rect 13495 10761 13504 10795
rect 13452 10752 13504 10761
rect 14004 10752 14056 10804
rect 14188 10752 14240 10804
rect 15384 10752 15436 10804
rect 1860 10659 1912 10668
rect 1860 10625 1869 10659
rect 1869 10625 1903 10659
rect 1903 10625 1912 10659
rect 1860 10616 1912 10625
rect 4344 10616 4396 10668
rect 5356 10616 5408 10668
rect 7932 10684 7984 10736
rect 10968 10727 11020 10736
rect 10968 10693 10977 10727
rect 10977 10693 11011 10727
rect 11011 10693 11020 10727
rect 10968 10684 11020 10693
rect 3608 10591 3660 10600
rect 2044 10523 2096 10532
rect 2044 10489 2053 10523
rect 2053 10489 2087 10523
rect 2087 10489 2096 10523
rect 2044 10480 2096 10489
rect 3608 10557 3617 10591
rect 3617 10557 3651 10591
rect 3651 10557 3660 10591
rect 3608 10548 3660 10557
rect 4252 10548 4304 10600
rect 9404 10616 9456 10668
rect 7748 10591 7800 10600
rect 7748 10557 7757 10591
rect 7757 10557 7791 10591
rect 7791 10557 7800 10591
rect 7748 10548 7800 10557
rect 5540 10480 5592 10532
rect 7840 10480 7892 10532
rect 6276 10455 6328 10464
rect 6276 10421 6285 10455
rect 6285 10421 6319 10455
rect 6319 10421 6328 10455
rect 6276 10412 6328 10421
rect 8024 10412 8076 10464
rect 12164 10548 12216 10600
rect 9588 10523 9640 10532
rect 9588 10489 9597 10523
rect 9597 10489 9631 10523
rect 9631 10489 9640 10523
rect 9588 10480 9640 10489
rect 11244 10480 11296 10532
rect 9772 10412 9824 10464
rect 10784 10412 10836 10464
rect 11704 10412 11756 10464
rect 11888 10412 11940 10464
rect 15844 10684 15896 10736
rect 17592 10684 17644 10736
rect 12440 10616 12492 10668
rect 13360 10616 13412 10668
rect 14188 10616 14240 10668
rect 14372 10659 14424 10668
rect 14372 10625 14381 10659
rect 14381 10625 14415 10659
rect 14415 10625 14424 10659
rect 14372 10616 14424 10625
rect 12716 10548 12768 10600
rect 19156 10548 19208 10600
rect 20628 10591 20680 10600
rect 20628 10557 20637 10591
rect 20637 10557 20671 10591
rect 20671 10557 20680 10591
rect 20628 10548 20680 10557
rect 22100 10548 22152 10600
rect 14096 10523 14148 10532
rect 14096 10489 14105 10523
rect 14105 10489 14139 10523
rect 14139 10489 14148 10523
rect 14096 10480 14148 10489
rect 12532 10412 12584 10464
rect 14004 10412 14056 10464
rect 14464 10412 14516 10464
rect 17500 10412 17552 10464
rect 20260 10455 20312 10464
rect 20260 10421 20269 10455
rect 20269 10421 20303 10455
rect 20303 10421 20312 10455
rect 20260 10412 20312 10421
rect 20536 10412 20588 10464
rect 22100 10455 22152 10464
rect 22100 10421 22109 10455
rect 22109 10421 22143 10455
rect 22143 10421 22152 10455
rect 22100 10412 22152 10421
rect 8982 10310 9034 10362
rect 9046 10310 9098 10362
rect 9110 10310 9162 10362
rect 9174 10310 9226 10362
rect 16982 10310 17034 10362
rect 17046 10310 17098 10362
rect 17110 10310 17162 10362
rect 17174 10310 17226 10362
rect 2044 10208 2096 10260
rect 3608 10251 3660 10260
rect 3608 10217 3617 10251
rect 3617 10217 3651 10251
rect 3651 10217 3660 10251
rect 3608 10208 3660 10217
rect 4068 10208 4120 10260
rect 5540 10208 5592 10260
rect 5632 10251 5684 10260
rect 5632 10217 5641 10251
rect 5641 10217 5675 10251
rect 5675 10217 5684 10251
rect 5632 10208 5684 10217
rect 7748 10208 7800 10260
rect 12716 10208 12768 10260
rect 13452 10208 13504 10260
rect 13912 10208 13964 10260
rect 14096 10208 14148 10260
rect 15752 10208 15804 10260
rect 3792 10140 3844 10192
rect 4160 10140 4212 10192
rect 2044 10072 2096 10124
rect 4344 10115 4396 10124
rect 4344 10081 4353 10115
rect 4353 10081 4387 10115
rect 4387 10081 4396 10115
rect 4344 10072 4396 10081
rect 5816 10115 5868 10124
rect 5816 10081 5825 10115
rect 5825 10081 5859 10115
rect 5859 10081 5868 10115
rect 5816 10072 5868 10081
rect 7104 10072 7156 10124
rect 8668 10140 8720 10192
rect 9588 10140 9640 10192
rect 13820 10183 13872 10192
rect 13820 10149 13829 10183
rect 13829 10149 13863 10183
rect 13863 10149 13872 10183
rect 14372 10183 14424 10192
rect 13820 10140 13872 10149
rect 14372 10149 14381 10183
rect 14381 10149 14415 10183
rect 14415 10149 14424 10183
rect 14372 10140 14424 10149
rect 20628 10140 20680 10192
rect 21456 10140 21508 10192
rect 7288 10072 7340 10124
rect 7748 10072 7800 10124
rect 7932 10072 7984 10124
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 10232 10072 10284 10124
rect 11796 10072 11848 10124
rect 15936 10115 15988 10124
rect 15936 10081 15945 10115
rect 15945 10081 15979 10115
rect 15979 10081 15988 10115
rect 15936 10072 15988 10081
rect 17592 10115 17644 10124
rect 2136 10047 2188 10056
rect 2136 10013 2145 10047
rect 2145 10013 2179 10047
rect 2179 10013 2188 10047
rect 2136 10004 2188 10013
rect 6368 10004 6420 10056
rect 8208 10004 8260 10056
rect 8576 10004 8628 10056
rect 1952 9936 2004 9988
rect 6828 9936 6880 9988
rect 8484 9936 8536 9988
rect 11060 10004 11112 10056
rect 11244 10047 11296 10056
rect 11244 10013 11253 10047
rect 11253 10013 11287 10047
rect 11287 10013 11296 10047
rect 11244 10004 11296 10013
rect 12164 10004 12216 10056
rect 11428 9936 11480 9988
rect 14464 10004 14516 10056
rect 15384 10047 15436 10056
rect 15384 10013 15393 10047
rect 15393 10013 15427 10047
rect 15427 10013 15436 10047
rect 15384 10004 15436 10013
rect 17592 10081 17601 10115
rect 17601 10081 17635 10115
rect 17635 10081 17644 10115
rect 17592 10072 17644 10081
rect 17500 10004 17552 10056
rect 17868 10047 17920 10056
rect 17868 10013 17877 10047
rect 17877 10013 17911 10047
rect 17911 10013 17920 10047
rect 17868 10004 17920 10013
rect 21824 10004 21876 10056
rect 5724 9868 5776 9920
rect 6368 9911 6420 9920
rect 6368 9877 6377 9911
rect 6377 9877 6411 9911
rect 6411 9877 6420 9911
rect 6368 9868 6420 9877
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 14372 9936 14424 9988
rect 21548 9979 21600 9988
rect 21548 9945 21557 9979
rect 21557 9945 21591 9979
rect 21591 9945 21600 9979
rect 21548 9936 21600 9945
rect 13636 9868 13688 9920
rect 4982 9766 5034 9818
rect 5046 9766 5098 9818
rect 5110 9766 5162 9818
rect 5174 9766 5226 9818
rect 12982 9766 13034 9818
rect 13046 9766 13098 9818
rect 13110 9766 13162 9818
rect 13174 9766 13226 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 2136 9707 2188 9716
rect 2136 9673 2145 9707
rect 2145 9673 2179 9707
rect 2179 9673 2188 9707
rect 2136 9664 2188 9673
rect 3792 9707 3844 9716
rect 3792 9673 3801 9707
rect 3801 9673 3835 9707
rect 3835 9673 3844 9707
rect 3792 9664 3844 9673
rect 4344 9664 4396 9716
rect 5816 9707 5868 9716
rect 5816 9673 5825 9707
rect 5825 9673 5859 9707
rect 5859 9673 5868 9707
rect 5816 9664 5868 9673
rect 7288 9664 7340 9716
rect 9772 9664 9824 9716
rect 10416 9664 10468 9716
rect 11060 9707 11112 9716
rect 2320 9596 2372 9648
rect 7564 9596 7616 9648
rect 7932 9596 7984 9648
rect 11060 9673 11069 9707
rect 11069 9673 11103 9707
rect 11103 9673 11112 9707
rect 11060 9664 11112 9673
rect 11428 9707 11480 9716
rect 11428 9673 11437 9707
rect 11437 9673 11471 9707
rect 11471 9673 11480 9707
rect 11428 9664 11480 9673
rect 11796 9707 11848 9716
rect 11796 9673 11805 9707
rect 11805 9673 11839 9707
rect 11839 9673 11848 9707
rect 11796 9664 11848 9673
rect 12164 9707 12216 9716
rect 12164 9673 12173 9707
rect 12173 9673 12207 9707
rect 12207 9673 12216 9707
rect 12164 9664 12216 9673
rect 13820 9664 13872 9716
rect 19156 9707 19208 9716
rect 19156 9673 19165 9707
rect 19165 9673 19199 9707
rect 19199 9673 19208 9707
rect 19156 9664 19208 9673
rect 20260 9707 20312 9716
rect 20260 9673 20269 9707
rect 20269 9673 20303 9707
rect 20303 9673 20312 9707
rect 20260 9664 20312 9673
rect 21456 9707 21508 9716
rect 21456 9673 21465 9707
rect 21465 9673 21499 9707
rect 21499 9673 21508 9707
rect 21456 9664 21508 9673
rect 21824 9707 21876 9716
rect 21824 9673 21833 9707
rect 21833 9673 21867 9707
rect 21867 9673 21876 9707
rect 21824 9664 21876 9673
rect 3424 9528 3476 9580
rect 4068 9528 4120 9580
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 9404 9528 9456 9580
rect 10784 9528 10836 9580
rect 12440 9596 12492 9648
rect 13912 9596 13964 9648
rect 15844 9596 15896 9648
rect 4620 9503 4672 9512
rect 4620 9469 4629 9503
rect 4629 9469 4663 9503
rect 4663 9469 4672 9503
rect 4620 9460 4672 9469
rect 8484 9435 8536 9444
rect 2044 9324 2096 9376
rect 2136 9324 2188 9376
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 4436 9367 4488 9376
rect 4436 9333 4445 9367
rect 4445 9333 4479 9367
rect 4479 9333 4488 9367
rect 8484 9401 8493 9435
rect 8493 9401 8527 9435
rect 8527 9401 8536 9435
rect 8484 9392 8536 9401
rect 8576 9435 8628 9444
rect 8576 9401 8585 9435
rect 8585 9401 8619 9435
rect 8619 9401 8628 9435
rect 8576 9392 8628 9401
rect 11244 9392 11296 9444
rect 4436 9324 4488 9333
rect 5264 9324 5316 9376
rect 7748 9367 7800 9376
rect 7748 9333 7757 9367
rect 7757 9333 7791 9367
rect 7791 9333 7800 9367
rect 7748 9324 7800 9333
rect 10508 9324 10560 9376
rect 13360 9460 13412 9512
rect 13636 9503 13688 9512
rect 13636 9469 13645 9503
rect 13645 9469 13679 9503
rect 13679 9469 13688 9503
rect 17592 9528 17644 9580
rect 17868 9528 17920 9580
rect 18236 9571 18288 9580
rect 18236 9537 18245 9571
rect 18245 9537 18279 9571
rect 18279 9537 18288 9571
rect 18236 9528 18288 9537
rect 20536 9571 20588 9580
rect 20536 9537 20545 9571
rect 20545 9537 20579 9571
rect 20579 9537 20588 9571
rect 20536 9528 20588 9537
rect 21548 9528 21600 9580
rect 13636 9460 13688 9469
rect 14740 9503 14792 9512
rect 14740 9469 14749 9503
rect 14749 9469 14783 9503
rect 14783 9469 14792 9503
rect 14740 9460 14792 9469
rect 14832 9392 14884 9444
rect 18788 9392 18840 9444
rect 15936 9367 15988 9376
rect 15936 9333 15945 9367
rect 15945 9333 15979 9367
rect 15979 9333 15988 9367
rect 15936 9324 15988 9333
rect 16488 9367 16540 9376
rect 16488 9333 16497 9367
rect 16497 9333 16531 9367
rect 16531 9333 16540 9367
rect 16488 9324 16540 9333
rect 17500 9324 17552 9376
rect 20260 9324 20312 9376
rect 8982 9222 9034 9274
rect 9046 9222 9098 9274
rect 9110 9222 9162 9274
rect 9174 9222 9226 9274
rect 16982 9222 17034 9274
rect 17046 9222 17098 9274
rect 17110 9222 17162 9274
rect 17174 9222 17226 9274
rect 112 9120 164 9172
rect 4620 9163 4672 9172
rect 4620 9129 4629 9163
rect 4629 9129 4663 9163
rect 4663 9129 4672 9163
rect 4620 9120 4672 9129
rect 5264 9163 5316 9172
rect 5264 9129 5273 9163
rect 5273 9129 5307 9163
rect 5307 9129 5316 9163
rect 5264 9120 5316 9129
rect 2044 9095 2096 9104
rect 2044 9061 2053 9095
rect 2053 9061 2087 9095
rect 2087 9061 2096 9095
rect 2044 9052 2096 9061
rect 6920 9120 6972 9172
rect 8484 9120 8536 9172
rect 10876 9120 10928 9172
rect 14464 9120 14516 9172
rect 14740 9163 14792 9172
rect 14740 9129 14749 9163
rect 14749 9129 14783 9163
rect 14783 9129 14792 9163
rect 14740 9120 14792 9129
rect 15660 9163 15712 9172
rect 15660 9129 15669 9163
rect 15669 9129 15703 9163
rect 15703 9129 15712 9163
rect 15660 9120 15712 9129
rect 16488 9120 16540 9172
rect 17592 9120 17644 9172
rect 18236 9163 18288 9172
rect 18236 9129 18245 9163
rect 18245 9129 18279 9163
rect 18279 9129 18288 9163
rect 18236 9120 18288 9129
rect 20536 9163 20588 9172
rect 20536 9129 20545 9163
rect 20545 9129 20579 9163
rect 20579 9129 20588 9163
rect 20536 9120 20588 9129
rect 3884 8984 3936 9036
rect 6092 9052 6144 9104
rect 13360 9095 13412 9104
rect 13360 9061 13369 9095
rect 13369 9061 13403 9095
rect 13403 9061 13412 9095
rect 13360 9052 13412 9061
rect 15936 9095 15988 9104
rect 15936 9061 15945 9095
rect 15945 9061 15979 9095
rect 15979 9061 15988 9095
rect 15936 9052 15988 9061
rect 16580 9052 16632 9104
rect 7932 8984 7984 9036
rect 9680 8984 9732 9036
rect 10600 8984 10652 9036
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 10508 8916 10560 8968
rect 2320 8848 2372 8900
rect 2872 8848 2924 8900
rect 5724 8848 5776 8900
rect 5908 8848 5960 8900
rect 11980 8984 12032 9036
rect 21456 8984 21508 9036
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 14556 8916 14608 8968
rect 15844 8959 15896 8968
rect 15844 8925 15853 8959
rect 15853 8925 15887 8959
rect 15887 8925 15896 8959
rect 15844 8916 15896 8925
rect 16212 8959 16264 8968
rect 16212 8925 16221 8959
rect 16221 8925 16255 8959
rect 16255 8925 16264 8959
rect 16212 8916 16264 8925
rect 13544 8848 13596 8900
rect 13820 8891 13872 8900
rect 13820 8857 13829 8891
rect 13829 8857 13863 8891
rect 13863 8857 13872 8891
rect 13820 8848 13872 8857
rect 17224 8848 17276 8900
rect 1400 8780 1452 8832
rect 6644 8780 6696 8832
rect 7840 8823 7892 8832
rect 7840 8789 7849 8823
rect 7849 8789 7883 8823
rect 7883 8789 7892 8823
rect 7840 8780 7892 8789
rect 4982 8678 5034 8730
rect 5046 8678 5098 8730
rect 5110 8678 5162 8730
rect 5174 8678 5226 8730
rect 12982 8678 13034 8730
rect 13046 8678 13098 8730
rect 13110 8678 13162 8730
rect 13174 8678 13226 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 2872 8576 2924 8628
rect 2044 8551 2096 8560
rect 2044 8517 2053 8551
rect 2053 8517 2087 8551
rect 2087 8517 2096 8551
rect 5632 8576 5684 8628
rect 10600 8619 10652 8628
rect 10600 8585 10609 8619
rect 10609 8585 10643 8619
rect 10643 8585 10652 8619
rect 10600 8576 10652 8585
rect 14556 8619 14608 8628
rect 14556 8585 14565 8619
rect 14565 8585 14599 8619
rect 14599 8585 14608 8619
rect 14556 8576 14608 8585
rect 15384 8619 15436 8628
rect 15384 8585 15393 8619
rect 15393 8585 15427 8619
rect 15427 8585 15436 8619
rect 15384 8576 15436 8585
rect 16580 8619 16632 8628
rect 16580 8585 16589 8619
rect 16589 8585 16623 8619
rect 16623 8585 16632 8619
rect 16580 8576 16632 8585
rect 21456 8619 21508 8628
rect 21456 8585 21465 8619
rect 21465 8585 21499 8619
rect 21499 8585 21508 8619
rect 21456 8576 21508 8585
rect 2044 8508 2096 8517
rect 3148 8508 3200 8560
rect 3608 8440 3660 8492
rect 8300 8508 8352 8560
rect 9404 8508 9456 8560
rect 11980 8551 12032 8560
rect 11980 8517 11989 8551
rect 11989 8517 12023 8551
rect 12023 8517 12032 8551
rect 11980 8508 12032 8517
rect 13820 8508 13872 8560
rect 16212 8551 16264 8560
rect 16212 8517 16221 8551
rect 16221 8517 16255 8551
rect 16255 8517 16264 8551
rect 16212 8508 16264 8517
rect 13268 8440 13320 8492
rect 13452 8440 13504 8492
rect 15660 8483 15712 8492
rect 15660 8449 15669 8483
rect 15669 8449 15703 8483
rect 15703 8449 15712 8483
rect 15660 8440 15712 8449
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 7840 8372 7892 8424
rect 22192 8576 22244 8628
rect 112 8236 164 8288
rect 3056 8279 3108 8288
rect 3056 8245 3065 8279
rect 3065 8245 3099 8279
rect 3099 8245 3108 8279
rect 4436 8304 4488 8356
rect 5356 8347 5408 8356
rect 5356 8313 5365 8347
rect 5365 8313 5399 8347
rect 5399 8313 5408 8347
rect 5356 8304 5408 8313
rect 5908 8347 5960 8356
rect 5908 8313 5917 8347
rect 5917 8313 5951 8347
rect 5951 8313 5960 8347
rect 5908 8304 5960 8313
rect 8024 8304 8076 8356
rect 9680 8347 9732 8356
rect 9680 8313 9689 8347
rect 9689 8313 9723 8347
rect 9723 8313 9732 8347
rect 9680 8304 9732 8313
rect 13728 8347 13780 8356
rect 13728 8313 13737 8347
rect 13737 8313 13771 8347
rect 13771 8313 13780 8347
rect 13728 8304 13780 8313
rect 6184 8279 6236 8288
rect 3056 8236 3108 8245
rect 6184 8245 6193 8279
rect 6193 8245 6227 8279
rect 6227 8245 6236 8279
rect 6184 8236 6236 8245
rect 8668 8279 8720 8288
rect 8668 8245 8677 8279
rect 8677 8245 8711 8279
rect 8711 8245 8720 8279
rect 8668 8236 8720 8245
rect 13360 8236 13412 8288
rect 15016 8279 15068 8288
rect 15016 8245 15025 8279
rect 15025 8245 15059 8279
rect 15059 8245 15068 8279
rect 15016 8236 15068 8245
rect 15384 8236 15436 8288
rect 16304 8236 16356 8288
rect 8982 8134 9034 8186
rect 9046 8134 9098 8186
rect 9110 8134 9162 8186
rect 9174 8134 9226 8186
rect 16982 8134 17034 8186
rect 17046 8134 17098 8186
rect 17110 8134 17162 8186
rect 17174 8134 17226 8186
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 7840 8075 7892 8084
rect 7840 8041 7849 8075
rect 7849 8041 7883 8075
rect 7883 8041 7892 8075
rect 7840 8032 7892 8041
rect 13452 8032 13504 8084
rect 15016 8032 15068 8084
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 17408 8032 17460 8084
rect 2412 7964 2464 8016
rect 6184 7964 6236 8016
rect 9680 8007 9732 8016
rect 9680 7973 9689 8007
rect 9689 7973 9723 8007
rect 9723 7973 9732 8007
rect 9680 7964 9732 7973
rect 12624 7964 12676 8016
rect 5356 7939 5408 7948
rect 2320 7828 2372 7880
rect 2504 7871 2556 7880
rect 2504 7837 2513 7871
rect 2513 7837 2547 7871
rect 2547 7837 2556 7871
rect 5356 7905 5365 7939
rect 5365 7905 5399 7939
rect 5399 7905 5408 7939
rect 5356 7896 5408 7905
rect 2504 7828 2556 7837
rect 7288 7896 7340 7948
rect 7564 7896 7616 7948
rect 9772 7939 9824 7948
rect 9772 7905 9781 7939
rect 9781 7905 9815 7939
rect 9815 7905 9824 7939
rect 9772 7896 9824 7905
rect 15384 7939 15436 7948
rect 15384 7905 15402 7939
rect 15402 7905 15436 7939
rect 15384 7896 15436 7905
rect 16212 7896 16264 7948
rect 21364 7896 21416 7948
rect 7472 7828 7524 7880
rect 12808 7828 12860 7880
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 1952 7735 2004 7744
rect 1952 7701 1961 7735
rect 1961 7701 1995 7735
rect 1995 7701 2004 7735
rect 1952 7692 2004 7701
rect 3608 7692 3660 7744
rect 3700 7692 3752 7744
rect 8852 7735 8904 7744
rect 8852 7701 8861 7735
rect 8861 7701 8895 7735
rect 8895 7701 8904 7735
rect 8852 7692 8904 7701
rect 10784 7735 10836 7744
rect 10784 7701 10793 7735
rect 10793 7701 10827 7735
rect 10827 7701 10836 7735
rect 10784 7692 10836 7701
rect 13636 7692 13688 7744
rect 14096 7735 14148 7744
rect 14096 7701 14105 7735
rect 14105 7701 14139 7735
rect 14139 7701 14148 7735
rect 14096 7692 14148 7701
rect 15568 7692 15620 7744
rect 4982 7590 5034 7642
rect 5046 7590 5098 7642
rect 5110 7590 5162 7642
rect 5174 7590 5226 7642
rect 12982 7590 13034 7642
rect 13046 7590 13098 7642
rect 13110 7590 13162 7642
rect 13174 7590 13226 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 2412 7488 2464 7540
rect 5724 7488 5776 7540
rect 7288 7488 7340 7540
rect 8668 7531 8720 7540
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 8668 7488 8720 7497
rect 8944 7488 8996 7540
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 10968 7488 11020 7540
rect 15384 7531 15436 7540
rect 5448 7463 5500 7472
rect 5448 7429 5457 7463
rect 5457 7429 5491 7463
rect 5491 7429 5500 7463
rect 5448 7420 5500 7429
rect 7748 7420 7800 7472
rect 9404 7463 9456 7472
rect 9404 7429 9413 7463
rect 9413 7429 9447 7463
rect 9447 7429 9456 7463
rect 9404 7420 9456 7429
rect 10600 7420 10652 7472
rect 2504 7352 2556 7404
rect 6276 7352 6328 7404
rect 7564 7352 7616 7404
rect 8668 7352 8720 7404
rect 10784 7352 10836 7404
rect 15384 7497 15393 7531
rect 15393 7497 15427 7531
rect 15427 7497 15436 7531
rect 15384 7488 15436 7497
rect 21364 7488 21416 7540
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 1676 7259 1728 7268
rect 1676 7225 1685 7259
rect 1685 7225 1719 7259
rect 1719 7225 1728 7259
rect 1676 7216 1728 7225
rect 1768 7259 1820 7268
rect 1768 7225 1777 7259
rect 1777 7225 1811 7259
rect 1811 7225 1820 7259
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 17960 7352 18012 7404
rect 1768 7216 1820 7225
rect 8852 7259 8904 7268
rect 3056 7191 3108 7200
rect 3056 7157 3065 7191
rect 3065 7157 3099 7191
rect 3099 7157 3108 7191
rect 8852 7225 8861 7259
rect 8861 7225 8895 7259
rect 8895 7225 8904 7259
rect 8852 7216 8904 7225
rect 8944 7259 8996 7268
rect 8944 7225 8953 7259
rect 8953 7225 8987 7259
rect 8987 7225 8996 7259
rect 8944 7216 8996 7225
rect 3056 7148 3108 7157
rect 4712 7148 4764 7200
rect 5080 7148 5132 7200
rect 6644 7191 6696 7200
rect 6644 7157 6653 7191
rect 6653 7157 6687 7191
rect 6687 7157 6696 7191
rect 6644 7148 6696 7157
rect 7472 7148 7524 7200
rect 11244 7216 11296 7268
rect 13544 7216 13596 7268
rect 14096 7284 14148 7336
rect 14740 7259 14792 7268
rect 10600 7191 10652 7200
rect 10600 7157 10609 7191
rect 10609 7157 10643 7191
rect 10643 7157 10652 7191
rect 10600 7148 10652 7157
rect 12624 7148 12676 7200
rect 12808 7148 12860 7200
rect 14740 7225 14749 7259
rect 14749 7225 14783 7259
rect 14783 7225 14792 7259
rect 14740 7216 14792 7225
rect 17500 7148 17552 7200
rect 19340 7284 19392 7336
rect 21272 7284 21324 7336
rect 18328 7191 18380 7200
rect 18328 7157 18337 7191
rect 18337 7157 18371 7191
rect 18371 7157 18380 7191
rect 18328 7148 18380 7157
rect 20352 7191 20404 7200
rect 20352 7157 20361 7191
rect 20361 7157 20395 7191
rect 20395 7157 20404 7191
rect 20352 7148 20404 7157
rect 8982 7046 9034 7098
rect 9046 7046 9098 7098
rect 9110 7046 9162 7098
rect 9174 7046 9226 7098
rect 16982 7046 17034 7098
rect 17046 7046 17098 7098
rect 17110 7046 17162 7098
rect 17174 7046 17226 7098
rect 2320 6944 2372 6996
rect 3148 6944 3200 6996
rect 5448 6944 5500 6996
rect 7288 6987 7340 6996
rect 7288 6953 7297 6987
rect 7297 6953 7331 6987
rect 7331 6953 7340 6987
rect 7288 6944 7340 6953
rect 7656 6944 7708 6996
rect 7472 6876 7524 6928
rect 1768 6851 1820 6860
rect 1768 6817 1777 6851
rect 1777 6817 1811 6851
rect 1811 6817 1820 6851
rect 1768 6808 1820 6817
rect 2412 6851 2464 6860
rect 2412 6817 2421 6851
rect 2421 6817 2455 6851
rect 2455 6817 2464 6851
rect 2412 6808 2464 6817
rect 4344 6851 4396 6860
rect 4344 6817 4353 6851
rect 4353 6817 4387 6851
rect 4387 6817 4396 6851
rect 4344 6808 4396 6817
rect 4252 6740 4304 6792
rect 5080 6808 5132 6860
rect 5724 6808 5776 6860
rect 6644 6808 6696 6860
rect 4712 6740 4764 6792
rect 10968 6944 11020 6996
rect 11612 6944 11664 6996
rect 12808 6987 12860 6996
rect 12808 6953 12817 6987
rect 12817 6953 12851 6987
rect 12851 6953 12860 6987
rect 12808 6944 12860 6953
rect 13360 6987 13412 6996
rect 13360 6953 13369 6987
rect 13369 6953 13403 6987
rect 13403 6953 13412 6987
rect 13360 6944 13412 6953
rect 17960 6944 18012 6996
rect 18788 6987 18840 6996
rect 18788 6953 18797 6987
rect 18797 6953 18831 6987
rect 18831 6953 18840 6987
rect 18788 6944 18840 6953
rect 19340 6987 19392 6996
rect 19340 6953 19349 6987
rect 19349 6953 19383 6987
rect 19383 6953 19392 6987
rect 19340 6944 19392 6953
rect 8208 6919 8260 6928
rect 8208 6885 8217 6919
rect 8217 6885 8251 6919
rect 8251 6885 8260 6919
rect 8208 6876 8260 6885
rect 11428 6876 11480 6928
rect 14096 6876 14148 6928
rect 16396 6919 16448 6928
rect 16396 6885 16405 6919
rect 16405 6885 16439 6919
rect 16439 6885 16448 6919
rect 16396 6876 16448 6885
rect 21272 6876 21324 6928
rect 9956 6851 10008 6860
rect 9956 6817 9965 6851
rect 9965 6817 9999 6851
rect 9999 6817 10008 6851
rect 9956 6808 10008 6817
rect 11244 6851 11296 6860
rect 11244 6817 11253 6851
rect 11253 6817 11287 6851
rect 11287 6817 11296 6851
rect 11244 6808 11296 6817
rect 4620 6672 4672 6724
rect 8852 6740 8904 6792
rect 9128 6740 9180 6792
rect 12164 6808 12216 6860
rect 12716 6808 12768 6860
rect 13636 6851 13688 6860
rect 13636 6817 13645 6851
rect 13645 6817 13679 6851
rect 13679 6817 13688 6851
rect 13636 6808 13688 6817
rect 18328 6808 18380 6860
rect 11612 6783 11664 6792
rect 11612 6749 11621 6783
rect 11621 6749 11655 6783
rect 11655 6749 11664 6783
rect 11612 6740 11664 6749
rect 16304 6783 16356 6792
rect 16304 6749 16313 6783
rect 16313 6749 16347 6783
rect 16347 6749 16356 6783
rect 16304 6740 16356 6749
rect 21456 6740 21508 6792
rect 8484 6672 8536 6724
rect 11060 6672 11112 6724
rect 11888 6672 11940 6724
rect 16856 6715 16908 6724
rect 16856 6681 16865 6715
rect 16865 6681 16899 6715
rect 16899 6681 16908 6715
rect 16856 6672 16908 6681
rect 4804 6604 4856 6656
rect 6184 6604 6236 6656
rect 8760 6604 8812 6656
rect 10876 6604 10928 6656
rect 12440 6647 12492 6656
rect 12440 6613 12449 6647
rect 12449 6613 12483 6647
rect 12483 6613 12492 6647
rect 12440 6604 12492 6613
rect 15016 6604 15068 6656
rect 21364 6604 21416 6656
rect 4982 6502 5034 6554
rect 5046 6502 5098 6554
rect 5110 6502 5162 6554
rect 5174 6502 5226 6554
rect 12982 6502 13034 6554
rect 13046 6502 13098 6554
rect 13110 6502 13162 6554
rect 13174 6502 13226 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 2412 6264 2464 6316
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 1952 6196 2004 6248
rect 3700 6400 3752 6452
rect 4712 6400 4764 6452
rect 6184 6443 6236 6452
rect 6184 6409 6193 6443
rect 6193 6409 6227 6443
rect 6227 6409 6236 6443
rect 6184 6400 6236 6409
rect 8208 6400 8260 6452
rect 8576 6400 8628 6452
rect 9956 6443 10008 6452
rect 9956 6409 9965 6443
rect 9965 6409 9999 6443
rect 9999 6409 10008 6443
rect 9956 6400 10008 6409
rect 4344 6332 4396 6384
rect 8116 6332 8168 6384
rect 10968 6400 11020 6452
rect 11888 6443 11940 6452
rect 11888 6409 11897 6443
rect 11897 6409 11931 6443
rect 11931 6409 11940 6443
rect 11888 6400 11940 6409
rect 12716 6443 12768 6452
rect 12716 6409 12725 6443
rect 12725 6409 12759 6443
rect 12759 6409 12768 6443
rect 12716 6400 12768 6409
rect 14832 6443 14884 6452
rect 14832 6409 14841 6443
rect 14841 6409 14875 6443
rect 14875 6409 14884 6443
rect 14832 6400 14884 6409
rect 15844 6443 15896 6452
rect 15844 6409 15853 6443
rect 15853 6409 15887 6443
rect 15887 6409 15896 6443
rect 15844 6400 15896 6409
rect 16396 6400 16448 6452
rect 18328 6400 18380 6452
rect 20352 6443 20404 6452
rect 20352 6409 20361 6443
rect 20361 6409 20395 6443
rect 20395 6409 20404 6443
rect 20352 6400 20404 6409
rect 21272 6400 21324 6452
rect 21364 6332 21416 6384
rect 3792 6196 3844 6248
rect 204 6128 256 6180
rect 112 6060 164 6112
rect 3608 6060 3660 6112
rect 7472 6264 7524 6316
rect 8852 6264 8904 6316
rect 14740 6264 14792 6316
rect 16304 6264 16356 6316
rect 18788 6264 18840 6316
rect 21456 6264 21508 6316
rect 4252 6239 4304 6248
rect 4252 6205 4261 6239
rect 4261 6205 4295 6239
rect 4295 6205 4304 6239
rect 4252 6196 4304 6205
rect 4804 6196 4856 6248
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 7288 6196 7340 6248
rect 7564 6196 7616 6248
rect 7932 6196 7984 6248
rect 10968 6239 11020 6248
rect 10968 6205 10977 6239
rect 10977 6205 11011 6239
rect 11011 6205 11020 6239
rect 10968 6196 11020 6205
rect 13360 6196 13412 6248
rect 5356 6171 5408 6180
rect 5356 6137 5365 6171
rect 5365 6137 5399 6171
rect 5399 6137 5408 6171
rect 5356 6128 5408 6137
rect 6368 6128 6420 6180
rect 8668 6128 8720 6180
rect 8760 6128 8812 6180
rect 9128 6171 9180 6180
rect 9128 6137 9137 6171
rect 9137 6137 9171 6171
rect 9171 6137 9180 6171
rect 10508 6171 10560 6180
rect 9128 6128 9180 6137
rect 10508 6137 10517 6171
rect 10517 6137 10551 6171
rect 10551 6137 10560 6171
rect 10508 6128 10560 6137
rect 12716 6128 12768 6180
rect 14832 6128 14884 6180
rect 7564 6060 7616 6112
rect 7840 6103 7892 6112
rect 7840 6069 7849 6103
rect 7849 6069 7883 6103
rect 7883 6069 7892 6103
rect 7840 6060 7892 6069
rect 13268 6103 13320 6112
rect 13268 6069 13277 6103
rect 13277 6069 13311 6103
rect 13311 6069 13320 6103
rect 13268 6060 13320 6069
rect 16672 6060 16724 6112
rect 20628 6171 20680 6180
rect 20628 6137 20637 6171
rect 20637 6137 20671 6171
rect 20671 6137 20680 6171
rect 20628 6128 20680 6137
rect 18052 6060 18104 6112
rect 20352 6060 20404 6112
rect 8982 5958 9034 6010
rect 9046 5958 9098 6010
rect 9110 5958 9162 6010
rect 9174 5958 9226 6010
rect 16982 5958 17034 6010
rect 17046 5958 17098 6010
rect 17110 5958 17162 6010
rect 17174 5958 17226 6010
rect 2044 5856 2096 5908
rect 8024 5899 8076 5908
rect 8024 5865 8033 5899
rect 8033 5865 8067 5899
rect 8067 5865 8076 5899
rect 8024 5856 8076 5865
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 8668 5856 8720 5908
rect 11244 5856 11296 5908
rect 13360 5899 13412 5908
rect 13360 5865 13369 5899
rect 13369 5865 13403 5899
rect 13403 5865 13412 5899
rect 13360 5856 13412 5865
rect 13636 5899 13688 5908
rect 13636 5865 13645 5899
rect 13645 5865 13679 5899
rect 13679 5865 13688 5899
rect 13636 5856 13688 5865
rect 14740 5856 14792 5908
rect 18788 5856 18840 5908
rect 20168 5899 20220 5908
rect 20168 5865 20177 5899
rect 20177 5865 20211 5899
rect 20211 5865 20220 5899
rect 20168 5856 20220 5865
rect 20444 5856 20496 5908
rect 20628 5899 20680 5908
rect 20628 5865 20637 5899
rect 20637 5865 20671 5899
rect 20671 5865 20680 5899
rect 20628 5856 20680 5865
rect 4252 5788 4304 5840
rect 12624 5788 12676 5840
rect 16580 5831 16632 5840
rect 16580 5797 16589 5831
rect 16589 5797 16623 5831
rect 16623 5797 16632 5831
rect 16580 5788 16632 5797
rect 2964 5720 3016 5772
rect 4344 5763 4396 5772
rect 4344 5729 4353 5763
rect 4353 5729 4387 5763
rect 4387 5729 4396 5763
rect 4344 5720 4396 5729
rect 4620 5763 4672 5772
rect 4620 5729 4629 5763
rect 4629 5729 4663 5763
rect 4663 5729 4672 5763
rect 4620 5720 4672 5729
rect 6000 5763 6052 5772
rect 6000 5729 6009 5763
rect 6009 5729 6043 5763
rect 6043 5729 6052 5763
rect 6000 5720 6052 5729
rect 6276 5763 6328 5772
rect 6276 5729 6285 5763
rect 6285 5729 6319 5763
rect 6319 5729 6328 5763
rect 6276 5720 6328 5729
rect 7840 5720 7892 5772
rect 10876 5763 10928 5772
rect 10876 5729 10885 5763
rect 10885 5729 10919 5763
rect 10919 5729 10928 5763
rect 10876 5720 10928 5729
rect 11428 5763 11480 5772
rect 11428 5729 11437 5763
rect 11437 5729 11471 5763
rect 11471 5729 11480 5763
rect 11428 5720 11480 5729
rect 21272 5788 21324 5840
rect 21732 5788 21784 5840
rect 1768 5695 1820 5704
rect 1768 5661 1777 5695
rect 1777 5661 1811 5695
rect 1811 5661 1820 5695
rect 1768 5652 1820 5661
rect 5356 5652 5408 5704
rect 5816 5652 5868 5704
rect 12440 5695 12492 5704
rect 12440 5661 12449 5695
rect 12449 5661 12483 5695
rect 12483 5661 12492 5695
rect 12440 5652 12492 5661
rect 16672 5652 16724 5704
rect 16856 5695 16908 5704
rect 16856 5661 16865 5695
rect 16865 5661 16899 5695
rect 16899 5661 16908 5695
rect 16856 5652 16908 5661
rect 6644 5516 6696 5568
rect 9404 5516 9456 5568
rect 4982 5414 5034 5466
rect 5046 5414 5098 5466
rect 5110 5414 5162 5466
rect 5174 5414 5226 5466
rect 12982 5414 13034 5466
rect 13046 5414 13098 5466
rect 13110 5414 13162 5466
rect 13174 5414 13226 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 2964 5355 3016 5364
rect 2964 5321 2973 5355
rect 2973 5321 3007 5355
rect 3007 5321 3016 5355
rect 2964 5312 3016 5321
rect 3792 5355 3844 5364
rect 3792 5321 3801 5355
rect 3801 5321 3835 5355
rect 3835 5321 3844 5355
rect 3792 5312 3844 5321
rect 6184 5312 6236 5364
rect 7288 5355 7340 5364
rect 20 5244 72 5296
rect 7288 5321 7297 5355
rect 7297 5321 7331 5355
rect 7331 5321 7340 5355
rect 7288 5312 7340 5321
rect 8024 5312 8076 5364
rect 8668 5312 8720 5364
rect 9404 5312 9456 5364
rect 12164 5355 12216 5364
rect 12164 5321 12173 5355
rect 12173 5321 12207 5355
rect 12207 5321 12216 5355
rect 12164 5312 12216 5321
rect 13360 5312 13412 5364
rect 15844 5355 15896 5364
rect 15844 5321 15853 5355
rect 15853 5321 15887 5355
rect 15887 5321 15896 5355
rect 15844 5312 15896 5321
rect 21272 5312 21324 5364
rect 10600 5287 10652 5296
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 4344 5176 4396 5228
rect 3792 5108 3844 5160
rect 4620 5108 4672 5160
rect 10600 5253 10609 5287
rect 10609 5253 10643 5287
rect 10643 5253 10652 5287
rect 10600 5244 10652 5253
rect 11796 5244 11848 5296
rect 6828 5176 6880 5228
rect 8116 5176 8168 5228
rect 8484 5176 8536 5228
rect 10508 5176 10560 5228
rect 10968 5176 11020 5228
rect 16856 5244 16908 5296
rect 13820 5219 13872 5228
rect 13820 5185 13829 5219
rect 13829 5185 13863 5219
rect 13863 5185 13872 5219
rect 13820 5176 13872 5185
rect 16580 5176 16632 5228
rect 20168 5219 20220 5228
rect 20168 5185 20177 5219
rect 20177 5185 20211 5219
rect 20211 5185 20220 5219
rect 20168 5176 20220 5185
rect 20444 5219 20496 5228
rect 20444 5185 20453 5219
rect 20453 5185 20487 5219
rect 20487 5185 20496 5219
rect 20444 5176 20496 5185
rect 4160 5040 4212 5092
rect 4804 5040 4856 5092
rect 6276 5108 6328 5160
rect 7748 5108 7800 5160
rect 15844 5108 15896 5160
rect 18144 5108 18196 5160
rect 6000 5040 6052 5092
rect 8116 5040 8168 5092
rect 11520 5083 11572 5092
rect 11520 5049 11529 5083
rect 11529 5049 11563 5083
rect 11563 5049 11572 5083
rect 11520 5040 11572 5049
rect 13452 5040 13504 5092
rect 18788 5040 18840 5092
rect 2412 5015 2464 5024
rect 2412 4981 2421 5015
rect 2421 4981 2455 5015
rect 2455 4981 2464 5015
rect 2412 4972 2464 4981
rect 3976 5015 4028 5024
rect 3976 4981 3985 5015
rect 3985 4981 4019 5015
rect 4019 4981 4028 5015
rect 3976 4972 4028 4981
rect 4988 5015 5040 5024
rect 4988 4981 4997 5015
rect 4997 4981 5031 5015
rect 5031 4981 5040 5015
rect 4988 4972 5040 4981
rect 5356 4972 5408 5024
rect 9496 4972 9548 5024
rect 9772 4972 9824 5024
rect 10876 4972 10928 5024
rect 12624 5015 12676 5024
rect 12624 4981 12633 5015
rect 12633 4981 12667 5015
rect 12667 4981 12676 5015
rect 12624 4972 12676 4981
rect 19892 5015 19944 5024
rect 19892 4981 19901 5015
rect 19901 4981 19935 5015
rect 19935 4981 19944 5015
rect 19892 4972 19944 4981
rect 8982 4870 9034 4922
rect 9046 4870 9098 4922
rect 9110 4870 9162 4922
rect 9174 4870 9226 4922
rect 16982 4870 17034 4922
rect 17046 4870 17098 4922
rect 17110 4870 17162 4922
rect 17174 4870 17226 4922
rect 2504 4768 2556 4820
rect 3056 4768 3108 4820
rect 2964 4700 3016 4752
rect 4620 4768 4672 4820
rect 4988 4768 5040 4820
rect 6000 4768 6052 4820
rect 7840 4768 7892 4820
rect 8484 4768 8536 4820
rect 10968 4768 11020 4820
rect 11520 4768 11572 4820
rect 15476 4768 15528 4820
rect 16672 4768 16724 4820
rect 4252 4700 4304 4752
rect 6828 4743 6880 4752
rect 6828 4709 6837 4743
rect 6837 4709 6871 4743
rect 6871 4709 6880 4743
rect 6828 4700 6880 4709
rect 11428 4700 11480 4752
rect 12440 4743 12492 4752
rect 12440 4709 12449 4743
rect 12449 4709 12483 4743
rect 12483 4709 12492 4743
rect 12440 4700 12492 4709
rect 13268 4743 13320 4752
rect 13268 4709 13277 4743
rect 13277 4709 13311 4743
rect 13311 4709 13320 4743
rect 13268 4700 13320 4709
rect 13820 4743 13872 4752
rect 13820 4709 13829 4743
rect 13829 4709 13863 4743
rect 13863 4709 13872 4743
rect 18144 4743 18196 4752
rect 13820 4700 13872 4709
rect 18144 4709 18153 4743
rect 18153 4709 18187 4743
rect 18187 4709 18196 4743
rect 18144 4700 18196 4709
rect 20812 4700 20864 4752
rect 5816 4632 5868 4684
rect 7656 4632 7708 4684
rect 9680 4675 9732 4684
rect 9680 4641 9689 4675
rect 9689 4641 9723 4675
rect 9723 4641 9732 4675
rect 9680 4632 9732 4641
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 2504 4564 2556 4616
rect 3976 4564 4028 4616
rect 9496 4564 9548 4616
rect 11336 4632 11388 4684
rect 17500 4675 17552 4684
rect 17500 4641 17509 4675
rect 17509 4641 17543 4675
rect 17543 4641 17552 4675
rect 17500 4632 17552 4641
rect 17868 4675 17920 4684
rect 17868 4641 17877 4675
rect 17877 4641 17911 4675
rect 17911 4641 17920 4675
rect 17868 4632 17920 4641
rect 20076 4632 20128 4684
rect 11244 4607 11296 4616
rect 11244 4573 11253 4607
rect 11253 4573 11287 4607
rect 11287 4573 11296 4607
rect 11244 4564 11296 4573
rect 12808 4564 12860 4616
rect 15292 4607 15344 4616
rect 15292 4573 15301 4607
rect 15301 4573 15335 4607
rect 15335 4573 15344 4607
rect 15292 4564 15344 4573
rect 21272 4564 21324 4616
rect 10140 4496 10192 4548
rect 20444 4496 20496 4548
rect 1860 4471 1912 4480
rect 1860 4437 1869 4471
rect 1869 4437 1903 4471
rect 1903 4437 1912 4471
rect 1860 4428 1912 4437
rect 3792 4428 3844 4480
rect 14464 4428 14516 4480
rect 16212 4471 16264 4480
rect 16212 4437 16221 4471
rect 16221 4437 16255 4471
rect 16255 4437 16264 4471
rect 16212 4428 16264 4437
rect 4982 4326 5034 4378
rect 5046 4326 5098 4378
rect 5110 4326 5162 4378
rect 5174 4326 5226 4378
rect 12982 4326 13034 4378
rect 13046 4326 13098 4378
rect 13110 4326 13162 4378
rect 13174 4326 13226 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 1768 4224 1820 4276
rect 2320 4224 2372 4276
rect 2964 4156 3016 4208
rect 4252 4224 4304 4276
rect 8024 4224 8076 4276
rect 9680 4267 9732 4276
rect 9680 4233 9689 4267
rect 9689 4233 9723 4267
rect 9723 4233 9732 4267
rect 9680 4224 9732 4233
rect 11336 4267 11388 4276
rect 11336 4233 11345 4267
rect 11345 4233 11379 4267
rect 11379 4233 11388 4267
rect 11336 4224 11388 4233
rect 12808 4267 12860 4276
rect 12808 4233 12817 4267
rect 12817 4233 12851 4267
rect 12851 4233 12860 4267
rect 12808 4224 12860 4233
rect 4804 4156 4856 4208
rect 7932 4156 7984 4208
rect 2504 4131 2556 4140
rect 2504 4097 2513 4131
rect 2513 4097 2547 4131
rect 2547 4097 2556 4131
rect 2504 4088 2556 4097
rect 5356 4088 5408 4140
rect 5908 4020 5960 4072
rect 15292 4224 15344 4276
rect 20076 4224 20128 4276
rect 21272 4267 21324 4276
rect 21272 4233 21281 4267
rect 21281 4233 21315 4267
rect 21315 4233 21324 4267
rect 21272 4224 21324 4233
rect 13268 4156 13320 4208
rect 9496 4020 9548 4072
rect 10140 4063 10192 4072
rect 10140 4029 10149 4063
rect 10149 4029 10183 4063
rect 10183 4029 10192 4063
rect 10140 4020 10192 4029
rect 12532 4020 12584 4072
rect 14464 4063 14516 4072
rect 14464 4029 14473 4063
rect 14473 4029 14507 4063
rect 14507 4029 14516 4063
rect 17868 4156 17920 4208
rect 16488 4131 16540 4140
rect 16488 4097 16497 4131
rect 16497 4097 16531 4131
rect 16531 4097 16540 4131
rect 16488 4088 16540 4097
rect 19892 4063 19944 4072
rect 14464 4020 14516 4029
rect 19892 4029 19901 4063
rect 19901 4029 19935 4063
rect 19935 4029 19944 4063
rect 19892 4020 19944 4029
rect 1860 3995 1912 4004
rect 1860 3961 1869 3995
rect 1869 3961 1903 3995
rect 1903 3961 1912 3995
rect 1860 3952 1912 3961
rect 3792 3995 3844 4004
rect 3792 3961 3801 3995
rect 3801 3961 3835 3995
rect 3835 3961 3844 3995
rect 3792 3952 3844 3961
rect 9312 3995 9364 4004
rect 9312 3961 9321 3995
rect 9321 3961 9355 3995
rect 9355 3961 9364 3995
rect 9312 3952 9364 3961
rect 10048 3995 10100 4004
rect 10048 3961 10057 3995
rect 10057 3961 10091 3995
rect 10091 3961 10100 3995
rect 10048 3952 10100 3961
rect 12624 3952 12676 4004
rect 15476 3952 15528 4004
rect 16120 3995 16172 4004
rect 16120 3961 16129 3995
rect 16129 3961 16163 3995
rect 16163 3961 16172 3995
rect 16120 3952 16172 3961
rect 16212 3995 16264 4004
rect 16212 3961 16221 3995
rect 16221 3961 16255 3995
rect 16255 3961 16264 3995
rect 16212 3952 16264 3961
rect 20812 3952 20864 4004
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 8300 3884 8352 3936
rect 11612 3884 11664 3936
rect 17500 3927 17552 3936
rect 17500 3893 17509 3927
rect 17509 3893 17543 3927
rect 17543 3893 17552 3927
rect 17500 3884 17552 3893
rect 8982 3782 9034 3834
rect 9046 3782 9098 3834
rect 9110 3782 9162 3834
rect 9174 3782 9226 3834
rect 16982 3782 17034 3834
rect 17046 3782 17098 3834
rect 17110 3782 17162 3834
rect 17174 3782 17226 3834
rect 112 3680 164 3732
rect 2320 3723 2372 3732
rect 2320 3689 2329 3723
rect 2329 3689 2363 3723
rect 2363 3689 2372 3723
rect 2320 3680 2372 3689
rect 3976 3680 4028 3732
rect 8392 3723 8444 3732
rect 8392 3689 8401 3723
rect 8401 3689 8435 3723
rect 8435 3689 8444 3723
rect 8392 3680 8444 3689
rect 9312 3680 9364 3732
rect 10048 3723 10100 3732
rect 1860 3612 1912 3664
rect 4620 3655 4672 3664
rect 4620 3621 4629 3655
rect 4629 3621 4663 3655
rect 4663 3621 4672 3655
rect 4620 3612 4672 3621
rect 2320 3544 2372 3596
rect 6920 3544 6972 3596
rect 8484 3544 8536 3596
rect 10048 3689 10057 3723
rect 10057 3689 10091 3723
rect 10091 3689 10100 3723
rect 10048 3680 10100 3689
rect 10140 3680 10192 3732
rect 11244 3680 11296 3732
rect 12532 3680 12584 3732
rect 16212 3680 16264 3732
rect 19892 3723 19944 3732
rect 19892 3689 19901 3723
rect 19901 3689 19935 3723
rect 19935 3689 19944 3723
rect 19892 3680 19944 3689
rect 11612 3655 11664 3664
rect 11612 3621 11621 3655
rect 11621 3621 11655 3655
rect 11655 3621 11664 3655
rect 11612 3612 11664 3621
rect 11704 3612 11756 3664
rect 15936 3655 15988 3664
rect 15936 3621 15945 3655
rect 15945 3621 15979 3655
rect 15979 3621 15988 3655
rect 15936 3612 15988 3621
rect 16120 3612 16172 3664
rect 20444 3612 20496 3664
rect 13452 3544 13504 3596
rect 13820 3544 13872 3596
rect 16488 3587 16540 3596
rect 16488 3553 16497 3587
rect 16497 3553 16531 3587
rect 16531 3553 16540 3587
rect 16488 3544 16540 3553
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 4804 3519 4856 3528
rect 4804 3485 4813 3519
rect 4813 3485 4847 3519
rect 4847 3485 4856 3519
rect 4804 3476 4856 3485
rect 10968 3476 11020 3528
rect 12808 3476 12860 3528
rect 15476 3476 15528 3528
rect 6828 3383 6880 3392
rect 6828 3349 6837 3383
rect 6837 3349 6871 3383
rect 6871 3349 6880 3383
rect 6828 3340 6880 3349
rect 9864 3340 9916 3392
rect 10416 3340 10468 3392
rect 11796 3340 11848 3392
rect 13360 3340 13412 3392
rect 4982 3238 5034 3290
rect 5046 3238 5098 3290
rect 5110 3238 5162 3290
rect 5174 3238 5226 3290
rect 12982 3238 13034 3290
rect 13046 3238 13098 3290
rect 13110 3238 13162 3290
rect 13174 3238 13226 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 1400 3136 1452 3188
rect 3792 3136 3844 3188
rect 10048 3179 10100 3188
rect 112 3000 164 3052
rect 2320 3043 2372 3052
rect 2320 3009 2329 3043
rect 2329 3009 2363 3043
rect 2363 3009 2372 3043
rect 2320 3000 2372 3009
rect 2504 2975 2556 2984
rect 2504 2941 2522 2975
rect 2522 2941 2556 2975
rect 2504 2932 2556 2941
rect 10048 3145 10057 3179
rect 10057 3145 10091 3179
rect 10091 3145 10100 3179
rect 10048 3136 10100 3145
rect 10416 3179 10468 3188
rect 10416 3145 10425 3179
rect 10425 3145 10459 3179
rect 10459 3145 10468 3179
rect 10416 3136 10468 3145
rect 13452 3179 13504 3188
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 13820 3136 13872 3188
rect 15476 3179 15528 3188
rect 15476 3145 15485 3179
rect 15485 3145 15519 3179
rect 15519 3145 15528 3179
rect 15476 3136 15528 3145
rect 4620 3000 4672 3052
rect 11152 3068 11204 3120
rect 8116 3000 8168 3052
rect 10232 3000 10284 3052
rect 10692 3000 10744 3052
rect 10968 3043 11020 3052
rect 10968 3009 10977 3043
rect 10977 3009 11011 3043
rect 11011 3009 11020 3043
rect 10968 3000 11020 3009
rect 12532 3043 12584 3052
rect 12532 3009 12541 3043
rect 12541 3009 12575 3043
rect 12575 3009 12584 3043
rect 12532 3000 12584 3009
rect 12808 3043 12860 3052
rect 12808 3009 12817 3043
rect 12817 3009 12851 3043
rect 12851 3009 12860 3043
rect 12808 3000 12860 3009
rect 6000 2864 6052 2916
rect 6828 2907 6880 2916
rect 6828 2873 6837 2907
rect 6837 2873 6871 2907
rect 6871 2873 6880 2907
rect 6828 2864 6880 2873
rect 16488 3068 16540 3120
rect 15936 3000 15988 3052
rect 16212 2975 16264 2984
rect 16212 2941 16221 2975
rect 16221 2941 16255 2975
rect 16255 2941 16264 2975
rect 16212 2932 16264 2941
rect 10416 2864 10468 2916
rect 12624 2907 12676 2916
rect 12624 2873 12633 2907
rect 12633 2873 12667 2907
rect 12667 2873 12676 2907
rect 12624 2864 12676 2873
rect 16580 2864 16632 2916
rect 6920 2796 6972 2848
rect 7748 2839 7800 2848
rect 7748 2805 7757 2839
rect 7757 2805 7791 2839
rect 7791 2805 7800 2839
rect 7748 2796 7800 2805
rect 8484 2796 8536 2848
rect 9404 2839 9456 2848
rect 9404 2805 9413 2839
rect 9413 2805 9447 2839
rect 9447 2805 9456 2839
rect 9404 2796 9456 2805
rect 11612 2839 11664 2848
rect 11612 2805 11621 2839
rect 11621 2805 11655 2839
rect 11655 2805 11664 2839
rect 11612 2796 11664 2805
rect 16028 2796 16080 2848
rect 19524 2796 19576 2848
rect 8982 2694 9034 2746
rect 9046 2694 9098 2746
rect 9110 2694 9162 2746
rect 9174 2694 9226 2746
rect 16982 2694 17034 2746
rect 17046 2694 17098 2746
rect 17110 2694 17162 2746
rect 17174 2694 17226 2746
rect 2228 2592 2280 2644
rect 9404 2592 9456 2644
rect 6000 2567 6052 2576
rect 6000 2533 6009 2567
rect 6009 2533 6043 2567
rect 6043 2533 6052 2567
rect 6000 2524 6052 2533
rect 9864 2567 9916 2576
rect 9864 2533 9873 2567
rect 9873 2533 9907 2567
rect 9907 2533 9916 2567
rect 9864 2524 9916 2533
rect 10692 2592 10744 2644
rect 21456 2592 21508 2644
rect 10968 2524 11020 2576
rect 12624 2567 12676 2576
rect 12624 2533 12633 2567
rect 12633 2533 12667 2567
rect 12667 2533 12676 2567
rect 12624 2524 12676 2533
rect 1860 2499 1912 2508
rect 1860 2465 1869 2499
rect 1869 2465 1903 2499
rect 1903 2465 1912 2499
rect 1860 2456 1912 2465
rect 4528 2499 4580 2508
rect 4528 2465 4537 2499
rect 4537 2465 4571 2499
rect 4571 2465 4580 2499
rect 4528 2456 4580 2465
rect 1032 2320 1084 2372
rect 7196 2456 7248 2508
rect 8300 2456 8352 2508
rect 7748 2388 7800 2440
rect 9864 2388 9916 2440
rect 11612 2456 11664 2508
rect 12808 2456 12860 2508
rect 15568 2456 15620 2508
rect 16580 2499 16632 2508
rect 16580 2465 16589 2499
rect 16589 2465 16623 2499
rect 16623 2465 16632 2499
rect 16580 2456 16632 2465
rect 9956 2320 10008 2372
rect 13268 2320 13320 2372
rect 15384 2252 15436 2304
rect 16856 2252 16908 2304
rect 17224 2252 17276 2304
rect 21272 2252 21324 2304
rect 22836 2252 22888 2304
rect 4982 2150 5034 2202
rect 5046 2150 5098 2202
rect 5110 2150 5162 2202
rect 5174 2150 5226 2202
rect 12982 2150 13034 2202
rect 13046 2150 13098 2202
rect 13110 2150 13162 2202
rect 13174 2150 13226 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
<< metal2 >>
rect 1214 23610 1270 24000
rect 3606 23610 3662 24000
rect 1214 23582 1624 23610
rect 1214 23520 1270 23582
rect 1214 21584 1270 21593
rect 1214 21519 1270 21528
rect 1228 19990 1256 21519
rect 1596 20602 1624 23582
rect 3436 23582 3662 23610
rect 3436 20602 3464 23582
rect 3606 23520 3662 23582
rect 5998 23610 6054 24000
rect 8390 23610 8446 24000
rect 10782 23610 10838 24000
rect 13174 23610 13230 24000
rect 5998 23582 6224 23610
rect 5998 23520 6054 23582
rect 5814 22808 5870 22817
rect 5814 22743 5870 22752
rect 4956 21788 5252 21808
rect 5012 21786 5036 21788
rect 5092 21786 5116 21788
rect 5172 21786 5196 21788
rect 5034 21734 5036 21786
rect 5098 21734 5110 21786
rect 5172 21734 5174 21786
rect 5012 21732 5036 21734
rect 5092 21732 5116 21734
rect 5172 21732 5196 21734
rect 4956 21712 5252 21732
rect 4956 20700 5252 20720
rect 5012 20698 5036 20700
rect 5092 20698 5116 20700
rect 5172 20698 5196 20700
rect 5034 20646 5036 20698
rect 5098 20646 5110 20698
rect 5172 20646 5174 20698
rect 5012 20644 5036 20646
rect 5092 20644 5116 20646
rect 5172 20644 5196 20646
rect 4956 20624 5252 20644
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 5828 20398 5856 22743
rect 5816 20392 5868 20398
rect 1306 20360 1362 20369
rect 5816 20334 5868 20340
rect 1306 20295 1362 20304
rect 1216 19984 1268 19990
rect 1216 19926 1268 19932
rect 1228 19514 1256 19926
rect 1216 19508 1268 19514
rect 1216 19450 1268 19456
rect 1214 19136 1270 19145
rect 1214 19071 1270 19080
rect 1228 18222 1256 19071
rect 1320 18834 1348 20295
rect 2044 20256 2096 20262
rect 2044 20198 2096 20204
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 1308 18828 1360 18834
rect 1308 18770 1360 18776
rect 1320 18426 1348 18770
rect 1308 18420 1360 18426
rect 1308 18362 1360 18368
rect 1216 18216 1268 18222
rect 1216 18158 1268 18164
rect 1490 18048 1546 18057
rect 1490 17983 1546 17992
rect 112 17740 164 17746
rect 112 17682 164 17688
rect 124 17377 152 17682
rect 110 17368 166 17377
rect 110 17303 166 17312
rect 1504 17134 1532 17983
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1467 17128 1532 17134
rect 1519 17088 1532 17128
rect 1467 17070 1519 17076
rect 1582 16416 1638 16425
rect 1582 16351 1638 16360
rect 1596 16250 1624 16351
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1412 15706 1440 15982
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1596 14618 1624 15438
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1688 12850 1716 17478
rect 1872 17338 1900 17682
rect 1860 17332 1912 17338
rect 1860 17274 1912 17280
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1780 13938 1808 16390
rect 1872 14550 1900 16934
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1964 15910 1992 16594
rect 1952 15904 2004 15910
rect 1952 15846 2004 15852
rect 1964 15473 1992 15846
rect 1950 15464 2006 15473
rect 1950 15399 2006 15408
rect 2056 15065 2084 20198
rect 3896 20058 3924 20198
rect 3884 20052 3936 20058
rect 3884 19994 3936 20000
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 2516 17202 2544 18022
rect 2884 17882 2912 19654
rect 4956 19612 5252 19632
rect 5012 19610 5036 19612
rect 5092 19610 5116 19612
rect 5172 19610 5196 19612
rect 5034 19558 5036 19610
rect 5098 19558 5110 19610
rect 5172 19558 5174 19610
rect 5012 19556 5036 19558
rect 5092 19556 5116 19558
rect 5172 19556 5196 19558
rect 4956 19536 5252 19556
rect 4956 18524 5252 18544
rect 5012 18522 5036 18524
rect 5092 18522 5116 18524
rect 5172 18522 5196 18524
rect 5034 18470 5036 18522
rect 5098 18470 5110 18522
rect 5172 18470 5174 18522
rect 5012 18468 5036 18470
rect 5092 18468 5116 18470
rect 5172 18468 5196 18470
rect 4956 18448 5252 18468
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2780 17740 2832 17746
rect 2780 17682 2832 17688
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 2516 16794 2544 17138
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2700 16726 2728 17478
rect 2792 17066 2820 17682
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5356 17536 5408 17542
rect 5356 17478 5408 17484
rect 4956 17436 5252 17456
rect 5012 17434 5036 17436
rect 5092 17434 5116 17436
rect 5172 17434 5196 17436
rect 5034 17382 5036 17434
rect 5098 17382 5110 17434
rect 5172 17382 5174 17434
rect 5012 17380 5036 17382
rect 5092 17380 5116 17382
rect 5172 17380 5196 17382
rect 4956 17360 5252 17380
rect 3148 17196 3200 17202
rect 3148 17138 3200 17144
rect 2780 17060 2832 17066
rect 2780 17002 2832 17008
rect 3160 16726 3188 17138
rect 5368 17066 5396 17478
rect 5644 17066 5672 17614
rect 3792 17060 3844 17066
rect 3792 17002 3844 17008
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 5632 17060 5684 17066
rect 5632 17002 5684 17008
rect 2688 16720 2740 16726
rect 2688 16662 2740 16668
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2240 15910 2268 16526
rect 2700 16250 2728 16662
rect 3804 16250 3832 17002
rect 5368 16658 5396 17002
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 4956 16348 5252 16368
rect 5012 16346 5036 16348
rect 5092 16346 5116 16348
rect 5172 16346 5196 16348
rect 5034 16294 5036 16346
rect 5098 16294 5110 16346
rect 5172 16294 5174 16346
rect 5012 16292 5036 16294
rect 5092 16292 5116 16294
rect 5172 16292 5196 16294
rect 4956 16272 5252 16292
rect 5368 16250 5396 16594
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 2228 15904 2280 15910
rect 2228 15846 2280 15852
rect 2042 15056 2098 15065
rect 2042 14991 2098 15000
rect 2136 14952 2188 14958
rect 2136 14894 2188 14900
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 2056 14550 2084 14758
rect 1860 14544 1912 14550
rect 1860 14486 1912 14492
rect 2044 14544 2096 14550
rect 2044 14486 2096 14492
rect 1872 14006 1900 14486
rect 2056 14074 2084 14486
rect 2148 14074 2176 14894
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 1860 14000 1912 14006
rect 1860 13942 1912 13948
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1780 13530 1808 13874
rect 2148 13802 2176 14010
rect 2136 13796 2188 13802
rect 2136 13738 2188 13744
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1780 12918 1808 13330
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1768 12912 1820 12918
rect 1768 12854 1820 12860
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1780 12374 1808 12854
rect 1872 12714 1900 13126
rect 1860 12708 1912 12714
rect 1860 12650 1912 12656
rect 2044 12708 2096 12714
rect 2044 12650 2096 12656
rect 1768 12368 1820 12374
rect 1768 12310 1820 12316
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1122 12064 1178 12073
rect 1122 11999 1178 12008
rect 1136 11762 1164 11999
rect 1124 11756 1176 11762
rect 1124 11698 1176 11704
rect 1688 11558 1716 12174
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1688 11354 1716 11494
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1780 11082 1808 12310
rect 2056 12238 2084 12650
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 1860 11280 1912 11286
rect 1860 11222 1912 11228
rect 1768 11076 1820 11082
rect 1768 11018 1820 11024
rect 1872 10674 1900 11222
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 18 10160 74 10169
rect 18 10095 74 10104
rect 32 5302 60 10095
rect 1964 9994 1992 11086
rect 2056 10538 2084 12174
rect 2044 10532 2096 10538
rect 2044 10474 2096 10480
rect 2056 10266 2084 10474
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 1952 9988 2004 9994
rect 1952 9930 2004 9936
rect 2056 9382 2084 10066
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2148 9722 2176 9998
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2148 9382 2176 9658
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 112 9172 164 9178
rect 112 9114 164 9120
rect 124 8945 152 9114
rect 2056 9110 2084 9318
rect 2044 9104 2096 9110
rect 2044 9046 2096 9052
rect 110 8936 166 8945
rect 110 8871 166 8880
rect 1400 8832 1452 8838
rect 1400 8774 1452 8780
rect 1412 8430 1440 8774
rect 2056 8566 2084 9046
rect 2044 8560 2096 8566
rect 2044 8502 2096 8508
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 112 8288 164 8294
rect 112 8230 164 8236
rect 124 7721 152 8230
rect 1676 7744 1728 7750
rect 110 7712 166 7721
rect 1676 7686 1728 7692
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 110 7647 166 7656
rect 1688 7274 1716 7686
rect 1676 7268 1728 7274
rect 1676 7210 1728 7216
rect 1768 7268 1820 7274
rect 1768 7210 1820 7216
rect 1780 6866 1808 7210
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 110 6624 166 6633
rect 166 6582 244 6610
rect 110 6559 166 6568
rect 216 6186 244 6582
rect 1964 6254 1992 7686
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 204 6180 256 6186
rect 204 6122 256 6128
rect 112 6112 164 6118
rect 112 6054 164 6060
rect 124 5409 152 6054
rect 110 5400 166 5409
rect 110 5335 166 5344
rect 20 5296 72 5302
rect 20 5238 72 5244
rect 110 4142 166 4151
rect 110 4077 166 4086
rect 124 3738 152 4077
rect 112 3732 164 3738
rect 112 3674 164 3680
rect 1412 3194 1440 6190
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1780 4282 1808 5646
rect 2056 5234 2084 5850
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1768 4276 1820 4282
rect 1768 4218 1820 4224
rect 1872 4010 1900 4422
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1872 3670 1900 3946
rect 1860 3664 1912 3670
rect 1860 3606 1912 3612
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 112 3052 164 3058
rect 112 2994 164 3000
rect 124 2961 152 2994
rect 110 2952 166 2961
rect 110 2887 166 2896
rect 2240 2650 2268 15846
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 2700 14822 2728 15506
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2608 13802 2636 14350
rect 2596 13796 2648 13802
rect 2596 13738 2648 13744
rect 2700 12986 2728 14758
rect 2792 13734 2820 15914
rect 2884 15706 2912 15982
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 2976 15162 3004 15506
rect 4724 15366 4752 15982
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 4724 15026 4752 15302
rect 4956 15260 5252 15280
rect 5012 15258 5036 15260
rect 5092 15258 5116 15260
rect 5172 15258 5196 15260
rect 5034 15206 5036 15258
rect 5098 15206 5110 15258
rect 5172 15206 5174 15258
rect 5012 15204 5036 15206
rect 5092 15204 5116 15206
rect 5172 15204 5196 15206
rect 4956 15184 5252 15204
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 4448 14482 4476 14894
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3804 13938 3832 14214
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 3148 13796 3200 13802
rect 3148 13738 3200 13744
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2976 12850 3004 13126
rect 3056 12912 3108 12918
rect 3056 12854 3108 12860
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 3068 12442 3096 12854
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2792 11694 2820 12038
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2596 11076 2648 11082
rect 2596 11018 2648 11024
rect 2608 10742 2636 11018
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2332 8906 2360 9590
rect 2320 8900 2372 8906
rect 2320 8842 2372 8848
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 2332 7886 2360 8842
rect 2884 8634 2912 8842
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3160 8566 3188 13738
rect 3804 13530 3832 13874
rect 4448 13814 4476 14418
rect 4356 13786 4476 13814
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 3700 13184 3752 13190
rect 3700 13126 3752 13132
rect 3712 12782 3740 13126
rect 4080 12986 4108 13330
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 4080 12306 4108 12582
rect 4264 12374 4292 13330
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3620 10606 3648 11494
rect 4080 11286 4108 12242
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4172 11354 4200 11630
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 4264 10606 4292 12310
rect 4356 11218 4384 13786
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4448 12918 4476 13670
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4448 12374 4476 12854
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4436 12368 4488 12374
rect 4436 12310 4488 12316
rect 4448 11558 4476 12310
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4356 10674 4384 11154
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 3620 10266 3648 10542
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 3804 9722 3832 10134
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 4080 9586 4108 10202
rect 4160 10192 4212 10198
rect 4264 10180 4292 10542
rect 4212 10152 4292 10180
rect 4160 10134 4212 10140
rect 4356 10130 4384 10610
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4356 9722 4384 10066
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3436 9489 3464 9522
rect 3422 9480 3478 9489
rect 3422 9415 3478 9424
rect 3436 9382 3464 9415
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 3148 8560 3200 8566
rect 3148 8502 3200 8508
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 2412 8016 2464 8022
rect 2412 7958 2464 7964
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2332 7002 2360 7822
rect 2424 7546 2452 7958
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2424 6866 2452 7482
rect 2516 7410 2544 7822
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 3068 7206 3096 8230
rect 3620 7750 3648 8434
rect 3896 8090 3924 8978
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2424 6322 2452 6802
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 2976 5370 3004 5714
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2424 4842 2452 4966
rect 2424 4826 2544 4842
rect 2424 4820 2556 4826
rect 2424 4814 2504 4820
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2332 4282 2360 4558
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2332 3738 2360 4218
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 2332 3058 2360 3538
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 2332 2961 2360 2994
rect 2318 2952 2374 2961
rect 2318 2887 2374 2896
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 1860 2508 1912 2514
rect 1860 2450 1912 2456
rect 1032 2372 1084 2378
rect 1032 2314 1084 2320
rect 754 82 810 480
rect 1044 82 1072 2314
rect 1872 2281 1900 2450
rect 1858 2272 1914 2281
rect 1858 2207 1914 2216
rect 754 54 1072 82
rect 2318 82 2374 480
rect 2424 82 2452 4814
rect 2504 4762 2556 4768
rect 2976 4758 3004 5306
rect 3068 4826 3096 7142
rect 3160 7002 3188 7278
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3620 6118 3648 7686
rect 3712 6458 3740 7686
rect 4356 6866 4384 9658
rect 4448 9382 4476 11494
rect 4540 11218 4568 12718
rect 4632 11898 4660 14894
rect 5644 14550 5672 14894
rect 5828 14550 5856 20198
rect 6196 18426 6224 23582
rect 8390 23582 8524 23610
rect 8390 23520 8446 23582
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8312 19174 8340 19654
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 6920 18828 6972 18834
rect 6920 18770 6972 18776
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5920 17678 5948 18226
rect 6196 18222 6224 18362
rect 6932 18358 6960 18770
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 5908 17672 5960 17678
rect 5908 17614 5960 17620
rect 5920 17202 5948 17614
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 6012 16998 6040 17750
rect 7944 17678 7972 18022
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 7932 17672 7984 17678
rect 7932 17614 7984 17620
rect 7944 17270 7972 17614
rect 7932 17264 7984 17270
rect 7932 17206 7984 17212
rect 8036 17134 8064 17750
rect 8128 17202 8156 18566
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8220 17338 8248 18022
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8116 17196 8168 17202
rect 8116 17138 8168 17144
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 6012 16726 6040 16934
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 8024 16720 8076 16726
rect 8024 16662 8076 16668
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 7116 15978 7144 16390
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7104 15972 7156 15978
rect 7104 15914 7156 15920
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6564 15638 6592 15846
rect 7116 15706 7144 15914
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 7196 15632 7248 15638
rect 7196 15574 7248 15580
rect 6092 15564 6144 15570
rect 6092 15506 6144 15512
rect 6104 15162 6132 15506
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6840 14958 6868 15302
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 5632 14544 5684 14550
rect 5632 14486 5684 14492
rect 5816 14544 5868 14550
rect 5816 14486 5868 14492
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 4956 14172 5252 14192
rect 5012 14170 5036 14172
rect 5092 14170 5116 14172
rect 5172 14170 5196 14172
rect 5034 14118 5036 14170
rect 5098 14118 5110 14170
rect 5172 14118 5174 14170
rect 5012 14116 5036 14118
rect 5092 14116 5116 14118
rect 5172 14116 5196 14118
rect 4956 14096 5252 14116
rect 5368 14074 5396 14350
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5736 13734 5764 14418
rect 5828 14074 5856 14486
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5736 13190 5764 13670
rect 6288 13530 6316 14758
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 6840 13870 6868 14486
rect 7116 14346 7144 15438
rect 7208 15162 7236 15574
rect 7392 15502 7420 16050
rect 8036 15910 8064 16662
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 8036 14890 8064 15846
rect 8024 14884 8076 14890
rect 8024 14826 8076 14832
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6840 13530 6868 13806
rect 7564 13796 7616 13802
rect 7564 13738 7616 13744
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 4956 13084 5252 13104
rect 5012 13082 5036 13084
rect 5092 13082 5116 13084
rect 5172 13082 5196 13084
rect 5034 13030 5036 13082
rect 5098 13030 5110 13082
rect 5172 13030 5174 13082
rect 5012 13028 5036 13030
rect 5092 13028 5116 13030
rect 5172 13028 5196 13030
rect 4956 13008 5252 13028
rect 5736 12782 5764 13126
rect 5920 12850 5948 13262
rect 6288 12918 6316 13466
rect 7576 13462 7604 13738
rect 7564 13456 7616 13462
rect 7564 13398 7616 13404
rect 7378 13288 7434 13297
rect 7378 13223 7434 13232
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6368 12912 6420 12918
rect 6368 12854 6420 12860
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5092 12442 5120 12718
rect 5460 12646 5488 12718
rect 6288 12714 6316 12854
rect 6276 12708 6328 12714
rect 6276 12650 6328 12656
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 4956 11996 5252 12016
rect 5012 11994 5036 11996
rect 5092 11994 5116 11996
rect 5172 11994 5196 11996
rect 5034 11942 5036 11994
rect 5098 11942 5110 11994
rect 5172 11942 5174 11994
rect 5012 11940 5036 11942
rect 5092 11940 5116 11942
rect 5172 11940 5196 11942
rect 4956 11920 5252 11940
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4724 11558 4752 11698
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4724 11354 4752 11494
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4540 10810 4568 11154
rect 4816 10810 4844 11766
rect 5368 11694 5396 12038
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 4956 10908 5252 10928
rect 5012 10906 5036 10908
rect 5092 10906 5116 10908
rect 5172 10906 5196 10908
rect 5034 10854 5036 10906
rect 5098 10854 5110 10906
rect 5172 10854 5174 10906
rect 5012 10852 5036 10854
rect 5092 10852 5116 10854
rect 5172 10852 5196 10854
rect 4956 10832 5252 10852
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4448 8362 4476 9318
rect 4632 9178 4660 9454
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 3700 6452 3752 6458
rect 3700 6394 3752 6400
rect 4264 6254 4292 6734
rect 4356 6390 4384 6802
rect 4724 6798 4752 7142
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 3792 6248 3844 6254
rect 3792 6190 3844 6196
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3804 5370 3832 6190
rect 4264 5846 4292 6190
rect 4252 5840 4304 5846
rect 4252 5782 4304 5788
rect 4356 5778 4384 6326
rect 4632 5778 4660 6666
rect 4724 6458 4752 6734
rect 4816 6662 4844 10746
rect 5368 10674 5396 11290
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 4956 9820 5252 9840
rect 5012 9818 5036 9820
rect 5092 9818 5116 9820
rect 5172 9818 5196 9820
rect 5034 9766 5036 9818
rect 5098 9766 5110 9818
rect 5172 9766 5174 9818
rect 5012 9764 5036 9766
rect 5092 9764 5116 9766
rect 5172 9764 5196 9766
rect 4956 9744 5252 9764
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5276 9178 5304 9318
rect 5264 9172 5316 9178
rect 5316 9132 5396 9160
rect 5264 9114 5316 9120
rect 4956 8732 5252 8752
rect 5012 8730 5036 8732
rect 5092 8730 5116 8732
rect 5172 8730 5196 8732
rect 5034 8678 5036 8730
rect 5098 8678 5110 8730
rect 5172 8678 5174 8730
rect 5012 8676 5036 8678
rect 5092 8676 5116 8678
rect 5172 8676 5196 8678
rect 4956 8656 5252 8676
rect 5368 8362 5396 9132
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5368 7954 5396 8298
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 4956 7644 5252 7664
rect 5012 7642 5036 7644
rect 5092 7642 5116 7644
rect 5172 7642 5196 7644
rect 5034 7590 5036 7642
rect 5098 7590 5110 7642
rect 5172 7590 5174 7642
rect 5012 7588 5036 7590
rect 5092 7588 5116 7590
rect 5172 7588 5196 7590
rect 4956 7568 5252 7588
rect 5460 7478 5488 10950
rect 5552 10538 5580 12242
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 5644 10810 5672 12174
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 5736 11626 5764 12038
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5736 11286 5764 11562
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5814 11112 5870 11121
rect 5814 11047 5870 11056
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5552 10266 5580 10474
rect 5644 10266 5672 10746
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5828 10130 5856 11047
rect 6104 11014 6132 12038
rect 6288 11558 6316 12174
rect 6380 12170 6408 12854
rect 6748 12782 6776 13126
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6288 11150 6316 11494
rect 6380 11218 6408 11630
rect 6472 11558 6500 12582
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6564 11354 6592 12718
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6288 10470 6316 11086
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5644 8634 5672 8910
rect 5736 8906 5764 9862
rect 5828 9722 5856 10066
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 6092 9104 6144 9110
rect 6144 9064 6224 9092
rect 6092 9046 6144 9052
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5920 8362 5948 8842
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 5092 6866 5120 7142
rect 5460 7002 5488 7414
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5736 6866 5764 7482
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4956 6556 5252 6576
rect 5012 6554 5036 6556
rect 5092 6554 5116 6556
rect 5172 6554 5196 6556
rect 5034 6502 5036 6554
rect 5098 6502 5110 6554
rect 5172 6502 5174 6554
rect 5012 6500 5036 6502
rect 5092 6500 5116 6502
rect 5172 6500 5196 6502
rect 4956 6480 5252 6500
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3804 5166 3832 5306
rect 4356 5234 4384 5714
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4632 5166 4660 5714
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 2964 4752 3016 4758
rect 2964 4694 3016 4700
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2516 4146 2544 4558
rect 2976 4214 3004 4694
rect 3988 4622 4016 4966
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2516 2990 2544 4082
rect 3804 4010 3832 4422
rect 3792 4004 3844 4010
rect 3792 3946 3844 3952
rect 3804 3194 3832 3946
rect 3988 3738 4016 4558
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 2318 54 2452 82
rect 3882 82 3938 480
rect 4172 82 4200 5034
rect 4632 4826 4660 5102
rect 4816 5098 4844 6190
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 5368 5710 5396 6122
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 4956 5468 5252 5488
rect 5012 5466 5036 5468
rect 5092 5466 5116 5468
rect 5172 5466 5196 5468
rect 5034 5414 5036 5466
rect 5098 5414 5110 5466
rect 5172 5414 5174 5466
rect 5012 5412 5036 5414
rect 5092 5412 5116 5414
rect 5172 5412 5196 5414
rect 4956 5392 5252 5412
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5000 4826 5028 4966
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4264 4282 4292 4694
rect 4956 4380 5252 4400
rect 5012 4378 5036 4380
rect 5092 4378 5116 4380
rect 5172 4378 5196 4380
rect 5034 4326 5036 4378
rect 5098 4326 5110 4378
rect 5172 4326 5174 4378
rect 5012 4324 5036 4326
rect 5092 4324 5116 4326
rect 5172 4324 5196 4326
rect 4956 4304 5252 4324
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4540 2514 4568 3470
rect 4632 3058 4660 3606
rect 4816 3534 4844 4150
rect 5368 4146 5396 4966
rect 5828 4690 5856 5646
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5828 3942 5856 4626
rect 5920 4078 5948 8298
rect 6196 8294 6224 9064
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6196 8022 6224 8230
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6288 7410 6316 10406
rect 6380 10062 6408 11154
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6564 10810 6592 10950
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6380 9926 6408 9998
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6196 6458 6224 6598
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 6012 5098 6040 5714
rect 6196 5370 6224 6394
rect 6380 6186 6408 9862
rect 6656 8838 6684 12582
rect 6748 11082 6776 12718
rect 7392 12306 7420 13223
rect 7576 12986 7604 13398
rect 8036 13326 8064 14214
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8116 13252 8168 13258
rect 8116 13194 8168 13200
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 8128 12646 8156 13194
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7300 11694 7328 12038
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7116 11286 7144 11630
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6840 9586 6868 9930
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6932 9178 6960 11018
rect 7116 11014 7144 11222
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7116 10130 7144 10950
rect 7300 10130 7328 11630
rect 7392 11354 7420 12242
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7300 9722 7328 10066
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 7300 7954 7328 9658
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7576 7954 7604 9590
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7300 7546 7328 7890
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6656 6866 6684 7142
rect 7300 7002 7328 7482
rect 7484 7206 7512 7822
rect 7576 7410 7604 7890
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6368 6180 6420 6186
rect 6368 6122 6420 6128
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6288 5166 6316 5714
rect 6656 5574 6684 6802
rect 7300 6254 7328 6938
rect 7484 6934 7512 7142
rect 7472 6928 7524 6934
rect 7472 6870 7524 6876
rect 7484 6322 7512 6870
rect 7576 6338 7604 7346
rect 7668 7002 7696 12038
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7852 11558 7880 11630
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7760 10266 7788 10542
rect 7852 10538 7880 11154
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7944 10742 7972 11086
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7748 10124 7800 10130
rect 7852 10112 7880 10474
rect 8036 10470 8064 10950
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 7800 10084 7880 10112
rect 7748 10066 7800 10072
rect 7748 9376 7800 9382
rect 7852 9364 7880 10084
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7944 9654 7972 10066
rect 7932 9648 7984 9654
rect 7932 9590 7984 9596
rect 7800 9336 7880 9364
rect 7748 9318 7800 9324
rect 7760 7478 7788 9318
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7852 8430 7880 8774
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7852 8090 7880 8366
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7472 6316 7524 6322
rect 7576 6310 7696 6338
rect 7472 6258 7524 6264
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6276 5160 6328 5166
rect 6276 5102 6328 5108
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 6012 4826 6040 5034
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6840 4758 6868 5170
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6840 4154 6868 4694
rect 6748 4126 6868 4154
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4956 3292 5252 3312
rect 5012 3290 5036 3292
rect 5092 3290 5116 3292
rect 5172 3290 5196 3292
rect 5034 3238 5036 3290
rect 5098 3238 5110 3290
rect 5172 3238 5174 3290
rect 5012 3236 5036 3238
rect 5092 3236 5116 3238
rect 5172 3236 5196 3238
rect 4956 3216 5252 3236
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4540 2417 4568 2450
rect 4526 2408 4582 2417
rect 4526 2343 4582 2352
rect 4956 2204 5252 2224
rect 5012 2202 5036 2204
rect 5092 2202 5116 2204
rect 5172 2202 5196 2204
rect 5034 2150 5036 2202
rect 5098 2150 5110 2202
rect 5172 2150 5174 2202
rect 5012 2148 5036 2150
rect 5092 2148 5116 2150
rect 5172 2148 5196 2150
rect 4956 2128 5252 2148
rect 3882 54 4200 82
rect 5538 82 5594 480
rect 5828 82 5856 3878
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 6012 2582 6040 2858
rect 6000 2576 6052 2582
rect 6000 2518 6052 2524
rect 6748 1193 6776 4126
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6840 2922 6868 3334
rect 6828 2916 6880 2922
rect 6828 2858 6880 2864
rect 6932 2854 6960 3538
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6734 1184 6790 1193
rect 6734 1119 6790 1128
rect 5538 54 5856 82
rect 6932 82 6960 2790
rect 7208 2514 7236 6190
rect 7300 5370 7328 6190
rect 7576 6118 7604 6190
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7668 4690 7696 6310
rect 7760 5166 7788 7414
rect 7944 6254 7972 8978
rect 8036 8362 8064 10406
rect 8128 8945 8156 12582
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8220 10062 8248 10950
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8114 8936 8170 8945
rect 8114 8871 8170 8880
rect 8312 8566 8340 19110
rect 8496 18970 8524 23582
rect 10704 23582 10838 23610
rect 8956 21244 9252 21264
rect 9012 21242 9036 21244
rect 9092 21242 9116 21244
rect 9172 21242 9196 21244
rect 9034 21190 9036 21242
rect 9098 21190 9110 21242
rect 9172 21190 9174 21242
rect 9012 21188 9036 21190
rect 9092 21188 9116 21190
rect 9172 21188 9196 21190
rect 8956 21168 9252 21188
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 8956 20156 9252 20176
rect 9012 20154 9036 20156
rect 9092 20154 9116 20156
rect 9172 20154 9196 20156
rect 9034 20102 9036 20154
rect 9098 20102 9110 20154
rect 9172 20102 9174 20154
rect 9012 20100 9036 20102
rect 9092 20100 9116 20102
rect 9172 20100 9196 20102
rect 8956 20080 9252 20100
rect 8956 19068 9252 19088
rect 9012 19066 9036 19068
rect 9092 19066 9116 19068
rect 9172 19066 9196 19068
rect 9034 19014 9036 19066
rect 9098 19014 9110 19066
rect 9172 19014 9174 19066
rect 9012 19012 9036 19014
rect 9092 19012 9116 19014
rect 9172 19012 9196 19014
rect 8956 18992 9252 19012
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8404 18154 8432 18566
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8392 18148 8444 18154
rect 8392 18090 8444 18096
rect 8404 17785 8432 18090
rect 8390 17776 8446 17785
rect 8390 17711 8446 17720
rect 8680 17678 8708 18226
rect 8956 17980 9252 18000
rect 9012 17978 9036 17980
rect 9092 17978 9116 17980
rect 9172 17978 9196 17980
rect 9034 17926 9036 17978
rect 9098 17926 9110 17978
rect 9172 17926 9174 17978
rect 9012 17924 9036 17926
rect 9092 17924 9116 17926
rect 9172 17924 9196 17926
rect 8956 17904 9252 17924
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8404 16794 8432 17070
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8404 15910 8432 16526
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8404 11898 8432 15846
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8496 11744 8524 12038
rect 8404 11716 8524 11744
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8220 6458 8248 6870
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5778 7880 6054
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7852 4826 7880 5714
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7944 4214 7972 6190
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8036 5370 8064 5850
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8036 4282 8064 5306
rect 8128 5234 8156 6326
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 8128 3058 8156 5034
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7760 2553 7788 2790
rect 7746 2544 7802 2553
rect 7196 2508 7248 2514
rect 8312 2514 8340 3878
rect 8404 3738 8432 11716
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10810 8524 10950
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8496 9994 8524 10746
rect 8680 10198 8708 17614
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8772 11286 8800 14554
rect 8864 13938 8892 17818
rect 8956 16892 9252 16912
rect 9012 16890 9036 16892
rect 9092 16890 9116 16892
rect 9172 16890 9196 16892
rect 9034 16838 9036 16890
rect 9098 16838 9110 16890
rect 9172 16838 9174 16890
rect 9012 16836 9036 16838
rect 9092 16836 9116 16838
rect 9172 16836 9196 16838
rect 8956 16816 9252 16836
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 8956 15804 9252 15824
rect 9012 15802 9036 15804
rect 9092 15802 9116 15804
rect 9172 15802 9196 15804
rect 9034 15750 9036 15802
rect 9098 15750 9110 15802
rect 9172 15750 9174 15802
rect 9012 15748 9036 15750
rect 9092 15748 9116 15750
rect 9172 15748 9196 15750
rect 8956 15728 9252 15748
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 8956 15065 8984 15098
rect 8942 15056 8998 15065
rect 9784 15026 9812 15982
rect 8942 14991 8998 15000
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 8956 14716 9252 14736
rect 9012 14714 9036 14716
rect 9092 14714 9116 14716
rect 9172 14714 9196 14716
rect 9034 14662 9036 14714
rect 9098 14662 9110 14714
rect 9172 14662 9174 14714
rect 9012 14660 9036 14662
rect 9092 14660 9116 14662
rect 9172 14660 9196 14662
rect 8956 14640 9252 14660
rect 9324 14618 9352 14894
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9416 14550 9444 14758
rect 9404 14544 9456 14550
rect 9404 14486 9456 14492
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8864 13530 8892 13874
rect 9416 13841 9444 14486
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9402 13832 9458 13841
rect 9312 13796 9364 13802
rect 9402 13767 9458 13776
rect 9678 13832 9734 13841
rect 9678 13767 9734 13776
rect 9312 13738 9364 13744
rect 8956 13628 9252 13648
rect 9012 13626 9036 13628
rect 9092 13626 9116 13628
rect 9172 13626 9196 13628
rect 9034 13574 9036 13626
rect 9098 13574 9110 13626
rect 9172 13574 9174 13626
rect 9012 13572 9036 13574
rect 9092 13572 9116 13574
rect 9172 13572 9196 13574
rect 8956 13552 9252 13572
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 9324 12986 9352 13738
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 8956 12540 9252 12560
rect 9012 12538 9036 12540
rect 9092 12538 9116 12540
rect 9172 12538 9196 12540
rect 9034 12486 9036 12538
rect 9098 12486 9110 12538
rect 9172 12486 9174 12538
rect 9012 12484 9036 12486
rect 9092 12484 9116 12486
rect 9172 12484 9196 12486
rect 8956 12464 9252 12484
rect 9324 12442 9352 12786
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9692 12306 9720 13767
rect 9784 13462 9812 14214
rect 9864 13796 9916 13802
rect 9864 13738 9916 13744
rect 9772 13456 9824 13462
rect 9772 13398 9824 13404
rect 9876 13326 9904 13738
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9692 11694 9720 12242
rect 9784 12102 9812 13262
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9692 11558 9720 11630
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 8956 11452 9252 11472
rect 9012 11450 9036 11452
rect 9092 11450 9116 11452
rect 9172 11450 9196 11452
rect 9034 11398 9036 11450
rect 9098 11398 9110 11450
rect 9172 11398 9174 11450
rect 9012 11396 9036 11398
rect 9092 11396 9116 11398
rect 9172 11396 9196 11398
rect 8956 11376 9252 11396
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9416 11014 9444 11154
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9416 10674 9444 10950
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 8956 10364 9252 10384
rect 9012 10362 9036 10364
rect 9092 10362 9116 10364
rect 9172 10362 9196 10364
rect 9034 10310 9036 10362
rect 9098 10310 9110 10362
rect 9172 10310 9174 10362
rect 9012 10308 9036 10310
rect 9092 10308 9116 10310
rect 9172 10308 9196 10310
rect 8956 10288 9252 10308
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8588 9450 8616 9998
rect 9416 9586 9444 10610
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9600 10198 9628 10474
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8496 9178 8524 9386
rect 8956 9276 9252 9296
rect 9012 9274 9036 9276
rect 9092 9274 9116 9276
rect 9172 9274 9196 9276
rect 9034 9222 9036 9274
rect 9098 9222 9110 9274
rect 9172 9222 9174 9274
rect 9012 9220 9036 9222
rect 9092 9220 9116 9222
rect 9172 9220 9196 9222
rect 8956 9200 9252 9220
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 9692 9042 9720 11494
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 10130 9812 10406
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9784 9722 9812 10066
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9968 9674 9996 20742
rect 10704 20602 10732 23582
rect 10782 23520 10838 23582
rect 12820 23582 13230 23610
rect 11152 21412 11204 21418
rect 11152 21354 11204 21360
rect 11164 21010 11192 21354
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 11164 20602 11192 20946
rect 12820 20602 12848 23582
rect 13174 23520 13230 23582
rect 15566 23610 15622 24000
rect 17958 23610 18014 24000
rect 20350 23610 20406 24000
rect 22742 23610 22798 24000
rect 15566 23582 15700 23610
rect 15566 23520 15622 23582
rect 12956 21788 13252 21808
rect 13012 21786 13036 21788
rect 13092 21786 13116 21788
rect 13172 21786 13196 21788
rect 13034 21734 13036 21786
rect 13098 21734 13110 21786
rect 13172 21734 13174 21786
rect 13012 21732 13036 21734
rect 13092 21732 13116 21734
rect 13172 21732 13196 21734
rect 12956 21712 13252 21732
rect 12956 20700 13252 20720
rect 13012 20698 13036 20700
rect 13092 20698 13116 20700
rect 13172 20698 13196 20700
rect 13034 20646 13036 20698
rect 13098 20646 13110 20698
rect 13172 20646 13174 20698
rect 13012 20644 13036 20646
rect 13092 20644 13116 20646
rect 13172 20644 13196 20646
rect 12956 20624 13252 20644
rect 10692 20596 10744 20602
rect 10692 20538 10744 20544
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10612 18426 10640 18702
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10152 17202 10180 17614
rect 10244 17338 10272 17750
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 10324 17060 10376 17066
rect 10324 17002 10376 17008
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 10060 15434 10088 15914
rect 10152 15706 10180 16594
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10048 15428 10100 15434
rect 10048 15370 10100 15376
rect 10060 15026 10088 15370
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 10152 14958 10180 15642
rect 10244 15570 10272 16526
rect 10336 16454 10364 17002
rect 10416 16720 10468 16726
rect 10416 16662 10468 16668
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10244 15094 10272 15506
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10060 14074 10088 14418
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10060 12986 10088 14010
rect 10232 13456 10284 13462
rect 10232 13398 10284 13404
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10048 12300 10100 12306
rect 10152 12288 10180 13126
rect 10244 12986 10272 13398
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 10100 12260 10180 12288
rect 10048 12242 10100 12248
rect 10060 11898 10088 12242
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10232 11824 10284 11830
rect 10232 11766 10284 11772
rect 10048 11620 10100 11626
rect 10048 11562 10100 11568
rect 10060 11218 10088 11562
rect 10244 11354 10272 11766
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10244 10130 10272 11290
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 9968 9646 10272 9674
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9404 8560 9456 8566
rect 9404 8502 9456 8508
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8680 7546 8708 8230
rect 8956 8188 9252 8208
rect 9012 8186 9036 8188
rect 9092 8186 9116 8188
rect 9172 8186 9196 8188
rect 9034 8134 9036 8186
rect 9098 8134 9110 8186
rect 9172 8134 9174 8186
rect 9012 8132 9036 8134
rect 9092 8132 9116 8134
rect 9172 8132 9196 8134
rect 8956 8112 9252 8132
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8496 5234 8524 6666
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8588 5914 8616 6394
rect 8680 6186 8708 7346
rect 8864 7274 8892 7686
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8956 7274 8984 7482
rect 9416 7478 9444 8502
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9692 8022 9720 8298
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9784 7546 9812 7890
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 8944 7268 8996 7274
rect 8944 7210 8996 7216
rect 8864 6798 8892 7210
rect 8956 7100 9252 7120
rect 9012 7098 9036 7100
rect 9092 7098 9116 7100
rect 9172 7098 9196 7100
rect 9034 7046 9036 7098
rect 9098 7046 9110 7098
rect 9172 7046 9174 7098
rect 9012 7044 9036 7046
rect 9092 7044 9116 7046
rect 9172 7044 9196 7046
rect 8956 7024 9252 7044
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8772 6186 8800 6598
rect 8864 6322 8892 6734
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 9140 6186 9168 6734
rect 9968 6458 9996 6802
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 8680 5914 8708 6122
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8680 5370 8708 5850
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8496 4826 8524 5170
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8496 2854 8524 3538
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 7746 2479 7802 2488
rect 8300 2508 8352 2514
rect 7196 2450 7248 2456
rect 7760 2446 7788 2479
rect 8300 2450 8352 2456
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7102 82 7158 480
rect 6932 54 7158 82
rect 8496 82 8524 2790
rect 8772 2009 8800 6122
rect 8956 6012 9252 6032
rect 9012 6010 9036 6012
rect 9092 6010 9116 6012
rect 9172 6010 9196 6012
rect 9034 5958 9036 6010
rect 9098 5958 9110 6010
rect 9172 5958 9174 6010
rect 9012 5956 9036 5958
rect 9092 5956 9116 5958
rect 9172 5956 9196 5958
rect 8956 5936 9252 5956
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5370 9444 5510
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9496 5024 9548 5030
rect 9772 5024 9824 5030
rect 9496 4966 9548 4972
rect 9692 4984 9772 5012
rect 8956 4924 9252 4944
rect 9012 4922 9036 4924
rect 9092 4922 9116 4924
rect 9172 4922 9196 4924
rect 9034 4870 9036 4922
rect 9098 4870 9110 4922
rect 9172 4870 9174 4922
rect 9012 4868 9036 4870
rect 9092 4868 9116 4870
rect 9172 4868 9196 4870
rect 8956 4848 9252 4868
rect 9508 4622 9536 4966
rect 9692 4690 9720 4984
rect 9772 4966 9824 4972
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9508 4078 9536 4558
rect 9692 4282 9720 4626
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 10152 4078 10180 4490
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 8956 3836 9252 3856
rect 9012 3834 9036 3836
rect 9092 3834 9116 3836
rect 9172 3834 9196 3836
rect 9034 3782 9036 3834
rect 9098 3782 9110 3834
rect 9172 3782 9174 3834
rect 9012 3780 9036 3782
rect 9092 3780 9116 3782
rect 9172 3780 9196 3782
rect 8956 3760 9252 3780
rect 9324 3738 9352 3946
rect 10060 3738 10088 3946
rect 10152 3738 10180 4014
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 8956 2748 9252 2768
rect 9012 2746 9036 2748
rect 9092 2746 9116 2748
rect 9172 2746 9196 2748
rect 9034 2694 9036 2746
rect 9098 2694 9110 2746
rect 9172 2694 9174 2746
rect 9012 2692 9036 2694
rect 9092 2692 9116 2694
rect 9172 2692 9196 2694
rect 8956 2672 9252 2692
rect 9416 2650 9444 2790
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 9876 2582 9904 3334
rect 10060 3194 10088 3674
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10244 3058 10272 9646
rect 10336 7993 10364 16390
rect 10428 15910 10456 16662
rect 10520 16250 10548 17274
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10428 14600 10456 15846
rect 10508 14612 10560 14618
rect 10428 14572 10508 14600
rect 10508 14554 10560 14560
rect 10520 14414 10548 14554
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10520 12782 10548 14350
rect 10704 13814 10732 20198
rect 12452 20058 12480 20334
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 11704 19916 11756 19922
rect 11704 19858 11756 19864
rect 11716 19514 11744 19858
rect 12956 19612 13252 19632
rect 13012 19610 13036 19612
rect 13092 19610 13116 19612
rect 13172 19610 13196 19612
rect 13034 19558 13036 19610
rect 13098 19558 13110 19610
rect 13172 19558 13174 19610
rect 13012 19556 13036 19558
rect 13092 19556 13116 19558
rect 13172 19556 13196 19558
rect 12956 19536 13252 19556
rect 15672 19514 15700 23582
rect 17696 23582 18014 23610
rect 16956 21244 17252 21264
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17034 21190 17036 21242
rect 17098 21190 17110 21242
rect 17172 21190 17174 21242
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 16956 21168 17252 21188
rect 17696 20602 17724 23582
rect 17958 23520 18014 23582
rect 20088 23582 20406 23610
rect 17684 20596 17736 20602
rect 17684 20538 17736 20544
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 10980 18630 11008 19246
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11164 18902 11192 19110
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10980 18154 11008 18566
rect 11164 18426 11192 18838
rect 11716 18698 11744 19450
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11716 18290 11744 18634
rect 12956 18524 13252 18544
rect 13012 18522 13036 18524
rect 13092 18522 13116 18524
rect 13172 18522 13196 18524
rect 13034 18470 13036 18522
rect 13098 18470 13110 18522
rect 13172 18470 13174 18522
rect 13012 18468 13036 18470
rect 13092 18468 13116 18470
rect 13172 18468 13196 18470
rect 12956 18448 13252 18468
rect 13372 18426 13400 18702
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 10888 17814 10916 18090
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10796 17066 10824 17614
rect 10888 17202 10916 17750
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10980 15706 11008 18090
rect 13372 18086 13400 18362
rect 13648 18290 13676 18770
rect 14844 18426 14872 19110
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13648 17814 13676 18226
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 14292 17814 14320 18090
rect 13636 17808 13688 17814
rect 13636 17750 13688 17756
rect 14280 17808 14332 17814
rect 16040 17785 16068 18566
rect 14280 17750 14332 17756
rect 16026 17776 16082 17785
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11716 17338 11744 17682
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13268 17604 13320 17610
rect 13268 17546 13320 17552
rect 12956 17436 13252 17456
rect 13012 17434 13036 17436
rect 13092 17434 13116 17436
rect 13172 17434 13196 17436
rect 13034 17382 13036 17434
rect 13098 17382 13110 17434
rect 13172 17382 13174 17434
rect 13012 17380 13036 17382
rect 13092 17380 13116 17382
rect 13172 17380 13196 17382
rect 12956 17360 13252 17380
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 13280 17202 13308 17546
rect 13556 17202 13584 17614
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 11888 16720 11940 16726
rect 11888 16662 11940 16668
rect 11900 16250 11928 16662
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 12268 15638 12296 15846
rect 12256 15632 12308 15638
rect 12256 15574 12308 15580
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 10704 13786 10916 13814
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10520 12646 10548 12718
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10428 11558 10456 11698
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10428 9722 10456 11494
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10520 9382 10548 12582
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11218 10732 12038
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10796 11014 10824 11630
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 10470 10824 10950
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10796 9586 10824 10406
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10520 8974 10548 9318
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10612 8634 10640 8978
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10322 7984 10378 7993
rect 10322 7919 10378 7928
rect 10796 7750 10824 9522
rect 10888 9178 10916 13786
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10980 11558 11008 12174
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10980 11132 11008 11494
rect 11060 11144 11112 11150
rect 10980 11104 11060 11132
rect 10980 10742 11008 11104
rect 11060 11086 11112 11092
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10600 7472 10652 7478
rect 10600 7414 10652 7420
rect 10612 7206 10640 7414
rect 10796 7410 10824 7686
rect 10980 7546 11008 10678
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 11072 9722 11100 9998
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10520 5234 10548 6122
rect 10612 5302 10640 7142
rect 10980 7002 11008 7482
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10888 5778 10916 6598
rect 10980 6458 11008 6938
rect 11072 6730 11100 9658
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10980 6254 11008 6394
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10600 5296 10652 5302
rect 10600 5238 10652 5244
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10888 5030 10916 5714
rect 10980 5234 11008 6190
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10980 4826 11008 5170
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10428 3194 10456 3334
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10428 2922 10456 3130
rect 10980 3058 11008 3470
rect 11164 3126 11192 15302
rect 12176 14958 12204 15438
rect 12268 15026 12296 15574
rect 12728 15366 12756 16526
rect 12820 16250 12848 16934
rect 12956 16348 13252 16368
rect 13012 16346 13036 16348
rect 13092 16346 13116 16348
rect 13172 16346 13196 16348
rect 13034 16294 13036 16346
rect 13098 16294 13110 16346
rect 13172 16294 13174 16346
rect 13012 16292 13036 16294
rect 13092 16292 13116 16294
rect 13172 16292 13196 16294
rect 12956 16272 13252 16292
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12820 15706 12848 16186
rect 13464 16182 13492 16934
rect 13556 16794 13584 17138
rect 13648 16998 13676 17750
rect 15384 17740 15436 17746
rect 16026 17711 16082 17720
rect 15384 17682 15436 17688
rect 15396 17338 15424 17682
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12956 15260 13252 15280
rect 13012 15258 13036 15260
rect 13092 15258 13116 15260
rect 13172 15258 13196 15260
rect 13034 15206 13036 15258
rect 13098 15206 13110 15258
rect 13172 15206 13174 15258
rect 13012 15204 13036 15206
rect 13092 15204 13116 15206
rect 13172 15204 13196 15206
rect 12956 15184 13252 15204
rect 13280 15026 13308 15982
rect 14554 15600 14610 15609
rect 14554 15535 14610 15544
rect 14568 15094 14596 15535
rect 14556 15088 14608 15094
rect 14556 15030 14608 15036
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 11992 14482 12020 14826
rect 12176 14550 12204 14894
rect 12452 14618 12480 14894
rect 14384 14618 14412 14894
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 11808 14074 11836 14418
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11992 13814 12020 14418
rect 12956 14172 13252 14192
rect 13012 14170 13036 14172
rect 13092 14170 13116 14172
rect 13172 14170 13196 14172
rect 13034 14118 13036 14170
rect 13098 14118 13110 14170
rect 13172 14118 13174 14170
rect 13012 14116 13036 14118
rect 13092 14116 13116 14118
rect 13172 14116 13196 14118
rect 12956 14096 13252 14116
rect 11992 13786 12204 13814
rect 12176 13734 12204 13786
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11256 12782 11284 13126
rect 11348 12850 11376 13262
rect 11428 12912 11480 12918
rect 11428 12854 11480 12860
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11348 12442 11376 12786
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11440 12306 11468 12854
rect 11532 12714 11560 13466
rect 11624 13326 11652 13670
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11256 11694 11284 12106
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11256 11014 11284 11630
rect 11532 11558 11560 12310
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11532 11286 11560 11494
rect 11716 11286 11744 13670
rect 12452 13190 12480 13670
rect 12544 13530 12572 13738
rect 13464 13734 13492 14418
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14752 14074 14780 14350
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14936 13938 14964 14214
rect 15488 14074 15516 14486
rect 15672 14414 15700 14894
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 15016 13796 15068 13802
rect 15016 13738 15068 13744
rect 13452 13728 13504 13734
rect 13452 13670 13504 13676
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12452 12782 12480 13126
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12820 12442 12848 13262
rect 12956 13084 13252 13104
rect 13012 13082 13036 13084
rect 13092 13082 13116 13084
rect 13172 13082 13196 13084
rect 13034 13030 13036 13082
rect 13098 13030 13110 13082
rect 13172 13030 13174 13082
rect 13012 13028 13036 13030
rect 13092 13028 13116 13030
rect 13172 13028 13196 13030
rect 12956 13008 13252 13028
rect 13280 12850 13308 13398
rect 13464 13326 13492 13670
rect 15028 13394 15056 13738
rect 15488 13530 15516 14010
rect 15672 13938 15700 14350
rect 16500 13938 16528 20198
rect 16956 20156 17252 20176
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17034 20102 17036 20154
rect 17098 20102 17110 20154
rect 17172 20102 17174 20154
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 16956 20080 17252 20100
rect 16956 19068 17252 19088
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17034 19014 17036 19066
rect 17098 19014 17110 19066
rect 17172 19014 17174 19066
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 16956 18992 17252 19012
rect 16956 17980 17252 18000
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17034 17926 17036 17978
rect 17098 17926 17110 17978
rect 17172 17926 17174 17978
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 16956 17904 17252 17924
rect 20088 17746 20116 23582
rect 20350 23520 20406 23582
rect 22480 23582 22798 23610
rect 21638 22672 21694 22681
rect 21638 22607 21694 22616
rect 20956 21788 21252 21808
rect 21012 21786 21036 21788
rect 21092 21786 21116 21788
rect 21172 21786 21196 21788
rect 21034 21734 21036 21786
rect 21098 21734 21110 21786
rect 21172 21734 21174 21786
rect 21012 21732 21036 21734
rect 21092 21732 21116 21734
rect 21172 21732 21196 21734
rect 20956 21712 21252 21732
rect 20956 20700 21252 20720
rect 21012 20698 21036 20700
rect 21092 20698 21116 20700
rect 21172 20698 21196 20700
rect 21034 20646 21036 20698
rect 21098 20646 21110 20698
rect 21172 20646 21174 20698
rect 21012 20644 21036 20646
rect 21092 20644 21116 20646
rect 21172 20644 21196 20646
rect 20956 20624 21252 20644
rect 21652 20602 21680 22607
rect 22480 20602 22508 23582
rect 22742 23520 22798 23582
rect 23570 21856 23626 21865
rect 23570 21791 23626 21800
rect 23584 21418 23612 21791
rect 23572 21412 23624 21418
rect 23572 21354 23624 21360
rect 21640 20596 21692 20602
rect 21640 20538 21692 20544
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 20076 17740 20128 17746
rect 20076 17682 20128 17688
rect 19340 17536 19392 17542
rect 19340 17478 19392 17484
rect 16956 16892 17252 16912
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17034 16838 17036 16890
rect 17098 16838 17110 16890
rect 17172 16838 17174 16890
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 16956 16816 17252 16836
rect 16956 15804 17252 15824
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17034 15750 17036 15802
rect 17098 15750 17110 15802
rect 17172 15750 17174 15802
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 16956 15728 17252 15748
rect 16956 14716 17252 14736
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17034 14662 17036 14714
rect 17098 14662 17110 14714
rect 17172 14662 17174 14714
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 16956 14640 17252 14660
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 16500 13530 16528 13874
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14292 12850 14320 13126
rect 15488 12986 15516 13330
rect 16592 12986 16620 13738
rect 16956 13628 17252 13648
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17034 13574 17036 13626
rect 17098 13574 17110 13626
rect 17172 13574 17174 13626
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 16956 13552 17252 13572
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11900 11898 11928 12038
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 12728 11558 12756 12242
rect 12956 11996 13252 12016
rect 13012 11994 13036 11996
rect 13092 11994 13116 11996
rect 13172 11994 13196 11996
rect 13034 11942 13036 11994
rect 13098 11942 13110 11994
rect 13172 11942 13174 11994
rect 13012 11940 13036 11942
rect 13092 11940 13116 11942
rect 13172 11940 13196 11942
rect 12956 11920 13252 11940
rect 13372 11558 13400 12242
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11256 10538 11284 10950
rect 11244 10532 11296 10538
rect 11244 10474 11296 10480
rect 11256 10062 11284 10474
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11244 9444 11296 9450
rect 11348 9432 11376 10950
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 11704 10464 11756 10470
rect 11888 10464 11940 10470
rect 11704 10406 11756 10412
rect 11808 10424 11888 10452
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11440 9722 11468 9930
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11296 9404 11376 9432
rect 11244 9386 11296 9392
rect 11256 7274 11284 9386
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11256 6866 11284 7210
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11256 5914 11284 6802
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11440 5778 11468 6870
rect 11624 6798 11652 6938
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11440 4758 11468 5714
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11532 4826 11560 5034
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11428 4752 11480 4758
rect 11428 4694 11480 4700
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11256 3738 11284 4558
rect 11348 4282 11376 4626
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11624 3670 11652 3878
rect 11716 3670 11744 10406
rect 11808 10130 11836 10424
rect 11888 10406 11940 10412
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11808 9722 11836 10066
rect 12176 10062 12204 10542
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12176 9722 12204 9998
rect 12452 9926 12480 10610
rect 12544 10470 12572 11154
rect 12728 10606 12756 11494
rect 12956 10908 13252 10928
rect 13012 10906 13036 10908
rect 13092 10906 13116 10908
rect 13172 10906 13196 10908
rect 13034 10854 13036 10906
rect 13098 10854 13110 10906
rect 13172 10854 13174 10906
rect 13012 10852 13036 10854
rect 13092 10852 13116 10854
rect 13172 10852 13196 10854
rect 12956 10832 13252 10852
rect 13372 10674 13400 11494
rect 13464 11286 13492 12650
rect 14292 12374 14320 12786
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 16224 12374 16252 12650
rect 16592 12442 16620 12718
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 16212 12368 16264 12374
rect 16212 12310 16264 12316
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 14200 11830 14228 12242
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 15672 11762 15700 12174
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 13452 11280 13504 11286
rect 13452 11222 13504 11228
rect 13464 10810 13492 11222
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12728 10266 12756 10542
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12452 9654 12480 9862
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11992 8566 12020 8978
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11900 6458 11928 6666
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 12176 5370 12204 6802
rect 12452 6662 12480 7278
rect 12636 7206 12664 7958
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12440 6656 12492 6662
rect 12492 6616 12572 6644
rect 12440 6598 12492 6604
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 10416 2916 10468 2922
rect 10416 2858 10468 2864
rect 10704 2650 10732 2994
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10980 2582 11008 2994
rect 11624 2854 11652 3606
rect 11808 3505 11836 5238
rect 12452 4758 12480 5646
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 12544 4078 12572 6616
rect 12636 6168 12664 7142
rect 12728 6866 12756 10202
rect 12956 9820 13252 9840
rect 13012 9818 13036 9820
rect 13092 9818 13116 9820
rect 13172 9818 13196 9820
rect 13034 9766 13036 9818
rect 13098 9766 13110 9818
rect 13172 9766 13174 9818
rect 13012 9764 13036 9766
rect 13092 9764 13116 9766
rect 13172 9764 13196 9766
rect 12956 9744 13252 9764
rect 13372 9518 13400 10610
rect 13464 10266 13492 10746
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13360 9104 13412 9110
rect 13360 9046 13412 9052
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 12956 8732 13252 8752
rect 13012 8730 13036 8732
rect 13092 8730 13116 8732
rect 13172 8730 13196 8732
rect 13034 8678 13036 8730
rect 13098 8678 13110 8730
rect 13172 8678 13174 8730
rect 13012 8676 13036 8678
rect 13092 8676 13116 8678
rect 13172 8676 13196 8678
rect 12956 8656 13252 8676
rect 13280 8498 13308 8910
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13372 8294 13400 9046
rect 13556 8906 13584 11562
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13832 10198 13860 11494
rect 14016 11218 14044 11630
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 14016 10810 14044 11154
rect 15396 10810 15424 11154
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 14016 10470 14044 10746
rect 14200 10674 14228 10746
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14096 10532 14148 10538
rect 14096 10474 14148 10480
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 14108 10266 14136 10474
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13648 9518 13676 9862
rect 13832 9722 13860 10134
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13924 9654 13952 10202
rect 14384 10198 14412 10610
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14372 10192 14424 10198
rect 14372 10134 14424 10140
rect 14384 9994 14412 10134
rect 14476 10062 14504 10406
rect 15764 10266 15792 12174
rect 16224 11626 16252 12310
rect 16868 12084 16896 13194
rect 17052 12782 17080 13398
rect 17328 13326 17356 13874
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 16956 12540 17252 12560
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17034 12486 17036 12538
rect 17098 12486 17110 12538
rect 17172 12486 17174 12538
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 16956 12464 17252 12484
rect 16948 12096 17000 12102
rect 16868 12056 16948 12084
rect 16948 12038 17000 12044
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 16960 11830 16988 12038
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 18340 11694 18368 12038
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 16212 11620 16264 11626
rect 16212 11562 16264 11568
rect 16956 11452 17252 11472
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17034 11398 17036 11450
rect 17098 11398 17110 11450
rect 17172 11398 17174 11450
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 16956 11376 17252 11396
rect 17880 11286 17908 11630
rect 18420 11620 18472 11626
rect 18420 11562 18472 11568
rect 18432 11354 18460 11562
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 15856 10742 15884 11154
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 17512 10470 17540 11086
rect 17604 10742 17632 11154
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 16956 10364 17252 10384
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17034 10310 17036 10362
rect 17098 10310 17110 10362
rect 17172 10310 17174 10362
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 16956 10288 17252 10308
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 14476 9178 14504 9998
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14752 9178 14780 9454
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12820 7206 12848 7822
rect 12956 7644 13252 7664
rect 13012 7642 13036 7644
rect 13092 7642 13116 7644
rect 13172 7642 13196 7644
rect 13034 7590 13036 7642
rect 13098 7590 13110 7642
rect 13172 7590 13174 7642
rect 13012 7588 13036 7590
rect 13092 7588 13116 7590
rect 13172 7588 13196 7590
rect 12956 7568 13252 7588
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12820 7002 12848 7142
rect 13372 7002 13400 8230
rect 13464 8090 13492 8434
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13556 7274 13584 8842
rect 13832 8566 13860 8842
rect 14568 8634 14596 8910
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13728 8356 13780 8362
rect 13648 8316 13728 8344
rect 13648 7750 13676 8316
rect 13728 8298 13780 8304
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 13544 7268 13596 7274
rect 13544 7210 13596 7216
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13648 6866 13676 7686
rect 14108 7342 14136 7686
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14108 6934 14136 7278
rect 14740 7268 14792 7274
rect 14740 7210 14792 7216
rect 14096 6928 14148 6934
rect 14096 6870 14148 6876
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 12728 6458 12756 6802
rect 12956 6556 13252 6576
rect 13012 6554 13036 6556
rect 13092 6554 13116 6556
rect 13172 6554 13196 6556
rect 13034 6502 13036 6554
rect 13098 6502 13110 6554
rect 13172 6502 13174 6554
rect 13012 6500 13036 6502
rect 13092 6500 13116 6502
rect 13172 6500 13196 6502
rect 12956 6480 13252 6500
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 12716 6180 12768 6186
rect 12636 6140 12716 6168
rect 12636 5846 12664 6140
rect 12716 6122 12768 6128
rect 13268 6112 13320 6118
rect 13268 6054 13320 6060
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12636 5030 12664 5782
rect 12956 5468 13252 5488
rect 13012 5466 13036 5468
rect 13092 5466 13116 5468
rect 13172 5466 13196 5468
rect 13034 5414 13036 5466
rect 13098 5414 13110 5466
rect 13172 5414 13174 5466
rect 13012 5412 13036 5414
rect 13092 5412 13116 5414
rect 13172 5412 13196 5414
rect 12956 5392 13252 5412
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12636 4010 12664 4966
rect 13280 4758 13308 6054
rect 13372 5914 13400 6190
rect 13648 5914 13676 6802
rect 14752 6322 14780 7210
rect 14844 6458 14872 9386
rect 15396 8634 15424 9998
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15396 8294 15424 8570
rect 15672 8498 15700 9114
rect 15856 8974 15884 9590
rect 15948 9382 15976 10066
rect 17512 10062 17540 10406
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17512 9382 17540 9998
rect 17604 9586 17632 10066
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17880 9586 17908 9998
rect 19168 9722 19196 10542
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 15948 9110 15976 9318
rect 16500 9178 16528 9318
rect 16956 9276 17252 9296
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17034 9222 17036 9274
rect 17098 9222 17110 9274
rect 17172 9222 17174 9274
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 16956 9200 17252 9220
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 15936 9104 15988 9110
rect 15936 9046 15988 9052
rect 16580 9104 16632 9110
rect 16580 9046 16632 9052
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15028 8090 15056 8230
rect 15856 8090 15884 8910
rect 16224 8566 16252 8910
rect 16592 8634 16620 9046
rect 17130 8936 17186 8945
rect 17224 8900 17276 8906
rect 17186 8880 17224 8888
rect 17130 8871 17224 8880
rect 17144 8860 17224 8871
rect 17224 8842 17276 8848
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16212 8560 16264 8566
rect 16212 8502 16264 8508
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15028 6662 15056 8026
rect 16224 7954 16252 8502
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 15396 7546 15424 7890
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14752 5914 14780 6258
rect 14844 6186 14872 6394
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 13372 5370 13400 5850
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13372 5080 13400 5306
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13452 5092 13504 5098
rect 13372 5052 13452 5080
rect 13452 5034 13504 5040
rect 13832 4758 13860 5170
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12820 4282 12848 4558
rect 12956 4380 13252 4400
rect 13012 4378 13036 4380
rect 13092 4378 13116 4380
rect 13172 4378 13196 4380
rect 13034 4326 13036 4378
rect 13098 4326 13110 4378
rect 13172 4326 13174 4378
rect 13012 4324 13036 4326
rect 13092 4324 13116 4326
rect 13172 4324 13196 4326
rect 12956 4304 13252 4324
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 13280 4214 13308 4694
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 11794 3496 11850 3505
rect 11794 3431 11850 3440
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 9876 2446 9904 2518
rect 11624 2514 11652 2790
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9956 2372 10008 2378
rect 9956 2314 10008 2320
rect 8758 2000 8814 2009
rect 8758 1935 8814 1944
rect 8758 82 8814 480
rect 8496 54 8814 82
rect 9968 82 9996 2314
rect 10322 82 10378 480
rect 9968 54 10378 82
rect 11808 82 11836 3334
rect 12544 3058 12572 3674
rect 13832 3602 13860 4694
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14476 4078 14504 4422
rect 15304 4282 15332 4558
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 15488 4010 15516 4762
rect 15476 4004 15528 4010
rect 15476 3946 15528 3952
rect 13452 3596 13504 3602
rect 13452 3538 13504 3544
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12820 3058 12848 3470
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 12956 3292 13252 3312
rect 13012 3290 13036 3292
rect 13092 3290 13116 3292
rect 13172 3290 13196 3292
rect 13034 3238 13036 3290
rect 13098 3238 13110 3290
rect 13172 3238 13174 3290
rect 13012 3236 13036 3238
rect 13092 3236 13116 3238
rect 13172 3236 13196 3238
rect 12956 3216 13252 3236
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 12636 2582 12664 2858
rect 12624 2576 12676 2582
rect 12624 2518 12676 2524
rect 12820 2514 12848 2994
rect 13372 2961 13400 3334
rect 13464 3194 13492 3538
rect 13832 3194 13860 3538
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15488 3194 15516 3470
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 13358 2952 13414 2961
rect 13358 2887 13414 2896
rect 15580 2514 15608 7686
rect 16316 6798 16344 8230
rect 16956 8188 17252 8208
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17034 8134 17036 8186
rect 17098 8134 17110 8186
rect 17172 8134 17174 8186
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 16956 8112 17252 8132
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17420 7993 17448 8026
rect 17406 7984 17462 7993
rect 17406 7919 17462 7928
rect 17512 7206 17540 9318
rect 17604 9178 17632 9522
rect 18248 9178 18276 9522
rect 19352 9489 19380 17478
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20456 12850 20484 16390
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20168 12640 20220 12646
rect 20168 12582 20220 12588
rect 20180 12374 20208 12582
rect 20456 12442 20484 12786
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20168 12368 20220 12374
rect 20168 12310 20220 12316
rect 19616 12300 19668 12306
rect 19616 12242 19668 12248
rect 19628 11898 19656 12242
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 20548 10554 20576 20198
rect 21270 19816 21326 19825
rect 21270 19751 21326 19760
rect 20956 19612 21252 19632
rect 21012 19610 21036 19612
rect 21092 19610 21116 19612
rect 21172 19610 21196 19612
rect 21034 19558 21036 19610
rect 21098 19558 21110 19610
rect 21172 19558 21174 19610
rect 21012 19556 21036 19558
rect 21092 19556 21116 19558
rect 21172 19556 21196 19558
rect 20956 19536 21252 19556
rect 21284 18834 21312 19751
rect 20812 18828 20864 18834
rect 20812 18770 20864 18776
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 20824 18426 20852 18770
rect 21270 18728 21326 18737
rect 21270 18663 21326 18672
rect 20956 18524 21252 18544
rect 21012 18522 21036 18524
rect 21092 18522 21116 18524
rect 21172 18522 21196 18524
rect 21034 18470 21036 18522
rect 21098 18470 21110 18522
rect 21172 18470 21174 18522
rect 21012 18468 21036 18470
rect 21092 18468 21116 18470
rect 21172 18468 21196 18470
rect 20956 18448 21252 18468
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 21284 17746 21312 18663
rect 21272 17740 21324 17746
rect 21272 17682 21324 17688
rect 20956 17436 21252 17456
rect 21012 17434 21036 17436
rect 21092 17434 21116 17436
rect 21172 17434 21196 17436
rect 21034 17382 21036 17434
rect 21098 17382 21110 17434
rect 21172 17382 21174 17434
rect 21012 17380 21036 17382
rect 21092 17380 21116 17382
rect 21172 17380 21196 17382
rect 20956 17360 21252 17380
rect 21284 17338 21312 17682
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21270 17096 21326 17105
rect 21270 17031 21326 17040
rect 21284 16658 21312 17031
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 20956 16348 21252 16368
rect 21012 16346 21036 16348
rect 21092 16346 21116 16348
rect 21172 16346 21196 16348
rect 21034 16294 21036 16346
rect 21098 16294 21110 16346
rect 21172 16294 21174 16346
rect 21012 16292 21036 16294
rect 21092 16292 21116 16294
rect 21172 16292 21196 16294
rect 20956 16272 21252 16292
rect 21284 16250 21312 16594
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 20956 15260 21252 15280
rect 21012 15258 21036 15260
rect 21092 15258 21116 15260
rect 21172 15258 21196 15260
rect 21034 15206 21036 15258
rect 21098 15206 21110 15258
rect 21172 15206 21174 15258
rect 21012 15204 21036 15206
rect 21092 15204 21116 15206
rect 21172 15204 21196 15206
rect 20956 15184 21252 15204
rect 21454 14240 21510 14249
rect 20956 14172 21252 14192
rect 21454 14175 21510 14184
rect 21012 14170 21036 14172
rect 21092 14170 21116 14172
rect 21172 14170 21196 14172
rect 21034 14118 21036 14170
rect 21098 14118 21110 14170
rect 21172 14118 21174 14170
rect 21012 14116 21036 14118
rect 21092 14116 21116 14118
rect 21172 14116 21196 14118
rect 20956 14096 21252 14116
rect 21468 13394 21496 14175
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20824 12374 20852 13126
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 21468 12986 21496 13330
rect 21456 12980 21508 12986
rect 21456 12922 21508 12928
rect 21088 12708 21140 12714
rect 21088 12650 21140 12656
rect 20812 12368 20864 12374
rect 20812 12310 20864 12316
rect 20824 11898 20852 12310
rect 21100 12238 21128 12650
rect 21732 12368 21784 12374
rect 21732 12310 21784 12316
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 21454 11928 21510 11937
rect 20812 11892 20864 11898
rect 21744 11898 21772 12310
rect 21454 11863 21510 11872
rect 21732 11892 21784 11898
rect 20812 11834 20864 11840
rect 21468 11830 21496 11863
rect 21732 11834 21784 11840
rect 21456 11824 21508 11830
rect 21456 11766 21508 11772
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 20456 10526 20576 10554
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20272 9722 20300 10406
rect 20260 9716 20312 9722
rect 20260 9658 20312 9664
rect 19338 9480 19394 9489
rect 18788 9444 18840 9450
rect 19338 9415 19394 9424
rect 18788 9386 18840 9392
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 16956 7100 17252 7120
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17034 7046 17036 7098
rect 17098 7046 17110 7098
rect 17172 7046 17174 7098
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 16956 7024 17252 7044
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15856 5370 15884 6394
rect 16316 6322 16344 6734
rect 16408 6458 16436 6870
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16580 5840 16632 5846
rect 16580 5782 16632 5788
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 15856 5166 15884 5306
rect 16592 5234 16620 5782
rect 16684 5710 16712 6054
rect 16868 5710 16896 6666
rect 16956 6012 17252 6032
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17034 5958 17036 6010
rect 17098 5958 17110 6010
rect 17172 5958 17174 6010
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 16956 5936 17252 5956
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 16684 4826 16712 5646
rect 16868 5302 16896 5646
rect 16856 5296 16908 5302
rect 16856 5238 16908 5244
rect 16956 4924 17252 4944
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17034 4870 17036 4922
rect 17098 4870 17110 4922
rect 17172 4870 17174 4922
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 16956 4848 17252 4868
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 17512 4690 17540 7142
rect 17972 7002 18000 7346
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 18340 6866 18368 7142
rect 18800 7002 18828 9386
rect 20272 9382 20300 9658
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19352 7002 19380 7278
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 18340 6458 18368 6802
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18800 6322 18828 6938
rect 20364 6458 20392 7142
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16224 4010 16252 4422
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16212 4004 16264 4010
rect 16212 3946 16264 3952
rect 16132 3670 16160 3946
rect 16224 3738 16252 3946
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 15948 3058 15976 3606
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 16224 2990 16252 3674
rect 16500 3602 16528 4082
rect 17512 3942 17540 4626
rect 17880 4214 17908 4626
rect 17868 4208 17920 4214
rect 17868 4150 17920 4156
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 16956 3836 17252 3856
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17034 3782 17036 3834
rect 17098 3782 17110 3834
rect 17172 3782 17174 3834
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 16956 3760 17252 3780
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16500 3126 16528 3538
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 16580 2916 16632 2922
rect 16580 2858 16632 2864
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 16040 2417 16068 2790
rect 16592 2514 16620 2858
rect 16956 2748 17252 2768
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17034 2694 17036 2746
rect 17098 2694 17110 2746
rect 17172 2694 17174 2746
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 16956 2672 17252 2692
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 16026 2408 16082 2417
rect 13268 2372 13320 2378
rect 16026 2343 16082 2352
rect 13268 2314 13320 2320
rect 12956 2204 13252 2224
rect 13012 2202 13036 2204
rect 13092 2202 13116 2204
rect 13172 2202 13196 2204
rect 13034 2150 13036 2202
rect 13098 2150 13110 2202
rect 13172 2150 13174 2202
rect 13012 2148 13036 2150
rect 13092 2148 13116 2150
rect 13172 2148 13196 2150
rect 12956 2128 13252 2148
rect 11886 82 11942 480
rect 11808 54 11942 82
rect 13280 82 13308 2314
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 13542 82 13598 480
rect 13280 54 13598 82
rect 754 0 810 54
rect 2318 0 2374 54
rect 3882 0 3938 54
rect 5538 0 5594 54
rect 7102 0 7158 54
rect 8758 0 8814 54
rect 10322 0 10378 54
rect 11886 0 11942 54
rect 13542 0 13598 54
rect 15106 82 15162 480
rect 15396 82 15424 2246
rect 15106 54 15424 82
rect 16762 82 16818 480
rect 16868 82 16896 2246
rect 17236 2009 17264 2246
rect 17222 2000 17278 2009
rect 17222 1935 17278 1944
rect 17512 1329 17540 3878
rect 17498 1320 17554 1329
rect 17498 1255 17554 1264
rect 16762 54 16896 82
rect 18064 82 18092 6054
rect 18800 5914 18828 6258
rect 20364 6118 20392 6394
rect 20352 6112 20404 6118
rect 20352 6054 20404 6060
rect 20456 5914 20484 10526
rect 20536 10464 20588 10470
rect 20536 10406 20588 10412
rect 20548 9586 20576 10406
rect 20640 10198 20668 10542
rect 20628 10192 20680 10198
rect 20628 10134 20680 10140
rect 21456 10192 21508 10198
rect 21456 10134 21508 10140
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 21468 9722 21496 10134
rect 21836 10062 21864 20198
rect 22190 12880 22246 12889
rect 22190 12815 22246 12824
rect 22100 10600 22152 10606
rect 22098 10568 22100 10577
rect 22152 10568 22154 10577
rect 22098 10503 22154 10512
rect 22112 10470 22140 10503
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 21824 10056 21876 10062
rect 21824 9998 21876 10004
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21456 9716 21508 9722
rect 21456 9658 21508 9664
rect 21560 9586 21588 9930
rect 21836 9722 21864 9998
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 21548 9580 21600 9586
rect 21548 9522 21600 9528
rect 20548 9178 20576 9522
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 21456 9036 21508 9042
rect 21456 8978 21508 8984
rect 21468 8809 21496 8978
rect 21454 8800 21510 8809
rect 20956 8732 21252 8752
rect 21454 8735 21510 8744
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 21468 8634 21496 8735
rect 22204 8634 22232 12815
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 21376 7721 21404 7890
rect 21362 7712 21418 7721
rect 20956 7644 21252 7664
rect 21362 7647 21418 7656
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 21376 7546 21404 7647
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 21284 6934 21312 7278
rect 21272 6928 21324 6934
rect 21272 6870 21324 6876
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 21284 6458 21312 6870
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21376 6390 21404 6598
rect 21364 6384 21416 6390
rect 21364 6326 21416 6332
rect 21468 6322 21496 6734
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 20628 6180 20680 6186
rect 20628 6122 20680 6128
rect 20640 5914 20668 6122
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18156 4758 18184 5102
rect 18800 5098 18828 5850
rect 20180 5234 20208 5850
rect 21272 5840 21324 5846
rect 21272 5782 21324 5788
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 21284 5370 21312 5782
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 20168 5228 20220 5234
rect 20168 5170 20220 5176
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 18788 5092 18840 5098
rect 18788 5034 18840 5040
rect 19892 5024 19944 5030
rect 19892 4966 19944 4972
rect 20074 4992 20130 5001
rect 18144 4752 18196 4758
rect 18144 4694 18196 4700
rect 19904 4078 19932 4966
rect 20074 4927 20130 4936
rect 20088 4690 20116 4927
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 20088 4282 20116 4626
rect 20456 4554 20484 5170
rect 20812 4752 20864 4758
rect 20812 4694 20864 4700
rect 20444 4548 20496 4554
rect 20444 4490 20496 4496
rect 20076 4276 20128 4282
rect 20076 4218 20128 4224
rect 19892 4072 19944 4078
rect 19892 4014 19944 4020
rect 19904 3738 19932 4014
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 20456 3670 20484 4490
rect 20824 4010 20852 4694
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 21284 4282 21312 4558
rect 21272 4276 21324 4282
rect 21272 4218 21324 4224
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 20444 3664 20496 3670
rect 20444 3606 20496 3612
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 19524 2848 19576 2854
rect 19524 2790 19576 2796
rect 18326 82 18382 480
rect 18064 54 18382 82
rect 19536 82 19564 2790
rect 21468 2650 21496 6258
rect 21730 5944 21786 5953
rect 21730 5879 21786 5888
rect 21744 5846 21772 5879
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 21456 2644 21508 2650
rect 21456 2586 21508 2592
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 22836 2304 22888 2310
rect 22836 2246 22888 2252
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 19890 82 19946 480
rect 19536 54 19946 82
rect 21284 82 21312 2246
rect 21546 82 21602 480
rect 21284 54 21602 82
rect 22848 82 22876 2246
rect 23110 82 23166 480
rect 22848 54 23166 82
rect 15106 0 15162 54
rect 16762 0 16818 54
rect 18326 0 18382 54
rect 19890 0 19946 54
rect 21546 0 21602 54
rect 23110 0 23166 54
<< via2 >>
rect 1214 21528 1270 21584
rect 5814 22752 5870 22808
rect 4956 21786 5012 21788
rect 5036 21786 5092 21788
rect 5116 21786 5172 21788
rect 5196 21786 5252 21788
rect 4956 21734 4982 21786
rect 4982 21734 5012 21786
rect 5036 21734 5046 21786
rect 5046 21734 5092 21786
rect 5116 21734 5162 21786
rect 5162 21734 5172 21786
rect 5196 21734 5226 21786
rect 5226 21734 5252 21786
rect 4956 21732 5012 21734
rect 5036 21732 5092 21734
rect 5116 21732 5172 21734
rect 5196 21732 5252 21734
rect 4956 20698 5012 20700
rect 5036 20698 5092 20700
rect 5116 20698 5172 20700
rect 5196 20698 5252 20700
rect 4956 20646 4982 20698
rect 4982 20646 5012 20698
rect 5036 20646 5046 20698
rect 5046 20646 5092 20698
rect 5116 20646 5162 20698
rect 5162 20646 5172 20698
rect 5196 20646 5226 20698
rect 5226 20646 5252 20698
rect 4956 20644 5012 20646
rect 5036 20644 5092 20646
rect 5116 20644 5172 20646
rect 5196 20644 5252 20646
rect 1306 20304 1362 20360
rect 1214 19080 1270 19136
rect 1490 17992 1546 18048
rect 110 17312 166 17368
rect 1582 16360 1638 16416
rect 1950 15408 2006 15464
rect 4956 19610 5012 19612
rect 5036 19610 5092 19612
rect 5116 19610 5172 19612
rect 5196 19610 5252 19612
rect 4956 19558 4982 19610
rect 4982 19558 5012 19610
rect 5036 19558 5046 19610
rect 5046 19558 5092 19610
rect 5116 19558 5162 19610
rect 5162 19558 5172 19610
rect 5196 19558 5226 19610
rect 5226 19558 5252 19610
rect 4956 19556 5012 19558
rect 5036 19556 5092 19558
rect 5116 19556 5172 19558
rect 5196 19556 5252 19558
rect 4956 18522 5012 18524
rect 5036 18522 5092 18524
rect 5116 18522 5172 18524
rect 5196 18522 5252 18524
rect 4956 18470 4982 18522
rect 4982 18470 5012 18522
rect 5036 18470 5046 18522
rect 5046 18470 5092 18522
rect 5116 18470 5162 18522
rect 5162 18470 5172 18522
rect 5196 18470 5226 18522
rect 5226 18470 5252 18522
rect 4956 18468 5012 18470
rect 5036 18468 5092 18470
rect 5116 18468 5172 18470
rect 5196 18468 5252 18470
rect 4956 17434 5012 17436
rect 5036 17434 5092 17436
rect 5116 17434 5172 17436
rect 5196 17434 5252 17436
rect 4956 17382 4982 17434
rect 4982 17382 5012 17434
rect 5036 17382 5046 17434
rect 5046 17382 5092 17434
rect 5116 17382 5162 17434
rect 5162 17382 5172 17434
rect 5196 17382 5226 17434
rect 5226 17382 5252 17434
rect 4956 17380 5012 17382
rect 5036 17380 5092 17382
rect 5116 17380 5172 17382
rect 5196 17380 5252 17382
rect 4956 16346 5012 16348
rect 5036 16346 5092 16348
rect 5116 16346 5172 16348
rect 5196 16346 5252 16348
rect 4956 16294 4982 16346
rect 4982 16294 5012 16346
rect 5036 16294 5046 16346
rect 5046 16294 5092 16346
rect 5116 16294 5162 16346
rect 5162 16294 5172 16346
rect 5196 16294 5226 16346
rect 5226 16294 5252 16346
rect 4956 16292 5012 16294
rect 5036 16292 5092 16294
rect 5116 16292 5172 16294
rect 5196 16292 5252 16294
rect 2042 15000 2098 15056
rect 1122 12008 1178 12064
rect 18 10104 74 10160
rect 110 8880 166 8936
rect 110 7656 166 7712
rect 110 6568 166 6624
rect 110 5344 166 5400
rect 110 4086 166 4142
rect 110 2896 166 2952
rect 4956 15258 5012 15260
rect 5036 15258 5092 15260
rect 5116 15258 5172 15260
rect 5196 15258 5252 15260
rect 4956 15206 4982 15258
rect 4982 15206 5012 15258
rect 5036 15206 5046 15258
rect 5046 15206 5092 15258
rect 5116 15206 5162 15258
rect 5162 15206 5172 15258
rect 5196 15206 5226 15258
rect 5226 15206 5252 15258
rect 4956 15204 5012 15206
rect 5036 15204 5092 15206
rect 5116 15204 5172 15206
rect 5196 15204 5252 15206
rect 3422 9424 3478 9480
rect 2318 2896 2374 2952
rect 1858 2216 1914 2272
rect 4956 14170 5012 14172
rect 5036 14170 5092 14172
rect 5116 14170 5172 14172
rect 5196 14170 5252 14172
rect 4956 14118 4982 14170
rect 4982 14118 5012 14170
rect 5036 14118 5046 14170
rect 5046 14118 5092 14170
rect 5116 14118 5162 14170
rect 5162 14118 5172 14170
rect 5196 14118 5226 14170
rect 5226 14118 5252 14170
rect 4956 14116 5012 14118
rect 5036 14116 5092 14118
rect 5116 14116 5172 14118
rect 5196 14116 5252 14118
rect 4956 13082 5012 13084
rect 5036 13082 5092 13084
rect 5116 13082 5172 13084
rect 5196 13082 5252 13084
rect 4956 13030 4982 13082
rect 4982 13030 5012 13082
rect 5036 13030 5046 13082
rect 5046 13030 5092 13082
rect 5116 13030 5162 13082
rect 5162 13030 5172 13082
rect 5196 13030 5226 13082
rect 5226 13030 5252 13082
rect 4956 13028 5012 13030
rect 5036 13028 5092 13030
rect 5116 13028 5172 13030
rect 5196 13028 5252 13030
rect 7378 13232 7434 13288
rect 4956 11994 5012 11996
rect 5036 11994 5092 11996
rect 5116 11994 5172 11996
rect 5196 11994 5252 11996
rect 4956 11942 4982 11994
rect 4982 11942 5012 11994
rect 5036 11942 5046 11994
rect 5046 11942 5092 11994
rect 5116 11942 5162 11994
rect 5162 11942 5172 11994
rect 5196 11942 5226 11994
rect 5226 11942 5252 11994
rect 4956 11940 5012 11942
rect 5036 11940 5092 11942
rect 5116 11940 5172 11942
rect 5196 11940 5252 11942
rect 4956 10906 5012 10908
rect 5036 10906 5092 10908
rect 5116 10906 5172 10908
rect 5196 10906 5252 10908
rect 4956 10854 4982 10906
rect 4982 10854 5012 10906
rect 5036 10854 5046 10906
rect 5046 10854 5092 10906
rect 5116 10854 5162 10906
rect 5162 10854 5172 10906
rect 5196 10854 5226 10906
rect 5226 10854 5252 10906
rect 4956 10852 5012 10854
rect 5036 10852 5092 10854
rect 5116 10852 5172 10854
rect 5196 10852 5252 10854
rect 4956 9818 5012 9820
rect 5036 9818 5092 9820
rect 5116 9818 5172 9820
rect 5196 9818 5252 9820
rect 4956 9766 4982 9818
rect 4982 9766 5012 9818
rect 5036 9766 5046 9818
rect 5046 9766 5092 9818
rect 5116 9766 5162 9818
rect 5162 9766 5172 9818
rect 5196 9766 5226 9818
rect 5226 9766 5252 9818
rect 4956 9764 5012 9766
rect 5036 9764 5092 9766
rect 5116 9764 5172 9766
rect 5196 9764 5252 9766
rect 4956 8730 5012 8732
rect 5036 8730 5092 8732
rect 5116 8730 5172 8732
rect 5196 8730 5252 8732
rect 4956 8678 4982 8730
rect 4982 8678 5012 8730
rect 5036 8678 5046 8730
rect 5046 8678 5092 8730
rect 5116 8678 5162 8730
rect 5162 8678 5172 8730
rect 5196 8678 5226 8730
rect 5226 8678 5252 8730
rect 4956 8676 5012 8678
rect 5036 8676 5092 8678
rect 5116 8676 5172 8678
rect 5196 8676 5252 8678
rect 4956 7642 5012 7644
rect 5036 7642 5092 7644
rect 5116 7642 5172 7644
rect 5196 7642 5252 7644
rect 4956 7590 4982 7642
rect 4982 7590 5012 7642
rect 5036 7590 5046 7642
rect 5046 7590 5092 7642
rect 5116 7590 5162 7642
rect 5162 7590 5172 7642
rect 5196 7590 5226 7642
rect 5226 7590 5252 7642
rect 4956 7588 5012 7590
rect 5036 7588 5092 7590
rect 5116 7588 5172 7590
rect 5196 7588 5252 7590
rect 5814 11056 5870 11112
rect 4956 6554 5012 6556
rect 5036 6554 5092 6556
rect 5116 6554 5172 6556
rect 5196 6554 5252 6556
rect 4956 6502 4982 6554
rect 4982 6502 5012 6554
rect 5036 6502 5046 6554
rect 5046 6502 5092 6554
rect 5116 6502 5162 6554
rect 5162 6502 5172 6554
rect 5196 6502 5226 6554
rect 5226 6502 5252 6554
rect 4956 6500 5012 6502
rect 5036 6500 5092 6502
rect 5116 6500 5172 6502
rect 5196 6500 5252 6502
rect 4956 5466 5012 5468
rect 5036 5466 5092 5468
rect 5116 5466 5172 5468
rect 5196 5466 5252 5468
rect 4956 5414 4982 5466
rect 4982 5414 5012 5466
rect 5036 5414 5046 5466
rect 5046 5414 5092 5466
rect 5116 5414 5162 5466
rect 5162 5414 5172 5466
rect 5196 5414 5226 5466
rect 5226 5414 5252 5466
rect 4956 5412 5012 5414
rect 5036 5412 5092 5414
rect 5116 5412 5172 5414
rect 5196 5412 5252 5414
rect 4956 4378 5012 4380
rect 5036 4378 5092 4380
rect 5116 4378 5172 4380
rect 5196 4378 5252 4380
rect 4956 4326 4982 4378
rect 4982 4326 5012 4378
rect 5036 4326 5046 4378
rect 5046 4326 5092 4378
rect 5116 4326 5162 4378
rect 5162 4326 5172 4378
rect 5196 4326 5226 4378
rect 5226 4326 5252 4378
rect 4956 4324 5012 4326
rect 5036 4324 5092 4326
rect 5116 4324 5172 4326
rect 5196 4324 5252 4326
rect 4956 3290 5012 3292
rect 5036 3290 5092 3292
rect 5116 3290 5172 3292
rect 5196 3290 5252 3292
rect 4956 3238 4982 3290
rect 4982 3238 5012 3290
rect 5036 3238 5046 3290
rect 5046 3238 5092 3290
rect 5116 3238 5162 3290
rect 5162 3238 5172 3290
rect 5196 3238 5226 3290
rect 5226 3238 5252 3290
rect 4956 3236 5012 3238
rect 5036 3236 5092 3238
rect 5116 3236 5172 3238
rect 5196 3236 5252 3238
rect 4526 2352 4582 2408
rect 4956 2202 5012 2204
rect 5036 2202 5092 2204
rect 5116 2202 5172 2204
rect 5196 2202 5252 2204
rect 4956 2150 4982 2202
rect 4982 2150 5012 2202
rect 5036 2150 5046 2202
rect 5046 2150 5092 2202
rect 5116 2150 5162 2202
rect 5162 2150 5172 2202
rect 5196 2150 5226 2202
rect 5226 2150 5252 2202
rect 4956 2148 5012 2150
rect 5036 2148 5092 2150
rect 5116 2148 5172 2150
rect 5196 2148 5252 2150
rect 6734 1128 6790 1184
rect 8114 8880 8170 8936
rect 8956 21242 9012 21244
rect 9036 21242 9092 21244
rect 9116 21242 9172 21244
rect 9196 21242 9252 21244
rect 8956 21190 8982 21242
rect 8982 21190 9012 21242
rect 9036 21190 9046 21242
rect 9046 21190 9092 21242
rect 9116 21190 9162 21242
rect 9162 21190 9172 21242
rect 9196 21190 9226 21242
rect 9226 21190 9252 21242
rect 8956 21188 9012 21190
rect 9036 21188 9092 21190
rect 9116 21188 9172 21190
rect 9196 21188 9252 21190
rect 8956 20154 9012 20156
rect 9036 20154 9092 20156
rect 9116 20154 9172 20156
rect 9196 20154 9252 20156
rect 8956 20102 8982 20154
rect 8982 20102 9012 20154
rect 9036 20102 9046 20154
rect 9046 20102 9092 20154
rect 9116 20102 9162 20154
rect 9162 20102 9172 20154
rect 9196 20102 9226 20154
rect 9226 20102 9252 20154
rect 8956 20100 9012 20102
rect 9036 20100 9092 20102
rect 9116 20100 9172 20102
rect 9196 20100 9252 20102
rect 8956 19066 9012 19068
rect 9036 19066 9092 19068
rect 9116 19066 9172 19068
rect 9196 19066 9252 19068
rect 8956 19014 8982 19066
rect 8982 19014 9012 19066
rect 9036 19014 9046 19066
rect 9046 19014 9092 19066
rect 9116 19014 9162 19066
rect 9162 19014 9172 19066
rect 9196 19014 9226 19066
rect 9226 19014 9252 19066
rect 8956 19012 9012 19014
rect 9036 19012 9092 19014
rect 9116 19012 9172 19014
rect 9196 19012 9252 19014
rect 8390 17720 8446 17776
rect 8956 17978 9012 17980
rect 9036 17978 9092 17980
rect 9116 17978 9172 17980
rect 9196 17978 9252 17980
rect 8956 17926 8982 17978
rect 8982 17926 9012 17978
rect 9036 17926 9046 17978
rect 9046 17926 9092 17978
rect 9116 17926 9162 17978
rect 9162 17926 9172 17978
rect 9196 17926 9226 17978
rect 9226 17926 9252 17978
rect 8956 17924 9012 17926
rect 9036 17924 9092 17926
rect 9116 17924 9172 17926
rect 9196 17924 9252 17926
rect 7746 2488 7802 2544
rect 8956 16890 9012 16892
rect 9036 16890 9092 16892
rect 9116 16890 9172 16892
rect 9196 16890 9252 16892
rect 8956 16838 8982 16890
rect 8982 16838 9012 16890
rect 9036 16838 9046 16890
rect 9046 16838 9092 16890
rect 9116 16838 9162 16890
rect 9162 16838 9172 16890
rect 9196 16838 9226 16890
rect 9226 16838 9252 16890
rect 8956 16836 9012 16838
rect 9036 16836 9092 16838
rect 9116 16836 9172 16838
rect 9196 16836 9252 16838
rect 8956 15802 9012 15804
rect 9036 15802 9092 15804
rect 9116 15802 9172 15804
rect 9196 15802 9252 15804
rect 8956 15750 8982 15802
rect 8982 15750 9012 15802
rect 9036 15750 9046 15802
rect 9046 15750 9092 15802
rect 9116 15750 9162 15802
rect 9162 15750 9172 15802
rect 9196 15750 9226 15802
rect 9226 15750 9252 15802
rect 8956 15748 9012 15750
rect 9036 15748 9092 15750
rect 9116 15748 9172 15750
rect 9196 15748 9252 15750
rect 8942 15000 8998 15056
rect 8956 14714 9012 14716
rect 9036 14714 9092 14716
rect 9116 14714 9172 14716
rect 9196 14714 9252 14716
rect 8956 14662 8982 14714
rect 8982 14662 9012 14714
rect 9036 14662 9046 14714
rect 9046 14662 9092 14714
rect 9116 14662 9162 14714
rect 9162 14662 9172 14714
rect 9196 14662 9226 14714
rect 9226 14662 9252 14714
rect 8956 14660 9012 14662
rect 9036 14660 9092 14662
rect 9116 14660 9172 14662
rect 9196 14660 9252 14662
rect 9402 13776 9458 13832
rect 9678 13776 9734 13832
rect 8956 13626 9012 13628
rect 9036 13626 9092 13628
rect 9116 13626 9172 13628
rect 9196 13626 9252 13628
rect 8956 13574 8982 13626
rect 8982 13574 9012 13626
rect 9036 13574 9046 13626
rect 9046 13574 9092 13626
rect 9116 13574 9162 13626
rect 9162 13574 9172 13626
rect 9196 13574 9226 13626
rect 9226 13574 9252 13626
rect 8956 13572 9012 13574
rect 9036 13572 9092 13574
rect 9116 13572 9172 13574
rect 9196 13572 9252 13574
rect 8956 12538 9012 12540
rect 9036 12538 9092 12540
rect 9116 12538 9172 12540
rect 9196 12538 9252 12540
rect 8956 12486 8982 12538
rect 8982 12486 9012 12538
rect 9036 12486 9046 12538
rect 9046 12486 9092 12538
rect 9116 12486 9162 12538
rect 9162 12486 9172 12538
rect 9196 12486 9226 12538
rect 9226 12486 9252 12538
rect 8956 12484 9012 12486
rect 9036 12484 9092 12486
rect 9116 12484 9172 12486
rect 9196 12484 9252 12486
rect 8956 11450 9012 11452
rect 9036 11450 9092 11452
rect 9116 11450 9172 11452
rect 9196 11450 9252 11452
rect 8956 11398 8982 11450
rect 8982 11398 9012 11450
rect 9036 11398 9046 11450
rect 9046 11398 9092 11450
rect 9116 11398 9162 11450
rect 9162 11398 9172 11450
rect 9196 11398 9226 11450
rect 9226 11398 9252 11450
rect 8956 11396 9012 11398
rect 9036 11396 9092 11398
rect 9116 11396 9172 11398
rect 9196 11396 9252 11398
rect 8956 10362 9012 10364
rect 9036 10362 9092 10364
rect 9116 10362 9172 10364
rect 9196 10362 9252 10364
rect 8956 10310 8982 10362
rect 8982 10310 9012 10362
rect 9036 10310 9046 10362
rect 9046 10310 9092 10362
rect 9116 10310 9162 10362
rect 9162 10310 9172 10362
rect 9196 10310 9226 10362
rect 9226 10310 9252 10362
rect 8956 10308 9012 10310
rect 9036 10308 9092 10310
rect 9116 10308 9172 10310
rect 9196 10308 9252 10310
rect 8956 9274 9012 9276
rect 9036 9274 9092 9276
rect 9116 9274 9172 9276
rect 9196 9274 9252 9276
rect 8956 9222 8982 9274
rect 8982 9222 9012 9274
rect 9036 9222 9046 9274
rect 9046 9222 9092 9274
rect 9116 9222 9162 9274
rect 9162 9222 9172 9274
rect 9196 9222 9226 9274
rect 9226 9222 9252 9274
rect 8956 9220 9012 9222
rect 9036 9220 9092 9222
rect 9116 9220 9172 9222
rect 9196 9220 9252 9222
rect 12956 21786 13012 21788
rect 13036 21786 13092 21788
rect 13116 21786 13172 21788
rect 13196 21786 13252 21788
rect 12956 21734 12982 21786
rect 12982 21734 13012 21786
rect 13036 21734 13046 21786
rect 13046 21734 13092 21786
rect 13116 21734 13162 21786
rect 13162 21734 13172 21786
rect 13196 21734 13226 21786
rect 13226 21734 13252 21786
rect 12956 21732 13012 21734
rect 13036 21732 13092 21734
rect 13116 21732 13172 21734
rect 13196 21732 13252 21734
rect 12956 20698 13012 20700
rect 13036 20698 13092 20700
rect 13116 20698 13172 20700
rect 13196 20698 13252 20700
rect 12956 20646 12982 20698
rect 12982 20646 13012 20698
rect 13036 20646 13046 20698
rect 13046 20646 13092 20698
rect 13116 20646 13162 20698
rect 13162 20646 13172 20698
rect 13196 20646 13226 20698
rect 13226 20646 13252 20698
rect 12956 20644 13012 20646
rect 13036 20644 13092 20646
rect 13116 20644 13172 20646
rect 13196 20644 13252 20646
rect 8956 8186 9012 8188
rect 9036 8186 9092 8188
rect 9116 8186 9172 8188
rect 9196 8186 9252 8188
rect 8956 8134 8982 8186
rect 8982 8134 9012 8186
rect 9036 8134 9046 8186
rect 9046 8134 9092 8186
rect 9116 8134 9162 8186
rect 9162 8134 9172 8186
rect 9196 8134 9226 8186
rect 9226 8134 9252 8186
rect 8956 8132 9012 8134
rect 9036 8132 9092 8134
rect 9116 8132 9172 8134
rect 9196 8132 9252 8134
rect 8956 7098 9012 7100
rect 9036 7098 9092 7100
rect 9116 7098 9172 7100
rect 9196 7098 9252 7100
rect 8956 7046 8982 7098
rect 8982 7046 9012 7098
rect 9036 7046 9046 7098
rect 9046 7046 9092 7098
rect 9116 7046 9162 7098
rect 9162 7046 9172 7098
rect 9196 7046 9226 7098
rect 9226 7046 9252 7098
rect 8956 7044 9012 7046
rect 9036 7044 9092 7046
rect 9116 7044 9172 7046
rect 9196 7044 9252 7046
rect 8956 6010 9012 6012
rect 9036 6010 9092 6012
rect 9116 6010 9172 6012
rect 9196 6010 9252 6012
rect 8956 5958 8982 6010
rect 8982 5958 9012 6010
rect 9036 5958 9046 6010
rect 9046 5958 9092 6010
rect 9116 5958 9162 6010
rect 9162 5958 9172 6010
rect 9196 5958 9226 6010
rect 9226 5958 9252 6010
rect 8956 5956 9012 5958
rect 9036 5956 9092 5958
rect 9116 5956 9172 5958
rect 9196 5956 9252 5958
rect 8956 4922 9012 4924
rect 9036 4922 9092 4924
rect 9116 4922 9172 4924
rect 9196 4922 9252 4924
rect 8956 4870 8982 4922
rect 8982 4870 9012 4922
rect 9036 4870 9046 4922
rect 9046 4870 9092 4922
rect 9116 4870 9162 4922
rect 9162 4870 9172 4922
rect 9196 4870 9226 4922
rect 9226 4870 9252 4922
rect 8956 4868 9012 4870
rect 9036 4868 9092 4870
rect 9116 4868 9172 4870
rect 9196 4868 9252 4870
rect 8956 3834 9012 3836
rect 9036 3834 9092 3836
rect 9116 3834 9172 3836
rect 9196 3834 9252 3836
rect 8956 3782 8982 3834
rect 8982 3782 9012 3834
rect 9036 3782 9046 3834
rect 9046 3782 9092 3834
rect 9116 3782 9162 3834
rect 9162 3782 9172 3834
rect 9196 3782 9226 3834
rect 9226 3782 9252 3834
rect 8956 3780 9012 3782
rect 9036 3780 9092 3782
rect 9116 3780 9172 3782
rect 9196 3780 9252 3782
rect 8956 2746 9012 2748
rect 9036 2746 9092 2748
rect 9116 2746 9172 2748
rect 9196 2746 9252 2748
rect 8956 2694 8982 2746
rect 8982 2694 9012 2746
rect 9036 2694 9046 2746
rect 9046 2694 9092 2746
rect 9116 2694 9162 2746
rect 9162 2694 9172 2746
rect 9196 2694 9226 2746
rect 9226 2694 9252 2746
rect 8956 2692 9012 2694
rect 9036 2692 9092 2694
rect 9116 2692 9172 2694
rect 9196 2692 9252 2694
rect 12956 19610 13012 19612
rect 13036 19610 13092 19612
rect 13116 19610 13172 19612
rect 13196 19610 13252 19612
rect 12956 19558 12982 19610
rect 12982 19558 13012 19610
rect 13036 19558 13046 19610
rect 13046 19558 13092 19610
rect 13116 19558 13162 19610
rect 13162 19558 13172 19610
rect 13196 19558 13226 19610
rect 13226 19558 13252 19610
rect 12956 19556 13012 19558
rect 13036 19556 13092 19558
rect 13116 19556 13172 19558
rect 13196 19556 13252 19558
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 16982 21242
rect 16982 21190 17012 21242
rect 17036 21190 17046 21242
rect 17046 21190 17092 21242
rect 17116 21190 17162 21242
rect 17162 21190 17172 21242
rect 17196 21190 17226 21242
rect 17226 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 12956 18522 13012 18524
rect 13036 18522 13092 18524
rect 13116 18522 13172 18524
rect 13196 18522 13252 18524
rect 12956 18470 12982 18522
rect 12982 18470 13012 18522
rect 13036 18470 13046 18522
rect 13046 18470 13092 18522
rect 13116 18470 13162 18522
rect 13162 18470 13172 18522
rect 13196 18470 13226 18522
rect 13226 18470 13252 18522
rect 12956 18468 13012 18470
rect 13036 18468 13092 18470
rect 13116 18468 13172 18470
rect 13196 18468 13252 18470
rect 12956 17434 13012 17436
rect 13036 17434 13092 17436
rect 13116 17434 13172 17436
rect 13196 17434 13252 17436
rect 12956 17382 12982 17434
rect 12982 17382 13012 17434
rect 13036 17382 13046 17434
rect 13046 17382 13092 17434
rect 13116 17382 13162 17434
rect 13162 17382 13172 17434
rect 13196 17382 13226 17434
rect 13226 17382 13252 17434
rect 12956 17380 13012 17382
rect 13036 17380 13092 17382
rect 13116 17380 13172 17382
rect 13196 17380 13252 17382
rect 10322 7928 10378 7984
rect 12956 16346 13012 16348
rect 13036 16346 13092 16348
rect 13116 16346 13172 16348
rect 13196 16346 13252 16348
rect 12956 16294 12982 16346
rect 12982 16294 13012 16346
rect 13036 16294 13046 16346
rect 13046 16294 13092 16346
rect 13116 16294 13162 16346
rect 13162 16294 13172 16346
rect 13196 16294 13226 16346
rect 13226 16294 13252 16346
rect 12956 16292 13012 16294
rect 13036 16292 13092 16294
rect 13116 16292 13172 16294
rect 13196 16292 13252 16294
rect 16026 17720 16082 17776
rect 12956 15258 13012 15260
rect 13036 15258 13092 15260
rect 13116 15258 13172 15260
rect 13196 15258 13252 15260
rect 12956 15206 12982 15258
rect 12982 15206 13012 15258
rect 13036 15206 13046 15258
rect 13046 15206 13092 15258
rect 13116 15206 13162 15258
rect 13162 15206 13172 15258
rect 13196 15206 13226 15258
rect 13226 15206 13252 15258
rect 12956 15204 13012 15206
rect 13036 15204 13092 15206
rect 13116 15204 13172 15206
rect 13196 15204 13252 15206
rect 14554 15544 14610 15600
rect 12956 14170 13012 14172
rect 13036 14170 13092 14172
rect 13116 14170 13172 14172
rect 13196 14170 13252 14172
rect 12956 14118 12982 14170
rect 12982 14118 13012 14170
rect 13036 14118 13046 14170
rect 13046 14118 13092 14170
rect 13116 14118 13162 14170
rect 13162 14118 13172 14170
rect 13196 14118 13226 14170
rect 13226 14118 13252 14170
rect 12956 14116 13012 14118
rect 13036 14116 13092 14118
rect 13116 14116 13172 14118
rect 13196 14116 13252 14118
rect 12956 13082 13012 13084
rect 13036 13082 13092 13084
rect 13116 13082 13172 13084
rect 13196 13082 13252 13084
rect 12956 13030 12982 13082
rect 12982 13030 13012 13082
rect 13036 13030 13046 13082
rect 13046 13030 13092 13082
rect 13116 13030 13162 13082
rect 13162 13030 13172 13082
rect 13196 13030 13226 13082
rect 13226 13030 13252 13082
rect 12956 13028 13012 13030
rect 13036 13028 13092 13030
rect 13116 13028 13172 13030
rect 13196 13028 13252 13030
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 16982 20154
rect 16982 20102 17012 20154
rect 17036 20102 17046 20154
rect 17046 20102 17092 20154
rect 17116 20102 17162 20154
rect 17162 20102 17172 20154
rect 17196 20102 17226 20154
rect 17226 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 16982 19066
rect 16982 19014 17012 19066
rect 17036 19014 17046 19066
rect 17046 19014 17092 19066
rect 17116 19014 17162 19066
rect 17162 19014 17172 19066
rect 17196 19014 17226 19066
rect 17226 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 16982 17978
rect 16982 17926 17012 17978
rect 17036 17926 17046 17978
rect 17046 17926 17092 17978
rect 17116 17926 17162 17978
rect 17162 17926 17172 17978
rect 17196 17926 17226 17978
rect 17226 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 21638 22616 21694 22672
rect 20956 21786 21012 21788
rect 21036 21786 21092 21788
rect 21116 21786 21172 21788
rect 21196 21786 21252 21788
rect 20956 21734 20982 21786
rect 20982 21734 21012 21786
rect 21036 21734 21046 21786
rect 21046 21734 21092 21786
rect 21116 21734 21162 21786
rect 21162 21734 21172 21786
rect 21196 21734 21226 21786
rect 21226 21734 21252 21786
rect 20956 21732 21012 21734
rect 21036 21732 21092 21734
rect 21116 21732 21172 21734
rect 21196 21732 21252 21734
rect 20956 20698 21012 20700
rect 21036 20698 21092 20700
rect 21116 20698 21172 20700
rect 21196 20698 21252 20700
rect 20956 20646 20982 20698
rect 20982 20646 21012 20698
rect 21036 20646 21046 20698
rect 21046 20646 21092 20698
rect 21116 20646 21162 20698
rect 21162 20646 21172 20698
rect 21196 20646 21226 20698
rect 21226 20646 21252 20698
rect 20956 20644 21012 20646
rect 21036 20644 21092 20646
rect 21116 20644 21172 20646
rect 21196 20644 21252 20646
rect 23570 21800 23626 21856
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 16982 16890
rect 16982 16838 17012 16890
rect 17036 16838 17046 16890
rect 17046 16838 17092 16890
rect 17116 16838 17162 16890
rect 17162 16838 17172 16890
rect 17196 16838 17226 16890
rect 17226 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 16982 15802
rect 16982 15750 17012 15802
rect 17036 15750 17046 15802
rect 17046 15750 17092 15802
rect 17116 15750 17162 15802
rect 17162 15750 17172 15802
rect 17196 15750 17226 15802
rect 17226 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 16982 14714
rect 16982 14662 17012 14714
rect 17036 14662 17046 14714
rect 17046 14662 17092 14714
rect 17116 14662 17162 14714
rect 17162 14662 17172 14714
rect 17196 14662 17226 14714
rect 17226 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 16982 13626
rect 16982 13574 17012 13626
rect 17036 13574 17046 13626
rect 17046 13574 17092 13626
rect 17116 13574 17162 13626
rect 17162 13574 17172 13626
rect 17196 13574 17226 13626
rect 17226 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 12956 11994 13012 11996
rect 13036 11994 13092 11996
rect 13116 11994 13172 11996
rect 13196 11994 13252 11996
rect 12956 11942 12982 11994
rect 12982 11942 13012 11994
rect 13036 11942 13046 11994
rect 13046 11942 13092 11994
rect 13116 11942 13162 11994
rect 13162 11942 13172 11994
rect 13196 11942 13226 11994
rect 13226 11942 13252 11994
rect 12956 11940 13012 11942
rect 13036 11940 13092 11942
rect 13116 11940 13172 11942
rect 13196 11940 13252 11942
rect 12956 10906 13012 10908
rect 13036 10906 13092 10908
rect 13116 10906 13172 10908
rect 13196 10906 13252 10908
rect 12956 10854 12982 10906
rect 12982 10854 13012 10906
rect 13036 10854 13046 10906
rect 13046 10854 13092 10906
rect 13116 10854 13162 10906
rect 13162 10854 13172 10906
rect 13196 10854 13226 10906
rect 13226 10854 13252 10906
rect 12956 10852 13012 10854
rect 13036 10852 13092 10854
rect 13116 10852 13172 10854
rect 13196 10852 13252 10854
rect 12956 9818 13012 9820
rect 13036 9818 13092 9820
rect 13116 9818 13172 9820
rect 13196 9818 13252 9820
rect 12956 9766 12982 9818
rect 12982 9766 13012 9818
rect 13036 9766 13046 9818
rect 13046 9766 13092 9818
rect 13116 9766 13162 9818
rect 13162 9766 13172 9818
rect 13196 9766 13226 9818
rect 13226 9766 13252 9818
rect 12956 9764 13012 9766
rect 13036 9764 13092 9766
rect 13116 9764 13172 9766
rect 13196 9764 13252 9766
rect 12956 8730 13012 8732
rect 13036 8730 13092 8732
rect 13116 8730 13172 8732
rect 13196 8730 13252 8732
rect 12956 8678 12982 8730
rect 12982 8678 13012 8730
rect 13036 8678 13046 8730
rect 13046 8678 13092 8730
rect 13116 8678 13162 8730
rect 13162 8678 13172 8730
rect 13196 8678 13226 8730
rect 13226 8678 13252 8730
rect 12956 8676 13012 8678
rect 13036 8676 13092 8678
rect 13116 8676 13172 8678
rect 13196 8676 13252 8678
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 16982 12538
rect 16982 12486 17012 12538
rect 17036 12486 17046 12538
rect 17046 12486 17092 12538
rect 17116 12486 17162 12538
rect 17162 12486 17172 12538
rect 17196 12486 17226 12538
rect 17226 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 16982 11450
rect 16982 11398 17012 11450
rect 17036 11398 17046 11450
rect 17046 11398 17092 11450
rect 17116 11398 17162 11450
rect 17162 11398 17172 11450
rect 17196 11398 17226 11450
rect 17226 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 16982 10362
rect 16982 10310 17012 10362
rect 17036 10310 17046 10362
rect 17046 10310 17092 10362
rect 17116 10310 17162 10362
rect 17162 10310 17172 10362
rect 17196 10310 17226 10362
rect 17226 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 12956 7642 13012 7644
rect 13036 7642 13092 7644
rect 13116 7642 13172 7644
rect 13196 7642 13252 7644
rect 12956 7590 12982 7642
rect 12982 7590 13012 7642
rect 13036 7590 13046 7642
rect 13046 7590 13092 7642
rect 13116 7590 13162 7642
rect 13162 7590 13172 7642
rect 13196 7590 13226 7642
rect 13226 7590 13252 7642
rect 12956 7588 13012 7590
rect 13036 7588 13092 7590
rect 13116 7588 13172 7590
rect 13196 7588 13252 7590
rect 12956 6554 13012 6556
rect 13036 6554 13092 6556
rect 13116 6554 13172 6556
rect 13196 6554 13252 6556
rect 12956 6502 12982 6554
rect 12982 6502 13012 6554
rect 13036 6502 13046 6554
rect 13046 6502 13092 6554
rect 13116 6502 13162 6554
rect 13162 6502 13172 6554
rect 13196 6502 13226 6554
rect 13226 6502 13252 6554
rect 12956 6500 13012 6502
rect 13036 6500 13092 6502
rect 13116 6500 13172 6502
rect 13196 6500 13252 6502
rect 12956 5466 13012 5468
rect 13036 5466 13092 5468
rect 13116 5466 13172 5468
rect 13196 5466 13252 5468
rect 12956 5414 12982 5466
rect 12982 5414 13012 5466
rect 13036 5414 13046 5466
rect 13046 5414 13092 5466
rect 13116 5414 13162 5466
rect 13162 5414 13172 5466
rect 13196 5414 13226 5466
rect 13226 5414 13252 5466
rect 12956 5412 13012 5414
rect 13036 5412 13092 5414
rect 13116 5412 13172 5414
rect 13196 5412 13252 5414
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 16982 9274
rect 16982 9222 17012 9274
rect 17036 9222 17046 9274
rect 17046 9222 17092 9274
rect 17116 9222 17162 9274
rect 17162 9222 17172 9274
rect 17196 9222 17226 9274
rect 17226 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 17130 8880 17186 8936
rect 12956 4378 13012 4380
rect 13036 4378 13092 4380
rect 13116 4378 13172 4380
rect 13196 4378 13252 4380
rect 12956 4326 12982 4378
rect 12982 4326 13012 4378
rect 13036 4326 13046 4378
rect 13046 4326 13092 4378
rect 13116 4326 13162 4378
rect 13162 4326 13172 4378
rect 13196 4326 13226 4378
rect 13226 4326 13252 4378
rect 12956 4324 13012 4326
rect 13036 4324 13092 4326
rect 13116 4324 13172 4326
rect 13196 4324 13252 4326
rect 11794 3440 11850 3496
rect 8758 1944 8814 2000
rect 12956 3290 13012 3292
rect 13036 3290 13092 3292
rect 13116 3290 13172 3292
rect 13196 3290 13252 3292
rect 12956 3238 12982 3290
rect 12982 3238 13012 3290
rect 13036 3238 13046 3290
rect 13046 3238 13092 3290
rect 13116 3238 13162 3290
rect 13162 3238 13172 3290
rect 13196 3238 13226 3290
rect 13226 3238 13252 3290
rect 12956 3236 13012 3238
rect 13036 3236 13092 3238
rect 13116 3236 13172 3238
rect 13196 3236 13252 3238
rect 13358 2896 13414 2952
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 16982 8186
rect 16982 8134 17012 8186
rect 17036 8134 17046 8186
rect 17046 8134 17092 8186
rect 17116 8134 17162 8186
rect 17162 8134 17172 8186
rect 17196 8134 17226 8186
rect 17226 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 17406 7928 17462 7984
rect 21270 19760 21326 19816
rect 20956 19610 21012 19612
rect 21036 19610 21092 19612
rect 21116 19610 21172 19612
rect 21196 19610 21252 19612
rect 20956 19558 20982 19610
rect 20982 19558 21012 19610
rect 21036 19558 21046 19610
rect 21046 19558 21092 19610
rect 21116 19558 21162 19610
rect 21162 19558 21172 19610
rect 21196 19558 21226 19610
rect 21226 19558 21252 19610
rect 20956 19556 21012 19558
rect 21036 19556 21092 19558
rect 21116 19556 21172 19558
rect 21196 19556 21252 19558
rect 21270 18672 21326 18728
rect 20956 18522 21012 18524
rect 21036 18522 21092 18524
rect 21116 18522 21172 18524
rect 21196 18522 21252 18524
rect 20956 18470 20982 18522
rect 20982 18470 21012 18522
rect 21036 18470 21046 18522
rect 21046 18470 21092 18522
rect 21116 18470 21162 18522
rect 21162 18470 21172 18522
rect 21196 18470 21226 18522
rect 21226 18470 21252 18522
rect 20956 18468 21012 18470
rect 21036 18468 21092 18470
rect 21116 18468 21172 18470
rect 21196 18468 21252 18470
rect 20956 17434 21012 17436
rect 21036 17434 21092 17436
rect 21116 17434 21172 17436
rect 21196 17434 21252 17436
rect 20956 17382 20982 17434
rect 20982 17382 21012 17434
rect 21036 17382 21046 17434
rect 21046 17382 21092 17434
rect 21116 17382 21162 17434
rect 21162 17382 21172 17434
rect 21196 17382 21226 17434
rect 21226 17382 21252 17434
rect 20956 17380 21012 17382
rect 21036 17380 21092 17382
rect 21116 17380 21172 17382
rect 21196 17380 21252 17382
rect 21270 17040 21326 17096
rect 20956 16346 21012 16348
rect 21036 16346 21092 16348
rect 21116 16346 21172 16348
rect 21196 16346 21252 16348
rect 20956 16294 20982 16346
rect 20982 16294 21012 16346
rect 21036 16294 21046 16346
rect 21046 16294 21092 16346
rect 21116 16294 21162 16346
rect 21162 16294 21172 16346
rect 21196 16294 21226 16346
rect 21226 16294 21252 16346
rect 20956 16292 21012 16294
rect 21036 16292 21092 16294
rect 21116 16292 21172 16294
rect 21196 16292 21252 16294
rect 20956 15258 21012 15260
rect 21036 15258 21092 15260
rect 21116 15258 21172 15260
rect 21196 15258 21252 15260
rect 20956 15206 20982 15258
rect 20982 15206 21012 15258
rect 21036 15206 21046 15258
rect 21046 15206 21092 15258
rect 21116 15206 21162 15258
rect 21162 15206 21172 15258
rect 21196 15206 21226 15258
rect 21226 15206 21252 15258
rect 20956 15204 21012 15206
rect 21036 15204 21092 15206
rect 21116 15204 21172 15206
rect 21196 15204 21252 15206
rect 21454 14184 21510 14240
rect 20956 14170 21012 14172
rect 21036 14170 21092 14172
rect 21116 14170 21172 14172
rect 21196 14170 21252 14172
rect 20956 14118 20982 14170
rect 20982 14118 21012 14170
rect 21036 14118 21046 14170
rect 21046 14118 21092 14170
rect 21116 14118 21162 14170
rect 21162 14118 21172 14170
rect 21196 14118 21226 14170
rect 21226 14118 21252 14170
rect 20956 14116 21012 14118
rect 21036 14116 21092 14118
rect 21116 14116 21172 14118
rect 21196 14116 21252 14118
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 21454 11872 21510 11928
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 19338 9424 19394 9480
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 16982 7098
rect 16982 7046 17012 7098
rect 17036 7046 17046 7098
rect 17046 7046 17092 7098
rect 17116 7046 17162 7098
rect 17162 7046 17172 7098
rect 17196 7046 17226 7098
rect 17226 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 16982 6010
rect 16982 5958 17012 6010
rect 17036 5958 17046 6010
rect 17046 5958 17092 6010
rect 17116 5958 17162 6010
rect 17162 5958 17172 6010
rect 17196 5958 17226 6010
rect 17226 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 16982 4922
rect 16982 4870 17012 4922
rect 17036 4870 17046 4922
rect 17046 4870 17092 4922
rect 17116 4870 17162 4922
rect 17162 4870 17172 4922
rect 17196 4870 17226 4922
rect 17226 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 16982 3834
rect 16982 3782 17012 3834
rect 17036 3782 17046 3834
rect 17046 3782 17092 3834
rect 17116 3782 17162 3834
rect 17162 3782 17172 3834
rect 17196 3782 17226 3834
rect 17226 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 16982 2746
rect 16982 2694 17012 2746
rect 17036 2694 17046 2746
rect 17046 2694 17092 2746
rect 17116 2694 17162 2746
rect 17162 2694 17172 2746
rect 17196 2694 17226 2746
rect 17226 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 16026 2352 16082 2408
rect 12956 2202 13012 2204
rect 13036 2202 13092 2204
rect 13116 2202 13172 2204
rect 13196 2202 13252 2204
rect 12956 2150 12982 2202
rect 12982 2150 13012 2202
rect 13036 2150 13046 2202
rect 13046 2150 13092 2202
rect 13116 2150 13162 2202
rect 13162 2150 13172 2202
rect 13196 2150 13226 2202
rect 13226 2150 13252 2202
rect 12956 2148 13012 2150
rect 13036 2148 13092 2150
rect 13116 2148 13172 2150
rect 13196 2148 13252 2150
rect 17222 1944 17278 2000
rect 17498 1264 17554 1320
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 22190 12824 22246 12880
rect 22098 10548 22100 10568
rect 22100 10548 22152 10568
rect 22152 10548 22154 10568
rect 22098 10512 22154 10548
rect 21454 8744 21510 8800
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 21362 7656 21418 7712
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 20074 4936 20130 4992
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 21730 5888 21786 5944
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
<< metal3 >>
rect 0 23264 480 23384
rect 62 22810 122 23264
rect 23520 23128 24000 23248
rect 5809 22810 5875 22813
rect 62 22808 5875 22810
rect 62 22752 5814 22808
rect 5870 22752 5875 22808
rect 62 22750 5875 22752
rect 5809 22747 5875 22750
rect 21633 22674 21699 22677
rect 23614 22674 23674 23128
rect 21633 22672 23674 22674
rect 21633 22616 21638 22672
rect 21694 22616 23674 22672
rect 21633 22614 23674 22616
rect 21633 22611 21699 22614
rect 0 22040 480 22160
rect 62 21586 122 22040
rect 23520 21858 24000 21888
rect 23484 21856 24000 21858
rect 23484 21800 23570 21856
rect 23626 21800 24000 21856
rect 23484 21798 24000 21800
rect 4944 21792 5264 21793
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 21727 5264 21728
rect 12944 21792 13264 21793
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 21727 13264 21728
rect 20944 21792 21264 21793
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 23520 21768 24000 21798
rect 20944 21727 21264 21728
rect 1209 21586 1275 21589
rect 62 21584 1275 21586
rect 62 21528 1214 21584
rect 1270 21528 1275 21584
rect 62 21526 1275 21528
rect 1209 21523 1275 21526
rect 8944 21248 9264 21249
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 21183 9264 21184
rect 16944 21248 17264 21249
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 21183 17264 21184
rect 0 20816 480 20936
rect 62 20362 122 20816
rect 4944 20704 5264 20705
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 20639 5264 20640
rect 12944 20704 13264 20705
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 20639 13264 20640
rect 20944 20704 21264 20705
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 20639 21264 20640
rect 1301 20362 1367 20365
rect 62 20360 1367 20362
rect 62 20304 1306 20360
rect 1362 20304 1367 20360
rect 62 20302 1367 20304
rect 1301 20299 1367 20302
rect 23520 20272 24000 20392
rect 8944 20160 9264 20161
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 20095 9264 20096
rect 16944 20160 17264 20161
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 20095 17264 20096
rect 21265 19818 21331 19821
rect 23614 19818 23674 20272
rect 21265 19816 23674 19818
rect 21265 19760 21270 19816
rect 21326 19760 23674 19816
rect 21265 19758 23674 19760
rect 21265 19755 21331 19758
rect 0 19592 480 19712
rect 4944 19616 5264 19617
rect 62 19138 122 19592
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 19551 5264 19552
rect 12944 19616 13264 19617
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 19551 13264 19552
rect 20944 19616 21264 19617
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 19551 21264 19552
rect 1209 19138 1275 19141
rect 62 19136 1275 19138
rect 62 19080 1214 19136
rect 1270 19080 1275 19136
rect 62 19078 1275 19080
rect 1209 19075 1275 19078
rect 8944 19072 9264 19073
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 19007 9264 19008
rect 16944 19072 17264 19073
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 19007 17264 19008
rect 23520 18912 24000 19032
rect 21265 18730 21331 18733
rect 23614 18730 23674 18912
rect 21265 18728 23674 18730
rect 21265 18672 21270 18728
rect 21326 18672 23674 18728
rect 21265 18670 23674 18672
rect 21265 18667 21331 18670
rect 0 18504 480 18624
rect 4944 18528 5264 18529
rect 62 18050 122 18504
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 18463 5264 18464
rect 12944 18528 13264 18529
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 18463 13264 18464
rect 20944 18528 21264 18529
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 18463 21264 18464
rect 1485 18050 1551 18053
rect 62 18048 1551 18050
rect 62 17992 1490 18048
rect 1546 17992 1551 18048
rect 62 17990 1551 17992
rect 1485 17987 1551 17990
rect 8944 17984 9264 17985
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 17919 9264 17920
rect 16944 17984 17264 17985
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 17919 17264 17920
rect 8385 17778 8451 17781
rect 16021 17778 16087 17781
rect 8385 17776 16087 17778
rect 8385 17720 8390 17776
rect 8446 17720 16026 17776
rect 16082 17720 16087 17776
rect 8385 17718 16087 17720
rect 8385 17715 8451 17718
rect 16021 17715 16087 17718
rect 23520 17552 24000 17672
rect 4944 17440 5264 17441
rect 0 17368 480 17400
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 17375 5264 17376
rect 12944 17440 13264 17441
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 17375 13264 17376
rect 20944 17440 21264 17441
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 17375 21264 17376
rect 0 17312 110 17368
rect 166 17312 480 17368
rect 0 17280 480 17312
rect 21265 17098 21331 17101
rect 23614 17098 23674 17552
rect 21265 17096 23674 17098
rect 21265 17040 21270 17096
rect 21326 17040 23674 17096
rect 21265 17038 23674 17040
rect 21265 17035 21331 17038
rect 8944 16896 9264 16897
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 16831 9264 16832
rect 16944 16896 17264 16897
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 16831 17264 16832
rect 54 16356 60 16420
rect 124 16418 130 16420
rect 1577 16418 1643 16421
rect 124 16416 1643 16418
rect 124 16360 1582 16416
rect 1638 16360 1643 16416
rect 124 16358 1643 16360
rect 124 16356 130 16358
rect 1577 16355 1643 16358
rect 4944 16352 5264 16353
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 16287 5264 16288
rect 12944 16352 13264 16353
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 16287 13264 16288
rect 20944 16352 21264 16353
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 16287 21264 16288
rect 0 16148 480 16176
rect 0 16084 60 16148
rect 124 16084 480 16148
rect 0 16056 480 16084
rect 23520 16056 24000 16176
rect 8944 15808 9264 15809
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 15743 9264 15744
rect 16944 15808 17264 15809
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 15743 17264 15744
rect 14549 15602 14615 15605
rect 23614 15602 23674 16056
rect 14549 15600 23674 15602
rect 14549 15544 14554 15600
rect 14610 15544 23674 15600
rect 14549 15542 23674 15544
rect 14549 15539 14615 15542
rect 1945 15466 2011 15469
rect 62 15464 2011 15466
rect 62 15408 1950 15464
rect 2006 15408 2011 15464
rect 62 15406 2011 15408
rect 62 14952 122 15406
rect 1945 15403 2011 15406
rect 4944 15264 5264 15265
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 15199 5264 15200
rect 12944 15264 13264 15265
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 15199 13264 15200
rect 20944 15264 21264 15265
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 15199 21264 15200
rect 2037 15058 2103 15061
rect 8937 15058 9003 15061
rect 2037 15056 9003 15058
rect 2037 15000 2042 15056
rect 2098 15000 8942 15056
rect 8998 15000 9003 15056
rect 2037 14998 9003 15000
rect 2037 14995 2103 14998
rect 8937 14995 9003 14998
rect 0 14832 480 14952
rect 8944 14720 9264 14721
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 14655 9264 14656
rect 16944 14720 17264 14721
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 23520 14696 24000 14816
rect 16944 14655 17264 14656
rect 21449 14242 21515 14245
rect 23614 14242 23674 14696
rect 21449 14240 23674 14242
rect 21449 14184 21454 14240
rect 21510 14184 23674 14240
rect 21449 14182 23674 14184
rect 21449 14179 21515 14182
rect 4944 14176 5264 14177
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 14111 5264 14112
rect 12944 14176 13264 14177
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 14111 13264 14112
rect 20944 14176 21264 14177
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 14111 21264 14112
rect 9397 13834 9463 13837
rect 9673 13834 9739 13837
rect 9270 13832 9739 13834
rect 9270 13776 9402 13832
rect 9458 13776 9678 13832
rect 9734 13776 9739 13832
rect 9270 13774 9739 13776
rect 9397 13771 9463 13774
rect 9673 13771 9739 13774
rect 0 13608 480 13728
rect 8944 13632 9264 13633
rect 62 13290 122 13608
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 13567 9264 13568
rect 16944 13632 17264 13633
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13567 17264 13568
rect 23520 13336 24000 13456
rect 7373 13290 7439 13293
rect 62 13288 7439 13290
rect 62 13232 7378 13288
rect 7434 13232 7439 13288
rect 62 13230 7439 13232
rect 7373 13227 7439 13230
rect 4944 13088 5264 13089
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 13023 5264 13024
rect 12944 13088 13264 13089
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 13023 13264 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 22185 12882 22251 12885
rect 23614 12882 23674 13336
rect 22185 12880 23674 12882
rect 22185 12824 22190 12880
rect 22246 12824 23674 12880
rect 22185 12822 23674 12824
rect 22185 12819 22251 12822
rect 0 12520 480 12640
rect 8944 12544 9264 12545
rect 62 12066 122 12520
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 12479 9264 12480
rect 16944 12544 17264 12545
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 12479 17264 12480
rect 1117 12066 1183 12069
rect 62 12064 1183 12066
rect 62 12008 1122 12064
rect 1178 12008 1183 12064
rect 62 12006 1183 12008
rect 1117 12003 1183 12006
rect 4944 12000 5264 12001
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 11935 5264 11936
rect 12944 12000 13264 12001
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 11935 13264 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 21449 11930 21515 11933
rect 23520 11930 24000 11960
rect 21449 11928 24000 11930
rect 21449 11872 21454 11928
rect 21510 11872 24000 11928
rect 21449 11870 24000 11872
rect 21449 11867 21515 11870
rect 23520 11840 24000 11870
rect 8944 11456 9264 11457
rect 0 11296 480 11416
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 11391 9264 11392
rect 16944 11456 17264 11457
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 11391 17264 11392
rect 62 11114 122 11296
rect 5809 11114 5875 11117
rect 62 11112 5875 11114
rect 62 11056 5814 11112
rect 5870 11056 5875 11112
rect 62 11054 5875 11056
rect 5809 11051 5875 11054
rect 4944 10912 5264 10913
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 10847 5264 10848
rect 12944 10912 13264 10913
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 10847 13264 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 22093 10570 22159 10573
rect 23520 10570 24000 10600
rect 22093 10568 24000 10570
rect 22093 10512 22098 10568
rect 22154 10512 24000 10568
rect 22093 10510 24000 10512
rect 22093 10507 22159 10510
rect 23520 10480 24000 10510
rect 8944 10368 9264 10369
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 10303 9264 10304
rect 16944 10368 17264 10369
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 10303 17264 10304
rect 0 10160 480 10192
rect 0 10104 18 10160
rect 74 10104 480 10160
rect 0 10072 480 10104
rect 4944 9824 5264 9825
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 9759 5264 9760
rect 12944 9824 13264 9825
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 9759 13264 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 3417 9482 3483 9485
rect 19333 9482 19399 9485
rect 3417 9480 19399 9482
rect 3417 9424 3422 9480
rect 3478 9424 19338 9480
rect 19394 9424 19399 9480
rect 3417 9422 19399 9424
rect 3417 9419 3483 9422
rect 19333 9419 19399 9422
rect 8944 9280 9264 9281
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 9215 9264 9216
rect 16944 9280 17264 9281
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 9215 17264 9216
rect 23520 9120 24000 9240
rect 0 8936 480 8968
rect 0 8880 110 8936
rect 166 8880 480 8936
rect 0 8848 480 8880
rect 8109 8938 8175 8941
rect 17125 8938 17191 8941
rect 8109 8936 17191 8938
rect 8109 8880 8114 8936
rect 8170 8880 17130 8936
rect 17186 8880 17191 8936
rect 8109 8878 17191 8880
rect 8109 8875 8175 8878
rect 17125 8875 17191 8878
rect 21449 8802 21515 8805
rect 23614 8802 23674 9120
rect 21449 8800 23674 8802
rect 21449 8744 21454 8800
rect 21510 8744 23674 8800
rect 21449 8742 23674 8744
rect 21449 8739 21515 8742
rect 4944 8736 5264 8737
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 8671 5264 8672
rect 12944 8736 13264 8737
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 8671 13264 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 8944 8192 9264 8193
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 8127 9264 8128
rect 16944 8192 17264 8193
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 8127 17264 8128
rect 10317 7986 10383 7989
rect 17401 7986 17467 7989
rect 10317 7984 17467 7986
rect 10317 7928 10322 7984
rect 10378 7928 17406 7984
rect 17462 7928 17467 7984
rect 10317 7926 17467 7928
rect 10317 7923 10383 7926
rect 17401 7923 17467 7926
rect 0 7712 480 7744
rect 0 7656 110 7712
rect 166 7656 480 7712
rect 0 7624 480 7656
rect 21357 7714 21423 7717
rect 23520 7714 24000 7744
rect 21357 7712 24000 7714
rect 21357 7656 21362 7712
rect 21418 7656 24000 7712
rect 21357 7654 24000 7656
rect 21357 7651 21423 7654
rect 4944 7648 5264 7649
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 7583 5264 7584
rect 12944 7648 13264 7649
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 7583 13264 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 23520 7624 24000 7654
rect 20944 7583 21264 7584
rect 8944 7104 9264 7105
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 7039 9264 7040
rect 16944 7104 17264 7105
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 7039 17264 7040
rect 0 6624 480 6656
rect 0 6568 110 6624
rect 166 6568 480 6624
rect 0 6536 480 6568
rect 4944 6560 5264 6561
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 6495 5264 6496
rect 12944 6560 13264 6561
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 6495 13264 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 23520 6264 24000 6384
rect 8944 6016 9264 6017
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 5951 9264 5952
rect 16944 6016 17264 6017
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 5951 17264 5952
rect 21725 5946 21791 5949
rect 23614 5946 23674 6264
rect 21725 5944 23674 5946
rect 21725 5888 21730 5944
rect 21786 5888 23674 5944
rect 21725 5886 23674 5888
rect 21725 5883 21791 5886
rect 4944 5472 5264 5473
rect 0 5400 480 5432
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 5407 5264 5408
rect 12944 5472 13264 5473
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 5407 13264 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 0 5344 110 5400
rect 166 5344 480 5400
rect 0 5312 480 5344
rect 20069 4994 20135 4997
rect 23520 4994 24000 5024
rect 20069 4992 24000 4994
rect 20069 4936 20074 4992
rect 20130 4936 24000 4992
rect 20069 4934 24000 4936
rect 20069 4931 20135 4934
rect 8944 4928 9264 4929
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 4863 9264 4864
rect 16944 4928 17264 4929
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 23520 4904 24000 4934
rect 16944 4863 17264 4864
rect 4944 4384 5264 4385
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 4319 5264 4320
rect 12944 4384 13264 4385
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 4319 13264 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 0 4142 480 4208
rect 0 4088 110 4142
rect 105 4086 110 4088
rect 166 4088 480 4142
rect 166 4086 252 4088
rect 105 4084 252 4086
rect 105 4081 171 4084
rect 8944 3840 9264 3841
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 3775 9264 3776
rect 16944 3840 17264 3841
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3775 17264 3776
rect 11789 3498 11855 3501
rect 23520 3498 24000 3528
rect 11789 3496 24000 3498
rect 11789 3440 11794 3496
rect 11850 3440 24000 3496
rect 11789 3438 24000 3440
rect 11789 3435 11855 3438
rect 23520 3408 24000 3438
rect 4944 3296 5264 3297
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 3231 5264 3232
rect 12944 3296 13264 3297
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 3231 13264 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 0 2952 480 2984
rect 0 2896 110 2952
rect 166 2896 480 2952
rect 0 2864 480 2896
rect 2313 2954 2379 2957
rect 13353 2954 13419 2957
rect 2313 2952 13419 2954
rect 2313 2896 2318 2952
rect 2374 2896 13358 2952
rect 13414 2896 13419 2952
rect 2313 2894 13419 2896
rect 2313 2891 2379 2894
rect 13353 2891 13419 2894
rect 8944 2752 9264 2753
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2687 9264 2688
rect 16944 2752 17264 2753
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2687 17264 2688
rect 7741 2546 7807 2549
rect 7741 2544 23674 2546
rect 7741 2488 7746 2544
rect 7802 2488 23674 2544
rect 7741 2486 23674 2488
rect 7741 2483 7807 2486
rect 4521 2410 4587 2413
rect 16021 2410 16087 2413
rect 4521 2408 16087 2410
rect 4521 2352 4526 2408
rect 4582 2352 16026 2408
rect 16082 2352 16087 2408
rect 4521 2350 16087 2352
rect 4521 2347 4587 2350
rect 16021 2347 16087 2350
rect 1853 2274 1919 2277
rect 62 2272 1919 2274
rect 62 2216 1858 2272
rect 1914 2216 1919 2272
rect 62 2214 1919 2216
rect 62 1760 122 2214
rect 1853 2211 1919 2214
rect 4944 2208 5264 2209
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2143 5264 2144
rect 12944 2208 13264 2209
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2143 13264 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 23614 2168 23674 2486
rect 20944 2143 21264 2144
rect 23520 2048 24000 2168
rect 8753 2002 8819 2005
rect 17217 2002 17283 2005
rect 8753 2000 17283 2002
rect 8753 1944 8758 2000
rect 8814 1944 17222 2000
rect 17278 1944 17283 2000
rect 8753 1942 17283 1944
rect 8753 1939 8819 1942
rect 17217 1939 17283 1942
rect 0 1640 480 1760
rect 17493 1322 17559 1325
rect 17493 1320 23674 1322
rect 17493 1264 17498 1320
rect 17554 1264 23674 1320
rect 17493 1262 23674 1264
rect 17493 1259 17559 1262
rect 6729 1186 6795 1189
rect 62 1184 6795 1186
rect 62 1128 6734 1184
rect 6790 1128 6795 1184
rect 62 1126 6795 1128
rect 62 672 122 1126
rect 6729 1123 6795 1126
rect 23614 808 23674 1262
rect 23520 688 24000 808
rect 0 552 480 672
<< via3 >>
rect 4952 21788 5016 21792
rect 4952 21732 4956 21788
rect 4956 21732 5012 21788
rect 5012 21732 5016 21788
rect 4952 21728 5016 21732
rect 5032 21788 5096 21792
rect 5032 21732 5036 21788
rect 5036 21732 5092 21788
rect 5092 21732 5096 21788
rect 5032 21728 5096 21732
rect 5112 21788 5176 21792
rect 5112 21732 5116 21788
rect 5116 21732 5172 21788
rect 5172 21732 5176 21788
rect 5112 21728 5176 21732
rect 5192 21788 5256 21792
rect 5192 21732 5196 21788
rect 5196 21732 5252 21788
rect 5252 21732 5256 21788
rect 5192 21728 5256 21732
rect 12952 21788 13016 21792
rect 12952 21732 12956 21788
rect 12956 21732 13012 21788
rect 13012 21732 13016 21788
rect 12952 21728 13016 21732
rect 13032 21788 13096 21792
rect 13032 21732 13036 21788
rect 13036 21732 13092 21788
rect 13092 21732 13096 21788
rect 13032 21728 13096 21732
rect 13112 21788 13176 21792
rect 13112 21732 13116 21788
rect 13116 21732 13172 21788
rect 13172 21732 13176 21788
rect 13112 21728 13176 21732
rect 13192 21788 13256 21792
rect 13192 21732 13196 21788
rect 13196 21732 13252 21788
rect 13252 21732 13256 21788
rect 13192 21728 13256 21732
rect 20952 21788 21016 21792
rect 20952 21732 20956 21788
rect 20956 21732 21012 21788
rect 21012 21732 21016 21788
rect 20952 21728 21016 21732
rect 21032 21788 21096 21792
rect 21032 21732 21036 21788
rect 21036 21732 21092 21788
rect 21092 21732 21096 21788
rect 21032 21728 21096 21732
rect 21112 21788 21176 21792
rect 21112 21732 21116 21788
rect 21116 21732 21172 21788
rect 21172 21732 21176 21788
rect 21112 21728 21176 21732
rect 21192 21788 21256 21792
rect 21192 21732 21196 21788
rect 21196 21732 21252 21788
rect 21252 21732 21256 21788
rect 21192 21728 21256 21732
rect 8952 21244 9016 21248
rect 8952 21188 8956 21244
rect 8956 21188 9012 21244
rect 9012 21188 9016 21244
rect 8952 21184 9016 21188
rect 9032 21244 9096 21248
rect 9032 21188 9036 21244
rect 9036 21188 9092 21244
rect 9092 21188 9096 21244
rect 9032 21184 9096 21188
rect 9112 21244 9176 21248
rect 9112 21188 9116 21244
rect 9116 21188 9172 21244
rect 9172 21188 9176 21244
rect 9112 21184 9176 21188
rect 9192 21244 9256 21248
rect 9192 21188 9196 21244
rect 9196 21188 9252 21244
rect 9252 21188 9256 21244
rect 9192 21184 9256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 4952 20700 5016 20704
rect 4952 20644 4956 20700
rect 4956 20644 5012 20700
rect 5012 20644 5016 20700
rect 4952 20640 5016 20644
rect 5032 20700 5096 20704
rect 5032 20644 5036 20700
rect 5036 20644 5092 20700
rect 5092 20644 5096 20700
rect 5032 20640 5096 20644
rect 5112 20700 5176 20704
rect 5112 20644 5116 20700
rect 5116 20644 5172 20700
rect 5172 20644 5176 20700
rect 5112 20640 5176 20644
rect 5192 20700 5256 20704
rect 5192 20644 5196 20700
rect 5196 20644 5252 20700
rect 5252 20644 5256 20700
rect 5192 20640 5256 20644
rect 12952 20700 13016 20704
rect 12952 20644 12956 20700
rect 12956 20644 13012 20700
rect 13012 20644 13016 20700
rect 12952 20640 13016 20644
rect 13032 20700 13096 20704
rect 13032 20644 13036 20700
rect 13036 20644 13092 20700
rect 13092 20644 13096 20700
rect 13032 20640 13096 20644
rect 13112 20700 13176 20704
rect 13112 20644 13116 20700
rect 13116 20644 13172 20700
rect 13172 20644 13176 20700
rect 13112 20640 13176 20644
rect 13192 20700 13256 20704
rect 13192 20644 13196 20700
rect 13196 20644 13252 20700
rect 13252 20644 13256 20700
rect 13192 20640 13256 20644
rect 20952 20700 21016 20704
rect 20952 20644 20956 20700
rect 20956 20644 21012 20700
rect 21012 20644 21016 20700
rect 20952 20640 21016 20644
rect 21032 20700 21096 20704
rect 21032 20644 21036 20700
rect 21036 20644 21092 20700
rect 21092 20644 21096 20700
rect 21032 20640 21096 20644
rect 21112 20700 21176 20704
rect 21112 20644 21116 20700
rect 21116 20644 21172 20700
rect 21172 20644 21176 20700
rect 21112 20640 21176 20644
rect 21192 20700 21256 20704
rect 21192 20644 21196 20700
rect 21196 20644 21252 20700
rect 21252 20644 21256 20700
rect 21192 20640 21256 20644
rect 8952 20156 9016 20160
rect 8952 20100 8956 20156
rect 8956 20100 9012 20156
rect 9012 20100 9016 20156
rect 8952 20096 9016 20100
rect 9032 20156 9096 20160
rect 9032 20100 9036 20156
rect 9036 20100 9092 20156
rect 9092 20100 9096 20156
rect 9032 20096 9096 20100
rect 9112 20156 9176 20160
rect 9112 20100 9116 20156
rect 9116 20100 9172 20156
rect 9172 20100 9176 20156
rect 9112 20096 9176 20100
rect 9192 20156 9256 20160
rect 9192 20100 9196 20156
rect 9196 20100 9252 20156
rect 9252 20100 9256 20156
rect 9192 20096 9256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 4952 19612 5016 19616
rect 4952 19556 4956 19612
rect 4956 19556 5012 19612
rect 5012 19556 5016 19612
rect 4952 19552 5016 19556
rect 5032 19612 5096 19616
rect 5032 19556 5036 19612
rect 5036 19556 5092 19612
rect 5092 19556 5096 19612
rect 5032 19552 5096 19556
rect 5112 19612 5176 19616
rect 5112 19556 5116 19612
rect 5116 19556 5172 19612
rect 5172 19556 5176 19612
rect 5112 19552 5176 19556
rect 5192 19612 5256 19616
rect 5192 19556 5196 19612
rect 5196 19556 5252 19612
rect 5252 19556 5256 19612
rect 5192 19552 5256 19556
rect 12952 19612 13016 19616
rect 12952 19556 12956 19612
rect 12956 19556 13012 19612
rect 13012 19556 13016 19612
rect 12952 19552 13016 19556
rect 13032 19612 13096 19616
rect 13032 19556 13036 19612
rect 13036 19556 13092 19612
rect 13092 19556 13096 19612
rect 13032 19552 13096 19556
rect 13112 19612 13176 19616
rect 13112 19556 13116 19612
rect 13116 19556 13172 19612
rect 13172 19556 13176 19612
rect 13112 19552 13176 19556
rect 13192 19612 13256 19616
rect 13192 19556 13196 19612
rect 13196 19556 13252 19612
rect 13252 19556 13256 19612
rect 13192 19552 13256 19556
rect 20952 19612 21016 19616
rect 20952 19556 20956 19612
rect 20956 19556 21012 19612
rect 21012 19556 21016 19612
rect 20952 19552 21016 19556
rect 21032 19612 21096 19616
rect 21032 19556 21036 19612
rect 21036 19556 21092 19612
rect 21092 19556 21096 19612
rect 21032 19552 21096 19556
rect 21112 19612 21176 19616
rect 21112 19556 21116 19612
rect 21116 19556 21172 19612
rect 21172 19556 21176 19612
rect 21112 19552 21176 19556
rect 21192 19612 21256 19616
rect 21192 19556 21196 19612
rect 21196 19556 21252 19612
rect 21252 19556 21256 19612
rect 21192 19552 21256 19556
rect 8952 19068 9016 19072
rect 8952 19012 8956 19068
rect 8956 19012 9012 19068
rect 9012 19012 9016 19068
rect 8952 19008 9016 19012
rect 9032 19068 9096 19072
rect 9032 19012 9036 19068
rect 9036 19012 9092 19068
rect 9092 19012 9096 19068
rect 9032 19008 9096 19012
rect 9112 19068 9176 19072
rect 9112 19012 9116 19068
rect 9116 19012 9172 19068
rect 9172 19012 9176 19068
rect 9112 19008 9176 19012
rect 9192 19068 9256 19072
rect 9192 19012 9196 19068
rect 9196 19012 9252 19068
rect 9252 19012 9256 19068
rect 9192 19008 9256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 4952 18524 5016 18528
rect 4952 18468 4956 18524
rect 4956 18468 5012 18524
rect 5012 18468 5016 18524
rect 4952 18464 5016 18468
rect 5032 18524 5096 18528
rect 5032 18468 5036 18524
rect 5036 18468 5092 18524
rect 5092 18468 5096 18524
rect 5032 18464 5096 18468
rect 5112 18524 5176 18528
rect 5112 18468 5116 18524
rect 5116 18468 5172 18524
rect 5172 18468 5176 18524
rect 5112 18464 5176 18468
rect 5192 18524 5256 18528
rect 5192 18468 5196 18524
rect 5196 18468 5252 18524
rect 5252 18468 5256 18524
rect 5192 18464 5256 18468
rect 12952 18524 13016 18528
rect 12952 18468 12956 18524
rect 12956 18468 13012 18524
rect 13012 18468 13016 18524
rect 12952 18464 13016 18468
rect 13032 18524 13096 18528
rect 13032 18468 13036 18524
rect 13036 18468 13092 18524
rect 13092 18468 13096 18524
rect 13032 18464 13096 18468
rect 13112 18524 13176 18528
rect 13112 18468 13116 18524
rect 13116 18468 13172 18524
rect 13172 18468 13176 18524
rect 13112 18464 13176 18468
rect 13192 18524 13256 18528
rect 13192 18468 13196 18524
rect 13196 18468 13252 18524
rect 13252 18468 13256 18524
rect 13192 18464 13256 18468
rect 20952 18524 21016 18528
rect 20952 18468 20956 18524
rect 20956 18468 21012 18524
rect 21012 18468 21016 18524
rect 20952 18464 21016 18468
rect 21032 18524 21096 18528
rect 21032 18468 21036 18524
rect 21036 18468 21092 18524
rect 21092 18468 21096 18524
rect 21032 18464 21096 18468
rect 21112 18524 21176 18528
rect 21112 18468 21116 18524
rect 21116 18468 21172 18524
rect 21172 18468 21176 18524
rect 21112 18464 21176 18468
rect 21192 18524 21256 18528
rect 21192 18468 21196 18524
rect 21196 18468 21252 18524
rect 21252 18468 21256 18524
rect 21192 18464 21256 18468
rect 8952 17980 9016 17984
rect 8952 17924 8956 17980
rect 8956 17924 9012 17980
rect 9012 17924 9016 17980
rect 8952 17920 9016 17924
rect 9032 17980 9096 17984
rect 9032 17924 9036 17980
rect 9036 17924 9092 17980
rect 9092 17924 9096 17980
rect 9032 17920 9096 17924
rect 9112 17980 9176 17984
rect 9112 17924 9116 17980
rect 9116 17924 9172 17980
rect 9172 17924 9176 17980
rect 9112 17920 9176 17924
rect 9192 17980 9256 17984
rect 9192 17924 9196 17980
rect 9196 17924 9252 17980
rect 9252 17924 9256 17980
rect 9192 17920 9256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 4952 17436 5016 17440
rect 4952 17380 4956 17436
rect 4956 17380 5012 17436
rect 5012 17380 5016 17436
rect 4952 17376 5016 17380
rect 5032 17436 5096 17440
rect 5032 17380 5036 17436
rect 5036 17380 5092 17436
rect 5092 17380 5096 17436
rect 5032 17376 5096 17380
rect 5112 17436 5176 17440
rect 5112 17380 5116 17436
rect 5116 17380 5172 17436
rect 5172 17380 5176 17436
rect 5112 17376 5176 17380
rect 5192 17436 5256 17440
rect 5192 17380 5196 17436
rect 5196 17380 5252 17436
rect 5252 17380 5256 17436
rect 5192 17376 5256 17380
rect 12952 17436 13016 17440
rect 12952 17380 12956 17436
rect 12956 17380 13012 17436
rect 13012 17380 13016 17436
rect 12952 17376 13016 17380
rect 13032 17436 13096 17440
rect 13032 17380 13036 17436
rect 13036 17380 13092 17436
rect 13092 17380 13096 17436
rect 13032 17376 13096 17380
rect 13112 17436 13176 17440
rect 13112 17380 13116 17436
rect 13116 17380 13172 17436
rect 13172 17380 13176 17436
rect 13112 17376 13176 17380
rect 13192 17436 13256 17440
rect 13192 17380 13196 17436
rect 13196 17380 13252 17436
rect 13252 17380 13256 17436
rect 13192 17376 13256 17380
rect 20952 17436 21016 17440
rect 20952 17380 20956 17436
rect 20956 17380 21012 17436
rect 21012 17380 21016 17436
rect 20952 17376 21016 17380
rect 21032 17436 21096 17440
rect 21032 17380 21036 17436
rect 21036 17380 21092 17436
rect 21092 17380 21096 17436
rect 21032 17376 21096 17380
rect 21112 17436 21176 17440
rect 21112 17380 21116 17436
rect 21116 17380 21172 17436
rect 21172 17380 21176 17436
rect 21112 17376 21176 17380
rect 21192 17436 21256 17440
rect 21192 17380 21196 17436
rect 21196 17380 21252 17436
rect 21252 17380 21256 17436
rect 21192 17376 21256 17380
rect 8952 16892 9016 16896
rect 8952 16836 8956 16892
rect 8956 16836 9012 16892
rect 9012 16836 9016 16892
rect 8952 16832 9016 16836
rect 9032 16892 9096 16896
rect 9032 16836 9036 16892
rect 9036 16836 9092 16892
rect 9092 16836 9096 16892
rect 9032 16832 9096 16836
rect 9112 16892 9176 16896
rect 9112 16836 9116 16892
rect 9116 16836 9172 16892
rect 9172 16836 9176 16892
rect 9112 16832 9176 16836
rect 9192 16892 9256 16896
rect 9192 16836 9196 16892
rect 9196 16836 9252 16892
rect 9252 16836 9256 16892
rect 9192 16832 9256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 60 16356 124 16420
rect 4952 16348 5016 16352
rect 4952 16292 4956 16348
rect 4956 16292 5012 16348
rect 5012 16292 5016 16348
rect 4952 16288 5016 16292
rect 5032 16348 5096 16352
rect 5032 16292 5036 16348
rect 5036 16292 5092 16348
rect 5092 16292 5096 16348
rect 5032 16288 5096 16292
rect 5112 16348 5176 16352
rect 5112 16292 5116 16348
rect 5116 16292 5172 16348
rect 5172 16292 5176 16348
rect 5112 16288 5176 16292
rect 5192 16348 5256 16352
rect 5192 16292 5196 16348
rect 5196 16292 5252 16348
rect 5252 16292 5256 16348
rect 5192 16288 5256 16292
rect 12952 16348 13016 16352
rect 12952 16292 12956 16348
rect 12956 16292 13012 16348
rect 13012 16292 13016 16348
rect 12952 16288 13016 16292
rect 13032 16348 13096 16352
rect 13032 16292 13036 16348
rect 13036 16292 13092 16348
rect 13092 16292 13096 16348
rect 13032 16288 13096 16292
rect 13112 16348 13176 16352
rect 13112 16292 13116 16348
rect 13116 16292 13172 16348
rect 13172 16292 13176 16348
rect 13112 16288 13176 16292
rect 13192 16348 13256 16352
rect 13192 16292 13196 16348
rect 13196 16292 13252 16348
rect 13252 16292 13256 16348
rect 13192 16288 13256 16292
rect 20952 16348 21016 16352
rect 20952 16292 20956 16348
rect 20956 16292 21012 16348
rect 21012 16292 21016 16348
rect 20952 16288 21016 16292
rect 21032 16348 21096 16352
rect 21032 16292 21036 16348
rect 21036 16292 21092 16348
rect 21092 16292 21096 16348
rect 21032 16288 21096 16292
rect 21112 16348 21176 16352
rect 21112 16292 21116 16348
rect 21116 16292 21172 16348
rect 21172 16292 21176 16348
rect 21112 16288 21176 16292
rect 21192 16348 21256 16352
rect 21192 16292 21196 16348
rect 21196 16292 21252 16348
rect 21252 16292 21256 16348
rect 21192 16288 21256 16292
rect 60 16084 124 16148
rect 8952 15804 9016 15808
rect 8952 15748 8956 15804
rect 8956 15748 9012 15804
rect 9012 15748 9016 15804
rect 8952 15744 9016 15748
rect 9032 15804 9096 15808
rect 9032 15748 9036 15804
rect 9036 15748 9092 15804
rect 9092 15748 9096 15804
rect 9032 15744 9096 15748
rect 9112 15804 9176 15808
rect 9112 15748 9116 15804
rect 9116 15748 9172 15804
rect 9172 15748 9176 15804
rect 9112 15744 9176 15748
rect 9192 15804 9256 15808
rect 9192 15748 9196 15804
rect 9196 15748 9252 15804
rect 9252 15748 9256 15804
rect 9192 15744 9256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 4952 15260 5016 15264
rect 4952 15204 4956 15260
rect 4956 15204 5012 15260
rect 5012 15204 5016 15260
rect 4952 15200 5016 15204
rect 5032 15260 5096 15264
rect 5032 15204 5036 15260
rect 5036 15204 5092 15260
rect 5092 15204 5096 15260
rect 5032 15200 5096 15204
rect 5112 15260 5176 15264
rect 5112 15204 5116 15260
rect 5116 15204 5172 15260
rect 5172 15204 5176 15260
rect 5112 15200 5176 15204
rect 5192 15260 5256 15264
rect 5192 15204 5196 15260
rect 5196 15204 5252 15260
rect 5252 15204 5256 15260
rect 5192 15200 5256 15204
rect 12952 15260 13016 15264
rect 12952 15204 12956 15260
rect 12956 15204 13012 15260
rect 13012 15204 13016 15260
rect 12952 15200 13016 15204
rect 13032 15260 13096 15264
rect 13032 15204 13036 15260
rect 13036 15204 13092 15260
rect 13092 15204 13096 15260
rect 13032 15200 13096 15204
rect 13112 15260 13176 15264
rect 13112 15204 13116 15260
rect 13116 15204 13172 15260
rect 13172 15204 13176 15260
rect 13112 15200 13176 15204
rect 13192 15260 13256 15264
rect 13192 15204 13196 15260
rect 13196 15204 13252 15260
rect 13252 15204 13256 15260
rect 13192 15200 13256 15204
rect 20952 15260 21016 15264
rect 20952 15204 20956 15260
rect 20956 15204 21012 15260
rect 21012 15204 21016 15260
rect 20952 15200 21016 15204
rect 21032 15260 21096 15264
rect 21032 15204 21036 15260
rect 21036 15204 21092 15260
rect 21092 15204 21096 15260
rect 21032 15200 21096 15204
rect 21112 15260 21176 15264
rect 21112 15204 21116 15260
rect 21116 15204 21172 15260
rect 21172 15204 21176 15260
rect 21112 15200 21176 15204
rect 21192 15260 21256 15264
rect 21192 15204 21196 15260
rect 21196 15204 21252 15260
rect 21252 15204 21256 15260
rect 21192 15200 21256 15204
rect 8952 14716 9016 14720
rect 8952 14660 8956 14716
rect 8956 14660 9012 14716
rect 9012 14660 9016 14716
rect 8952 14656 9016 14660
rect 9032 14716 9096 14720
rect 9032 14660 9036 14716
rect 9036 14660 9092 14716
rect 9092 14660 9096 14716
rect 9032 14656 9096 14660
rect 9112 14716 9176 14720
rect 9112 14660 9116 14716
rect 9116 14660 9172 14716
rect 9172 14660 9176 14716
rect 9112 14656 9176 14660
rect 9192 14716 9256 14720
rect 9192 14660 9196 14716
rect 9196 14660 9252 14716
rect 9252 14660 9256 14716
rect 9192 14656 9256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 4952 14172 5016 14176
rect 4952 14116 4956 14172
rect 4956 14116 5012 14172
rect 5012 14116 5016 14172
rect 4952 14112 5016 14116
rect 5032 14172 5096 14176
rect 5032 14116 5036 14172
rect 5036 14116 5092 14172
rect 5092 14116 5096 14172
rect 5032 14112 5096 14116
rect 5112 14172 5176 14176
rect 5112 14116 5116 14172
rect 5116 14116 5172 14172
rect 5172 14116 5176 14172
rect 5112 14112 5176 14116
rect 5192 14172 5256 14176
rect 5192 14116 5196 14172
rect 5196 14116 5252 14172
rect 5252 14116 5256 14172
rect 5192 14112 5256 14116
rect 12952 14172 13016 14176
rect 12952 14116 12956 14172
rect 12956 14116 13012 14172
rect 13012 14116 13016 14172
rect 12952 14112 13016 14116
rect 13032 14172 13096 14176
rect 13032 14116 13036 14172
rect 13036 14116 13092 14172
rect 13092 14116 13096 14172
rect 13032 14112 13096 14116
rect 13112 14172 13176 14176
rect 13112 14116 13116 14172
rect 13116 14116 13172 14172
rect 13172 14116 13176 14172
rect 13112 14112 13176 14116
rect 13192 14172 13256 14176
rect 13192 14116 13196 14172
rect 13196 14116 13252 14172
rect 13252 14116 13256 14172
rect 13192 14112 13256 14116
rect 20952 14172 21016 14176
rect 20952 14116 20956 14172
rect 20956 14116 21012 14172
rect 21012 14116 21016 14172
rect 20952 14112 21016 14116
rect 21032 14172 21096 14176
rect 21032 14116 21036 14172
rect 21036 14116 21092 14172
rect 21092 14116 21096 14172
rect 21032 14112 21096 14116
rect 21112 14172 21176 14176
rect 21112 14116 21116 14172
rect 21116 14116 21172 14172
rect 21172 14116 21176 14172
rect 21112 14112 21176 14116
rect 21192 14172 21256 14176
rect 21192 14116 21196 14172
rect 21196 14116 21252 14172
rect 21252 14116 21256 14172
rect 21192 14112 21256 14116
rect 8952 13628 9016 13632
rect 8952 13572 8956 13628
rect 8956 13572 9012 13628
rect 9012 13572 9016 13628
rect 8952 13568 9016 13572
rect 9032 13628 9096 13632
rect 9032 13572 9036 13628
rect 9036 13572 9092 13628
rect 9092 13572 9096 13628
rect 9032 13568 9096 13572
rect 9112 13628 9176 13632
rect 9112 13572 9116 13628
rect 9116 13572 9172 13628
rect 9172 13572 9176 13628
rect 9112 13568 9176 13572
rect 9192 13628 9256 13632
rect 9192 13572 9196 13628
rect 9196 13572 9252 13628
rect 9252 13572 9256 13628
rect 9192 13568 9256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 4952 13084 5016 13088
rect 4952 13028 4956 13084
rect 4956 13028 5012 13084
rect 5012 13028 5016 13084
rect 4952 13024 5016 13028
rect 5032 13084 5096 13088
rect 5032 13028 5036 13084
rect 5036 13028 5092 13084
rect 5092 13028 5096 13084
rect 5032 13024 5096 13028
rect 5112 13084 5176 13088
rect 5112 13028 5116 13084
rect 5116 13028 5172 13084
rect 5172 13028 5176 13084
rect 5112 13024 5176 13028
rect 5192 13084 5256 13088
rect 5192 13028 5196 13084
rect 5196 13028 5252 13084
rect 5252 13028 5256 13084
rect 5192 13024 5256 13028
rect 12952 13084 13016 13088
rect 12952 13028 12956 13084
rect 12956 13028 13012 13084
rect 13012 13028 13016 13084
rect 12952 13024 13016 13028
rect 13032 13084 13096 13088
rect 13032 13028 13036 13084
rect 13036 13028 13092 13084
rect 13092 13028 13096 13084
rect 13032 13024 13096 13028
rect 13112 13084 13176 13088
rect 13112 13028 13116 13084
rect 13116 13028 13172 13084
rect 13172 13028 13176 13084
rect 13112 13024 13176 13028
rect 13192 13084 13256 13088
rect 13192 13028 13196 13084
rect 13196 13028 13252 13084
rect 13252 13028 13256 13084
rect 13192 13024 13256 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 8952 12540 9016 12544
rect 8952 12484 8956 12540
rect 8956 12484 9012 12540
rect 9012 12484 9016 12540
rect 8952 12480 9016 12484
rect 9032 12540 9096 12544
rect 9032 12484 9036 12540
rect 9036 12484 9092 12540
rect 9092 12484 9096 12540
rect 9032 12480 9096 12484
rect 9112 12540 9176 12544
rect 9112 12484 9116 12540
rect 9116 12484 9172 12540
rect 9172 12484 9176 12540
rect 9112 12480 9176 12484
rect 9192 12540 9256 12544
rect 9192 12484 9196 12540
rect 9196 12484 9252 12540
rect 9252 12484 9256 12540
rect 9192 12480 9256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 4952 11996 5016 12000
rect 4952 11940 4956 11996
rect 4956 11940 5012 11996
rect 5012 11940 5016 11996
rect 4952 11936 5016 11940
rect 5032 11996 5096 12000
rect 5032 11940 5036 11996
rect 5036 11940 5092 11996
rect 5092 11940 5096 11996
rect 5032 11936 5096 11940
rect 5112 11996 5176 12000
rect 5112 11940 5116 11996
rect 5116 11940 5172 11996
rect 5172 11940 5176 11996
rect 5112 11936 5176 11940
rect 5192 11996 5256 12000
rect 5192 11940 5196 11996
rect 5196 11940 5252 11996
rect 5252 11940 5256 11996
rect 5192 11936 5256 11940
rect 12952 11996 13016 12000
rect 12952 11940 12956 11996
rect 12956 11940 13012 11996
rect 13012 11940 13016 11996
rect 12952 11936 13016 11940
rect 13032 11996 13096 12000
rect 13032 11940 13036 11996
rect 13036 11940 13092 11996
rect 13092 11940 13096 11996
rect 13032 11936 13096 11940
rect 13112 11996 13176 12000
rect 13112 11940 13116 11996
rect 13116 11940 13172 11996
rect 13172 11940 13176 11996
rect 13112 11936 13176 11940
rect 13192 11996 13256 12000
rect 13192 11940 13196 11996
rect 13196 11940 13252 11996
rect 13252 11940 13256 11996
rect 13192 11936 13256 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 8952 11452 9016 11456
rect 8952 11396 8956 11452
rect 8956 11396 9012 11452
rect 9012 11396 9016 11452
rect 8952 11392 9016 11396
rect 9032 11452 9096 11456
rect 9032 11396 9036 11452
rect 9036 11396 9092 11452
rect 9092 11396 9096 11452
rect 9032 11392 9096 11396
rect 9112 11452 9176 11456
rect 9112 11396 9116 11452
rect 9116 11396 9172 11452
rect 9172 11396 9176 11452
rect 9112 11392 9176 11396
rect 9192 11452 9256 11456
rect 9192 11396 9196 11452
rect 9196 11396 9252 11452
rect 9252 11396 9256 11452
rect 9192 11392 9256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 4952 10908 5016 10912
rect 4952 10852 4956 10908
rect 4956 10852 5012 10908
rect 5012 10852 5016 10908
rect 4952 10848 5016 10852
rect 5032 10908 5096 10912
rect 5032 10852 5036 10908
rect 5036 10852 5092 10908
rect 5092 10852 5096 10908
rect 5032 10848 5096 10852
rect 5112 10908 5176 10912
rect 5112 10852 5116 10908
rect 5116 10852 5172 10908
rect 5172 10852 5176 10908
rect 5112 10848 5176 10852
rect 5192 10908 5256 10912
rect 5192 10852 5196 10908
rect 5196 10852 5252 10908
rect 5252 10852 5256 10908
rect 5192 10848 5256 10852
rect 12952 10908 13016 10912
rect 12952 10852 12956 10908
rect 12956 10852 13012 10908
rect 13012 10852 13016 10908
rect 12952 10848 13016 10852
rect 13032 10908 13096 10912
rect 13032 10852 13036 10908
rect 13036 10852 13092 10908
rect 13092 10852 13096 10908
rect 13032 10848 13096 10852
rect 13112 10908 13176 10912
rect 13112 10852 13116 10908
rect 13116 10852 13172 10908
rect 13172 10852 13176 10908
rect 13112 10848 13176 10852
rect 13192 10908 13256 10912
rect 13192 10852 13196 10908
rect 13196 10852 13252 10908
rect 13252 10852 13256 10908
rect 13192 10848 13256 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 8952 10364 9016 10368
rect 8952 10308 8956 10364
rect 8956 10308 9012 10364
rect 9012 10308 9016 10364
rect 8952 10304 9016 10308
rect 9032 10364 9096 10368
rect 9032 10308 9036 10364
rect 9036 10308 9092 10364
rect 9092 10308 9096 10364
rect 9032 10304 9096 10308
rect 9112 10364 9176 10368
rect 9112 10308 9116 10364
rect 9116 10308 9172 10364
rect 9172 10308 9176 10364
rect 9112 10304 9176 10308
rect 9192 10364 9256 10368
rect 9192 10308 9196 10364
rect 9196 10308 9252 10364
rect 9252 10308 9256 10364
rect 9192 10304 9256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 4952 9820 5016 9824
rect 4952 9764 4956 9820
rect 4956 9764 5012 9820
rect 5012 9764 5016 9820
rect 4952 9760 5016 9764
rect 5032 9820 5096 9824
rect 5032 9764 5036 9820
rect 5036 9764 5092 9820
rect 5092 9764 5096 9820
rect 5032 9760 5096 9764
rect 5112 9820 5176 9824
rect 5112 9764 5116 9820
rect 5116 9764 5172 9820
rect 5172 9764 5176 9820
rect 5112 9760 5176 9764
rect 5192 9820 5256 9824
rect 5192 9764 5196 9820
rect 5196 9764 5252 9820
rect 5252 9764 5256 9820
rect 5192 9760 5256 9764
rect 12952 9820 13016 9824
rect 12952 9764 12956 9820
rect 12956 9764 13012 9820
rect 13012 9764 13016 9820
rect 12952 9760 13016 9764
rect 13032 9820 13096 9824
rect 13032 9764 13036 9820
rect 13036 9764 13092 9820
rect 13092 9764 13096 9820
rect 13032 9760 13096 9764
rect 13112 9820 13176 9824
rect 13112 9764 13116 9820
rect 13116 9764 13172 9820
rect 13172 9764 13176 9820
rect 13112 9760 13176 9764
rect 13192 9820 13256 9824
rect 13192 9764 13196 9820
rect 13196 9764 13252 9820
rect 13252 9764 13256 9820
rect 13192 9760 13256 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 8952 9276 9016 9280
rect 8952 9220 8956 9276
rect 8956 9220 9012 9276
rect 9012 9220 9016 9276
rect 8952 9216 9016 9220
rect 9032 9276 9096 9280
rect 9032 9220 9036 9276
rect 9036 9220 9092 9276
rect 9092 9220 9096 9276
rect 9032 9216 9096 9220
rect 9112 9276 9176 9280
rect 9112 9220 9116 9276
rect 9116 9220 9172 9276
rect 9172 9220 9176 9276
rect 9112 9216 9176 9220
rect 9192 9276 9256 9280
rect 9192 9220 9196 9276
rect 9196 9220 9252 9276
rect 9252 9220 9256 9276
rect 9192 9216 9256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 4952 8732 5016 8736
rect 4952 8676 4956 8732
rect 4956 8676 5012 8732
rect 5012 8676 5016 8732
rect 4952 8672 5016 8676
rect 5032 8732 5096 8736
rect 5032 8676 5036 8732
rect 5036 8676 5092 8732
rect 5092 8676 5096 8732
rect 5032 8672 5096 8676
rect 5112 8732 5176 8736
rect 5112 8676 5116 8732
rect 5116 8676 5172 8732
rect 5172 8676 5176 8732
rect 5112 8672 5176 8676
rect 5192 8732 5256 8736
rect 5192 8676 5196 8732
rect 5196 8676 5252 8732
rect 5252 8676 5256 8732
rect 5192 8672 5256 8676
rect 12952 8732 13016 8736
rect 12952 8676 12956 8732
rect 12956 8676 13012 8732
rect 13012 8676 13016 8732
rect 12952 8672 13016 8676
rect 13032 8732 13096 8736
rect 13032 8676 13036 8732
rect 13036 8676 13092 8732
rect 13092 8676 13096 8732
rect 13032 8672 13096 8676
rect 13112 8732 13176 8736
rect 13112 8676 13116 8732
rect 13116 8676 13172 8732
rect 13172 8676 13176 8732
rect 13112 8672 13176 8676
rect 13192 8732 13256 8736
rect 13192 8676 13196 8732
rect 13196 8676 13252 8732
rect 13252 8676 13256 8732
rect 13192 8672 13256 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 8952 8188 9016 8192
rect 8952 8132 8956 8188
rect 8956 8132 9012 8188
rect 9012 8132 9016 8188
rect 8952 8128 9016 8132
rect 9032 8188 9096 8192
rect 9032 8132 9036 8188
rect 9036 8132 9092 8188
rect 9092 8132 9096 8188
rect 9032 8128 9096 8132
rect 9112 8188 9176 8192
rect 9112 8132 9116 8188
rect 9116 8132 9172 8188
rect 9172 8132 9176 8188
rect 9112 8128 9176 8132
rect 9192 8188 9256 8192
rect 9192 8132 9196 8188
rect 9196 8132 9252 8188
rect 9252 8132 9256 8188
rect 9192 8128 9256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 4952 7644 5016 7648
rect 4952 7588 4956 7644
rect 4956 7588 5012 7644
rect 5012 7588 5016 7644
rect 4952 7584 5016 7588
rect 5032 7644 5096 7648
rect 5032 7588 5036 7644
rect 5036 7588 5092 7644
rect 5092 7588 5096 7644
rect 5032 7584 5096 7588
rect 5112 7644 5176 7648
rect 5112 7588 5116 7644
rect 5116 7588 5172 7644
rect 5172 7588 5176 7644
rect 5112 7584 5176 7588
rect 5192 7644 5256 7648
rect 5192 7588 5196 7644
rect 5196 7588 5252 7644
rect 5252 7588 5256 7644
rect 5192 7584 5256 7588
rect 12952 7644 13016 7648
rect 12952 7588 12956 7644
rect 12956 7588 13012 7644
rect 13012 7588 13016 7644
rect 12952 7584 13016 7588
rect 13032 7644 13096 7648
rect 13032 7588 13036 7644
rect 13036 7588 13092 7644
rect 13092 7588 13096 7644
rect 13032 7584 13096 7588
rect 13112 7644 13176 7648
rect 13112 7588 13116 7644
rect 13116 7588 13172 7644
rect 13172 7588 13176 7644
rect 13112 7584 13176 7588
rect 13192 7644 13256 7648
rect 13192 7588 13196 7644
rect 13196 7588 13252 7644
rect 13252 7588 13256 7644
rect 13192 7584 13256 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 8952 7100 9016 7104
rect 8952 7044 8956 7100
rect 8956 7044 9012 7100
rect 9012 7044 9016 7100
rect 8952 7040 9016 7044
rect 9032 7100 9096 7104
rect 9032 7044 9036 7100
rect 9036 7044 9092 7100
rect 9092 7044 9096 7100
rect 9032 7040 9096 7044
rect 9112 7100 9176 7104
rect 9112 7044 9116 7100
rect 9116 7044 9172 7100
rect 9172 7044 9176 7100
rect 9112 7040 9176 7044
rect 9192 7100 9256 7104
rect 9192 7044 9196 7100
rect 9196 7044 9252 7100
rect 9252 7044 9256 7100
rect 9192 7040 9256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 4952 6556 5016 6560
rect 4952 6500 4956 6556
rect 4956 6500 5012 6556
rect 5012 6500 5016 6556
rect 4952 6496 5016 6500
rect 5032 6556 5096 6560
rect 5032 6500 5036 6556
rect 5036 6500 5092 6556
rect 5092 6500 5096 6556
rect 5032 6496 5096 6500
rect 5112 6556 5176 6560
rect 5112 6500 5116 6556
rect 5116 6500 5172 6556
rect 5172 6500 5176 6556
rect 5112 6496 5176 6500
rect 5192 6556 5256 6560
rect 5192 6500 5196 6556
rect 5196 6500 5252 6556
rect 5252 6500 5256 6556
rect 5192 6496 5256 6500
rect 12952 6556 13016 6560
rect 12952 6500 12956 6556
rect 12956 6500 13012 6556
rect 13012 6500 13016 6556
rect 12952 6496 13016 6500
rect 13032 6556 13096 6560
rect 13032 6500 13036 6556
rect 13036 6500 13092 6556
rect 13092 6500 13096 6556
rect 13032 6496 13096 6500
rect 13112 6556 13176 6560
rect 13112 6500 13116 6556
rect 13116 6500 13172 6556
rect 13172 6500 13176 6556
rect 13112 6496 13176 6500
rect 13192 6556 13256 6560
rect 13192 6500 13196 6556
rect 13196 6500 13252 6556
rect 13252 6500 13256 6556
rect 13192 6496 13256 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 8952 6012 9016 6016
rect 8952 5956 8956 6012
rect 8956 5956 9012 6012
rect 9012 5956 9016 6012
rect 8952 5952 9016 5956
rect 9032 6012 9096 6016
rect 9032 5956 9036 6012
rect 9036 5956 9092 6012
rect 9092 5956 9096 6012
rect 9032 5952 9096 5956
rect 9112 6012 9176 6016
rect 9112 5956 9116 6012
rect 9116 5956 9172 6012
rect 9172 5956 9176 6012
rect 9112 5952 9176 5956
rect 9192 6012 9256 6016
rect 9192 5956 9196 6012
rect 9196 5956 9252 6012
rect 9252 5956 9256 6012
rect 9192 5952 9256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 4952 5468 5016 5472
rect 4952 5412 4956 5468
rect 4956 5412 5012 5468
rect 5012 5412 5016 5468
rect 4952 5408 5016 5412
rect 5032 5468 5096 5472
rect 5032 5412 5036 5468
rect 5036 5412 5092 5468
rect 5092 5412 5096 5468
rect 5032 5408 5096 5412
rect 5112 5468 5176 5472
rect 5112 5412 5116 5468
rect 5116 5412 5172 5468
rect 5172 5412 5176 5468
rect 5112 5408 5176 5412
rect 5192 5468 5256 5472
rect 5192 5412 5196 5468
rect 5196 5412 5252 5468
rect 5252 5412 5256 5468
rect 5192 5408 5256 5412
rect 12952 5468 13016 5472
rect 12952 5412 12956 5468
rect 12956 5412 13012 5468
rect 13012 5412 13016 5468
rect 12952 5408 13016 5412
rect 13032 5468 13096 5472
rect 13032 5412 13036 5468
rect 13036 5412 13092 5468
rect 13092 5412 13096 5468
rect 13032 5408 13096 5412
rect 13112 5468 13176 5472
rect 13112 5412 13116 5468
rect 13116 5412 13172 5468
rect 13172 5412 13176 5468
rect 13112 5408 13176 5412
rect 13192 5468 13256 5472
rect 13192 5412 13196 5468
rect 13196 5412 13252 5468
rect 13252 5412 13256 5468
rect 13192 5408 13256 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 8952 4924 9016 4928
rect 8952 4868 8956 4924
rect 8956 4868 9012 4924
rect 9012 4868 9016 4924
rect 8952 4864 9016 4868
rect 9032 4924 9096 4928
rect 9032 4868 9036 4924
rect 9036 4868 9092 4924
rect 9092 4868 9096 4924
rect 9032 4864 9096 4868
rect 9112 4924 9176 4928
rect 9112 4868 9116 4924
rect 9116 4868 9172 4924
rect 9172 4868 9176 4924
rect 9112 4864 9176 4868
rect 9192 4924 9256 4928
rect 9192 4868 9196 4924
rect 9196 4868 9252 4924
rect 9252 4868 9256 4924
rect 9192 4864 9256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 4952 4380 5016 4384
rect 4952 4324 4956 4380
rect 4956 4324 5012 4380
rect 5012 4324 5016 4380
rect 4952 4320 5016 4324
rect 5032 4380 5096 4384
rect 5032 4324 5036 4380
rect 5036 4324 5092 4380
rect 5092 4324 5096 4380
rect 5032 4320 5096 4324
rect 5112 4380 5176 4384
rect 5112 4324 5116 4380
rect 5116 4324 5172 4380
rect 5172 4324 5176 4380
rect 5112 4320 5176 4324
rect 5192 4380 5256 4384
rect 5192 4324 5196 4380
rect 5196 4324 5252 4380
rect 5252 4324 5256 4380
rect 5192 4320 5256 4324
rect 12952 4380 13016 4384
rect 12952 4324 12956 4380
rect 12956 4324 13012 4380
rect 13012 4324 13016 4380
rect 12952 4320 13016 4324
rect 13032 4380 13096 4384
rect 13032 4324 13036 4380
rect 13036 4324 13092 4380
rect 13092 4324 13096 4380
rect 13032 4320 13096 4324
rect 13112 4380 13176 4384
rect 13112 4324 13116 4380
rect 13116 4324 13172 4380
rect 13172 4324 13176 4380
rect 13112 4320 13176 4324
rect 13192 4380 13256 4384
rect 13192 4324 13196 4380
rect 13196 4324 13252 4380
rect 13252 4324 13256 4380
rect 13192 4320 13256 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 8952 3836 9016 3840
rect 8952 3780 8956 3836
rect 8956 3780 9012 3836
rect 9012 3780 9016 3836
rect 8952 3776 9016 3780
rect 9032 3836 9096 3840
rect 9032 3780 9036 3836
rect 9036 3780 9092 3836
rect 9092 3780 9096 3836
rect 9032 3776 9096 3780
rect 9112 3836 9176 3840
rect 9112 3780 9116 3836
rect 9116 3780 9172 3836
rect 9172 3780 9176 3836
rect 9112 3776 9176 3780
rect 9192 3836 9256 3840
rect 9192 3780 9196 3836
rect 9196 3780 9252 3836
rect 9252 3780 9256 3836
rect 9192 3776 9256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 4952 3292 5016 3296
rect 4952 3236 4956 3292
rect 4956 3236 5012 3292
rect 5012 3236 5016 3292
rect 4952 3232 5016 3236
rect 5032 3292 5096 3296
rect 5032 3236 5036 3292
rect 5036 3236 5092 3292
rect 5092 3236 5096 3292
rect 5032 3232 5096 3236
rect 5112 3292 5176 3296
rect 5112 3236 5116 3292
rect 5116 3236 5172 3292
rect 5172 3236 5176 3292
rect 5112 3232 5176 3236
rect 5192 3292 5256 3296
rect 5192 3236 5196 3292
rect 5196 3236 5252 3292
rect 5252 3236 5256 3292
rect 5192 3232 5256 3236
rect 12952 3292 13016 3296
rect 12952 3236 12956 3292
rect 12956 3236 13012 3292
rect 13012 3236 13016 3292
rect 12952 3232 13016 3236
rect 13032 3292 13096 3296
rect 13032 3236 13036 3292
rect 13036 3236 13092 3292
rect 13092 3236 13096 3292
rect 13032 3232 13096 3236
rect 13112 3292 13176 3296
rect 13112 3236 13116 3292
rect 13116 3236 13172 3292
rect 13172 3236 13176 3292
rect 13112 3232 13176 3236
rect 13192 3292 13256 3296
rect 13192 3236 13196 3292
rect 13196 3236 13252 3292
rect 13252 3236 13256 3292
rect 13192 3232 13256 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 8952 2748 9016 2752
rect 8952 2692 8956 2748
rect 8956 2692 9012 2748
rect 9012 2692 9016 2748
rect 8952 2688 9016 2692
rect 9032 2748 9096 2752
rect 9032 2692 9036 2748
rect 9036 2692 9092 2748
rect 9092 2692 9096 2748
rect 9032 2688 9096 2692
rect 9112 2748 9176 2752
rect 9112 2692 9116 2748
rect 9116 2692 9172 2748
rect 9172 2692 9176 2748
rect 9112 2688 9176 2692
rect 9192 2748 9256 2752
rect 9192 2692 9196 2748
rect 9196 2692 9252 2748
rect 9252 2692 9256 2748
rect 9192 2688 9256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 4952 2204 5016 2208
rect 4952 2148 4956 2204
rect 4956 2148 5012 2204
rect 5012 2148 5016 2204
rect 4952 2144 5016 2148
rect 5032 2204 5096 2208
rect 5032 2148 5036 2204
rect 5036 2148 5092 2204
rect 5092 2148 5096 2204
rect 5032 2144 5096 2148
rect 5112 2204 5176 2208
rect 5112 2148 5116 2204
rect 5116 2148 5172 2204
rect 5172 2148 5176 2204
rect 5112 2144 5176 2148
rect 5192 2204 5256 2208
rect 5192 2148 5196 2204
rect 5196 2148 5252 2204
rect 5252 2148 5256 2204
rect 5192 2144 5256 2148
rect 12952 2204 13016 2208
rect 12952 2148 12956 2204
rect 12956 2148 13012 2204
rect 13012 2148 13016 2204
rect 12952 2144 13016 2148
rect 13032 2204 13096 2208
rect 13032 2148 13036 2204
rect 13036 2148 13092 2204
rect 13092 2148 13096 2204
rect 13032 2144 13096 2148
rect 13112 2204 13176 2208
rect 13112 2148 13116 2204
rect 13116 2148 13172 2204
rect 13172 2148 13176 2204
rect 13112 2144 13176 2148
rect 13192 2204 13256 2208
rect 13192 2148 13196 2204
rect 13196 2148 13252 2204
rect 13252 2148 13256 2204
rect 13192 2144 13256 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
<< metal4 >>
rect 4944 21792 5264 21808
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 20704 5264 21728
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 19616 5264 20640
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 18528 5264 19552
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 17440 5264 18464
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 59 16420 125 16421
rect 59 16356 60 16420
rect 124 16356 125 16420
rect 59 16355 125 16356
rect 62 16149 122 16355
rect 4944 16352 5264 17376
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 59 16148 125 16149
rect 59 16084 60 16148
rect 124 16084 125 16148
rect 59 16083 125 16084
rect 4944 15264 5264 16288
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 14176 5264 15200
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 13088 5264 14112
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 12000 5264 13024
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 10912 5264 11936
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 9824 5264 10848
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 8736 5264 9760
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 7648 5264 8672
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 6560 5264 7584
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 5472 5264 6496
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 4384 5264 5408
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 3296 5264 4320
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 2208 5264 3232
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2128 5264 2144
rect 8944 21248 9264 21808
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 20160 9264 21184
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 19072 9264 20096
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 17984 9264 19008
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 16896 9264 17920
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 15808 9264 16832
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 14720 9264 15744
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 13632 9264 14656
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 12544 9264 13568
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 11456 9264 12480
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 10368 9264 11392
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 9280 9264 10304
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 8192 9264 9216
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 7104 9264 8128
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 6016 9264 7040
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 4928 9264 5952
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 3840 9264 4864
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 2752 9264 3776
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2128 9264 2688
rect 12944 21792 13264 21808
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 20704 13264 21728
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 19616 13264 20640
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 18528 13264 19552
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 17440 13264 18464
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 16352 13264 17376
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 15264 13264 16288
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 14176 13264 15200
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 13088 13264 14112
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 12000 13264 13024
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 10912 13264 11936
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 9824 13264 10848
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 8736 13264 9760
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 7648 13264 8672
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 6560 13264 7584
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 5472 13264 6496
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 4384 13264 5408
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 3296 13264 4320
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 2208 13264 3232
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2128 13264 2144
rect 16944 21248 17264 21808
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 17984 17264 19008
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 12544 17264 13568
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8192 17264 9216
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 7104 17264 8128
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 2752 17264 3776
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2128 17264 2688
rect 20944 21792 21264 21808
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 20704 21264 21728
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 19616 21264 20640
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 18528 21264 19552
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 17440 21264 18464
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 16352 21264 17376
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 15264 21264 16288
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 14176 21264 15200
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 13088 21264 14112
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
use scs8hd_fill_2  FILLER_1_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_10
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_10 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_22 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3128 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_17
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_21
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 774 592
use scs8hd_inv_8  _112_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_30 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_32 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_38
timestamp 1586364061
transform 1 0 4600 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_29
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 314 592
use scs8hd_inv_8  _083_
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_42
timestamp 1586364061
transform 1 0 4968 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_43
timestamp 1586364061
transform 1 0 5060 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_47
timestamp 1586364061
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use scs8hd_or2_4  _122_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 682 592
use scs8hd_nand2_4  _126_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_69
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _204_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_1_73
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_79
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 406 592
use scs8hd_inv_8  _094_
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_94
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_115
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_111
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_111
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_119
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _093_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_140
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_149
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_149 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 314 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_160
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_164
timestamp 1586364061
transform 1 0 16192 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_166
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 17112 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_172
timestamp 1586364061
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_176
timestamp 1586364061
transform 1 0 17296 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_170
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_184
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_182
timestamp 1586364061
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_190
timestamp 1586364061
transform 1 0 18584 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19964 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_194
timestamp 1586364061
transform 1 0 18952 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_206
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_212
timestamp 1586364061
transform 1 0 20608 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_221
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_218
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 22816 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 22816 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_225
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_1_230
timestamp 1586364061
transform 1 0 22264 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_11
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 130 592
use scs8hd_conb_1  _186_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_14
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_18
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_30
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_45
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_57
timestamp 1586364061
transform 1 0 6348 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_61
timestamp 1586364061
transform 1 0 6716 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_75
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_104
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_108
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_121
timestamp 1586364061
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_133
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_152
timestamp 1586364061
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 15548 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use scs8hd_conb_1  _191_
timestamp 1586364061
transform 1 0 17296 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_168
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_172
timestamp 1586364061
transform 1 0 16928 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_179
timestamp 1586364061
transform 1 0 17572 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_191
timestamp 1586364061
transform 1 0 18676 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 22816 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_16
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_20
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_26
timestamp 1586364061
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3864 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_43
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_65
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_69
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 774 592
use scs8hd_nor2_4  _138_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_94
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_3_109
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_113
timestamp 1586364061
transform 1 0 11500 0 1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_3_121
timestamp 1586364061
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_conb_1  _184_
timestamp 1586364061
transform 1 0 12880 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_131
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 866 592
use scs8hd_decap_4  FILLER_3_149
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_153
timestamp 1586364061
transform 1 0 15180 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_inv_8  _102_
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_200
timestamp 1586364061
transform 1 0 19504 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_212
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_217
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_221
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 22816 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  FILLER_4_9
timestamp 1586364061
transform 1 0 1932 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_21
timestamp 1586364061
transform 1 0 3036 0 -1 4896
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _080_
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_43
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__D
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_60
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_64
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_73
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_83
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use scs8hd_conb_1  _195_
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_113
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_4  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_139
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_151
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_165
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 17388 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_169
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_198
timestamp 1586364061
transform 1 0 19320 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 22816 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_232
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_21
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_26
timestamp 1586364061
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 3680 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 5888 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_43
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_50
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_54
timestamp 1586364061
transform 1 0 6072 0 1 4896
box -38 -48 406 592
use scs8hd_or4_4  _173_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_58
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__D
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_79
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_82
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_or4_4  _136_
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 406 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_101
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_142
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_146
timestamp 1586364061
transform 1 0 14536 0 1 4896
box -38 -48 1142 592
use scs8hd_inv_8  _108_
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_158
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_170
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18308 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_180
timestamp 1586364061
transform 1 0 17664 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20056 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_198
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_215
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_219
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 22816 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_231
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _111_
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_16
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_19
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_20
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 3128 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_24
timestamp 1586364061
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_24
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_37
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 314 592
use scs8hd_or2_4  _121_
timestamp 1586364061
transform 1 0 5336 0 1 5984
box -38 -48 682 592
use scs8hd_nand2_4  _148_
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_48
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_42
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_59
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__173__C
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__C
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_64
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use scs8hd_nor3_4  _177_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 1 5984
box -38 -48 1234 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_82
timestamp 1586364061
transform 1 0 8648 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_76
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_80
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__C
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_94
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _081_
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_115
timestamp 1586364061
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_111
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_115
timestamp 1586364061
transform 1 0 11684 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__D
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 11868 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_119
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_119
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 1050 592
use scs8hd_inv_8  _107_
timestamp 1586364061
transform 1 0 12972 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__158__C
timestamp 1586364061
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_134
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_138
timestamp 1586364061
transform 1 0 13800 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_127
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_7_142
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_161
timestamp 1586364061
transform 1 0 15916 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_166
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_175
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_173
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_177
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18768 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_189
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_190
timestamp 1586364061
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_201
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_194
timestamp 1586364061
transform 1 0 18952 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_202
timestamp 1586364061
transform 1 0 19688 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_207
timestamp 1586364061
transform 1 0 20148 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20332 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_208
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_218
timestamp 1586364061
transform 1 0 21160 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 22816 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 22816 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_230
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_224
timestamp 1586364061
transform 1 0 21712 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 130 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3128 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_16
timestamp 1586364061
transform 1 0 2576 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_20
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_24
timestamp 1586364061
transform 1 0 3312 0 -1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 3680 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_30
timestamp 1586364061
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use scs8hd_or4_4  _164_
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_46
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_69
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_8  _120_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use scs8hd_or4_4  _158_
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_8  _087_
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_139
timestamp 1586364061
transform 1 0 13892 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_8_151
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_162
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_173
timestamp 1586364061
transform 1 0 17020 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_181
timestamp 1586364061
transform 1 0 17756 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_199
timestamp 1586364061
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_211
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 22816 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_232
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_14
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_18
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__D
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_33
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_37
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_40
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_or4_4  _167_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__D
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _179_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__176__C
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__C
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_65
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_69
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_73
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_92
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_96
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 314 592
use scs8hd_or4_4  _127_
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__D
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_101
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 590 592
use scs8hd_nor2_4  _160_
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 866 592
use scs8hd_decap_4  FILLER_9_149
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_168
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 1142 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 774 592
use scs8hd_inv_8  _088_
timestamp 1586364061
transform 1 0 20056 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_201
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_215
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_219
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 22816 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_231
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_20
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_25
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_35
timestamp 1586364061
transform 1 0 4324 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_39
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_8  _103_
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 4968 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_53
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 774 592
use scs8hd_nor3_4  _176_
timestamp 1586364061
transform 1 0 6900 0 -1 8160
box -38 -48 1234 592
use scs8hd_fill_2  FILLER_10_61
timestamp 1586364061
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_82
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_8  _119_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_85
timestamp 1586364061
transform 1 0 8924 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_107
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12512 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_10_119
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_123
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_135
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_139
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_142
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_146
timestamp 1586364061
transform 1 0 14536 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_157
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_161
timestamp 1586364061
transform 1 0 15916 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_173
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_185
timestamp 1586364061
transform 1 0 18124 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_197
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_209
timestamp 1586364061
transform 1 0 20332 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_218
timestamp 1586364061
transform 1 0 21160 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 22816 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_230
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_83
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_87
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _182_
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_100
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_104
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 406 592
use scs8hd_conb_1  _192_
timestamp 1586364061
transform 1 0 12512 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11868 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_111
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 590 592
use scs8hd_decap_3  FILLER_11_119
timestamp 1586364061
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_127
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_133
timestamp 1586364061
transform 1 0 13340 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_144
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_148
timestamp 1586364061
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_152
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_166
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_170
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_182
timestamp 1586364061
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_214
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_218
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 22816 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21712 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_222
timestamp 1586364061
transform 1 0 21528 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_226
timestamp 1586364061
transform 1 0 21896 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_17
timestamp 1586364061
transform 1 0 2668 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_29
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_40
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5520 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_46
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use scs8hd_conb_1  _178_
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_57
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 406 592
use scs8hd_conb_1  _181_
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_74
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_6  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 590 592
use scs8hd_inv_8  _084_
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_12_99
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_109
timestamp 1586364061
transform 1 0 11132 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_120
timestamp 1586364061
transform 1 0 12144 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_12_128
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_12_150
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15548 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_168
timestamp 1586364061
transform 1 0 16560 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_12_176
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_184
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_188
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_200
timestamp 1586364061
transform 1 0 19504 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_208
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_212
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_218
timestamp 1586364061
transform 1 0 21160 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 22816 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_230
timestamp 1586364061
transform 1 0 22264 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_9
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_9
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _114_
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 3496 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_22
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_26
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_20
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_24
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_28
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_30
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 1050 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__D
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__C
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_43
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_47
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_54
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_62
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_58
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__D
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__C
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_conb_1  _180_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_69
timestamp 1586364061
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_65
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__C
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use scs8hd_nor3_4  _174_
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 1234 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_73
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_77
timestamp 1586364061
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_81
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_8  _117_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__D
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_88
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_93
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_85
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_89
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_8  _082_
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use scs8hd_or4_4  _145_
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__C
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 590 592
use scs8hd_decap_4  FILLER_14_119
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _146_
timestamp 1586364061
transform 1 0 13156 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_133
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_144
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use scs8hd_inv_8  _099_
timestamp 1586364061
transform 1 0 15364 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_163
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_164
timestamp 1586364061
transform 1 0 16192 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 866 592
use scs8hd_conb_1  _190_
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_176
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_172
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_180
timestamp 1586364061
transform 1 0 17664 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_183
timestamp 1586364061
transform 1 0 17940 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_205
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_195
timestamp 1586364061
transform 1 0 19044 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_207
timestamp 1586364061
transform 1 0 20148 0 -1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_219
timestamp 1586364061
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 22816 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 22816 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_223
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_227
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_232
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_inv_8  _115_
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_18
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_22
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_35
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 314 592
use scs8hd_or4_4  _152_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_68
timestamp 1586364061
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_83
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_87
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__C
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_100
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_105
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_109
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_or4_4  _161_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_15_149
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 406 592
use scs8hd_conb_1  _185_
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_153
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_172
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_176
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_180
timestamp 1586364061
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_inv_8  _100_
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_202
timestamp 1586364061
transform 1 0 19688 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_214
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 22816 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_225
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_16
timestamp 1586364061
transform 1 0 2576 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_20
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _171_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_28
timestamp 1586364061
transform 1 0 3680 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use scs8hd_or4_4  _142_
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_61
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_70
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_74
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_16_96
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 222 592
use scs8hd_or4_4  _133_
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 10120 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__C
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_100
timestamp 1586364061
transform 1 0 10304 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_104
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__161__D
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__D
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_116
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_120
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _163_
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  FILLER_16_171
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_183
timestamp 1586364061
transform 1 0 17940 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_189
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_201
timestamp 1586364061
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 22816 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_6
timestamp 1586364061
transform 1 0 1656 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_10
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2668 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_14
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_28
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 406 592
use scs8hd_decap_4  FILLER_17_34
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_40
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_nor3_4  _175_
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__C
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_77
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_87
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_91
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _139_
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__D
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_116
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_120
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _109_
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 13340 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_127
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_131
timestamp 1586364061
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_144
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_148
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_161
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_165
timestamp 1586364061
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_169
timestamp 1586364061
transform 1 0 16652 0 1 11424
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_198
timestamp 1586364061
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_202
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_210
timestamp 1586364061
transform 1 0 20424 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_218
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 22816 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_222
timestamp 1586364061
transform 1 0 21528 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_226
timestamp 1586364061
transform 1 0 21896 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2668 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_14
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_19
timestamp 1586364061
transform 1 0 2852 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _170_
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_43
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_47
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__170__D
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_60
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_71
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_18_83
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _155_
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__139__D
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 774 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_127
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_131
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_135
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_169
timestamp 1586364061
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_173
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18308 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_185
timestamp 1586364061
transform 1 0 18124 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_189
timestamp 1586364061
transform 1 0 18492 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_8  _110_
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_211
timestamp 1586364061
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 22816 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_232
timestamp 1586364061
transform 1 0 22448 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_8  _116_
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_18
timestamp 1586364061
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_14
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_18
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_14
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2576 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_26
timestamp 1586364061
transform 1 0 3496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_22
timestamp 1586364061
transform 1 0 3128 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_22
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _172_
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_29
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5888 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_46
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_65
timestamp 1586364061
transform 1 0 7084 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_69
timestamp 1586364061
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_73
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_97
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_101
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_107
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_138
timestamp 1586364061
transform 1 0 13800 0 -1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_140
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_142
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_151
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_8  _105_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_8  _106_
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_154
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_158
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 590 592
use scs8hd_decap_3  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_192
timestamp 1586364061
transform 1 0 18768 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_204
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_204
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20332 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_218
timestamp 1586364061
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_212
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 22816 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 22816 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_19_222
timestamp 1586364061
transform 1 0 21528 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_230
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_17
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_21
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_25
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 6072 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5704 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_44
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_48
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_52
timestamp 1586364061
transform 1 0 5888 0 1 13600
box -38 -48 222 592
use scs8hd_inv_8  _098_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_56
timestamp 1586364061
transform 1 0 6256 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_60
timestamp 1586364061
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_21_83
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 1142 592
use scs8hd_conb_1  _188_
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_136
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_144
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_158
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_162
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 22816 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_16
timestamp 1586364061
transform 1 0 2576 0 -1 14688
box -38 -48 1142 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_28
timestamp 1586364061
transform 1 0 3680 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_40
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_71
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_8  _096_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_87
timestamp 1586364061
transform 1 0 9108 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_90
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_110
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_121
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_8  FILLER_22_134
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 774 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_151
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_175
timestamp 1586364061
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_187
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_199
timestamp 1586364061
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_211
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 22816 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 590 592
use scs8hd_inv_8  _104_
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_16
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_20
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_24
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_29
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_42
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_46
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_23_49
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 1142 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_85
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_101
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_105
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 590 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_111
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 1142 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_148
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_152
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_163
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 22816 0 1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_6
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_10
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4692 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_38
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 590 592
use scs8hd_inv_8  _097_
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 590 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_73
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_24_108
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12144 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_131
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_147
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 22816 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 590 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_30
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_50
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_54
timestamp 1586364061
transform 1 0 6072 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_58
timestamp 1586364061
transform 1 0 6440 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_73
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_77
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_81
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_85
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_88
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_103
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_107
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12512 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_115
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _092_
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_139
timestamp 1586364061
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_152
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_164
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_25_176
timestamp 1586364061
transform 1 0 17296 0 1 15776
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_182
timestamp 1586364061
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_214
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_217
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 22816 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_25_229
timestamp 1586364061
transform 1 0 22172 0 1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_6
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_6
timestamp 1586364061
transform 1 0 1656 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_10
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_14
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_25
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_29
timestamp 1586364061
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_33
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_37
timestamp 1586364061
transform 1 0 4508 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_40
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _086_
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_54
timestamp 1586364061
transform 1 0 6072 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_62
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_66
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_65
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 314 592
use scs8hd_inv_8  _118_
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_70
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_83
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_87
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_91
timestamp 1586364061
transform 1 0 9476 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_94
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_118
timestamp 1586364061
transform 1 0 11960 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_124
timestamp 1586364061
transform 1 0 12512 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_111
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_27_116
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 590 592
use scs8hd_decap_6  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_134
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_138
timestamp 1586364061
transform 1 0 13800 0 -1 16864
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_140
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_144
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_152
timestamp 1586364061
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_156
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_168
timestamp 1586364061
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_180
timestamp 1586364061
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_218
timestamp 1586364061
transform 1 0 21160 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_214
timestamp 1586364061
transform 1 0 20792 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_217
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 22816 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 22816 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_230
timestamp 1586364061
transform 1 0 22264 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_229
timestamp 1586364061
transform 1 0 22172 0 1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_6
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_8  _085_
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5520 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_46
timestamp 1586364061
transform 1 0 5336 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_57
timestamp 1586364061
transform 1 0 6348 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_82
timestamp 1586364061
transform 1 0 8648 0 -1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_90
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 11592 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_123
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_133
timestamp 1586364061
transform 1 0 13340 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_143
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_151
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_157
timestamp 1586364061
transform 1 0 15548 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_169
timestamp 1586364061
transform 1 0 16652 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_181
timestamp 1586364061
transform 1 0 17756 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_193
timestamp 1586364061
transform 1 0 18860 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_205
timestamp 1586364061
transform 1 0 19964 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_213
timestamp 1586364061
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_218
timestamp 1586364061
transform 1 0 21160 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 22816 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_230
timestamp 1586364061
transform 1 0 22264 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_6
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_10
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_14
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_26
timestamp 1586364061
transform 1 0 3496 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_65
timestamp 1586364061
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_69
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__213__A
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_73
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_87
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _194_
timestamp 1586364061
transform 1 0 12512 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_127
timestamp 1586364061
transform 1 0 12788 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_131
timestamp 1586364061
transform 1 0 13156 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_144
timestamp 1586364061
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_148
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_155
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_214
timestamp 1586364061
transform 1 0 20792 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_217
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 22816 0 1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_29_229
timestamp 1586364061
transform 1 0 22172 0 1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_18
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_buf_2  _213_
timestamp 1586364061
transform 1 0 6900 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_6  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_62
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_67
timestamp 1586364061
transform 1 0 7268 0 -1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_75
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use scs8hd_conb_1  _193_
timestamp 1586364061
transform 1 0 10028 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_100
timestamp 1586364061
transform 1 0 10304 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_104
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_8  _091_
timestamp 1586364061
transform 1 0 13340 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_4  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_8  FILLER_30_142
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_150
timestamp 1586364061
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_218
timestamp 1586364061
transform 1 0 21160 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 22816 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_230
timestamp 1586364061
transform 1 0 22264 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_19
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_31
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_43
timestamp 1586364061
transform 1 0 5060 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_31_55
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8280 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_31_80
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_92
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 774 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 10672 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 10488 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_100
timestamp 1586364061
transform 1 0 10304 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_113
timestamp 1586364061
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_117
timestamp 1586364061
transform 1 0 11868 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 590 592
use scs8hd_buf_2  _210_
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_141
timestamp 1586364061
transform 1 0 14076 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_146
timestamp 1586364061
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_150
timestamp 1586364061
transform 1 0 14904 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_162
timestamp 1586364061
transform 1 0 16008 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_174
timestamp 1586364061
transform 1 0 17112 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_182
timestamp 1586364061
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 22816 0 1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_18
timestamp 1586364061
transform 1 0 2760 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_30
timestamp 1586364061
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_76
timestamp 1586364061
transform 1 0 8096 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_81
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_89
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_114
timestamp 1586364061
transform 1 0 11592 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_126
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_138
timestamp 1586364061
transform 1 0 13800 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_32_150
timestamp 1586364061
transform 1 0 14904 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 22816 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 590 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_11
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 3772 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_31
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_43
timestamp 1586364061
transform 1 0 5060 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_49
timestamp 1586364061
transform 1 0 5612 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _212_
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__212__A
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_106
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_109
timestamp 1586364061
transform 1 0 11132 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _211_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_121
timestamp 1586364061
transform 1 0 12236 0 -1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__211__A
timestamp 1586364061
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_127
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_131
timestamp 1586364061
transform 1 0 13156 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_133
timestamp 1586364061
transform 1 0 13340 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_143
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_155
timestamp 1586364061
transform 1 0 15364 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_167
timestamp 1586364061
transform 1 0 16468 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_173
timestamp 1586364061
transform 1 0 17020 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_177
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20516 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20976 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_214
timestamp 1586364061
transform 1 0 20792 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_218
timestamp 1586364061
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21528 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 22816 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 22816 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_225
timestamp 1586364061
transform 1 0 21804 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_229
timestamp 1586364061
transform 1 0 22172 0 1 20128
box -38 -48 406 592
use scs8hd_decap_6  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_63
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_125
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_137
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 22816 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 314 592
<< labels >>
rlabel metal3 s 23520 688 24000 808 6 address[0]
port 0 nsew default input
rlabel metal3 s 23520 2048 24000 2168 6 address[1]
port 1 nsew default input
rlabel metal3 s 23520 3408 24000 3528 6 address[2]
port 2 nsew default input
rlabel metal3 s 0 552 480 672 6 address[3]
port 3 nsew default input
rlabel metal2 s 3882 0 3938 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 5538 0 5594 480 6 address[5]
port 5 nsew default input
rlabel metal3 s 23520 4904 24000 5024 6 chanx_right_in[0]
port 6 nsew default input
rlabel metal3 s 0 1640 480 1760 6 chanx_right_in[1]
port 7 nsew default input
rlabel metal3 s 23520 6264 24000 6384 6 chanx_right_in[2]
port 8 nsew default input
rlabel metal3 s 23520 7624 24000 7744 6 chanx_right_in[3]
port 9 nsew default input
rlabel metal3 s 0 2864 480 2984 6 chanx_right_in[4]
port 10 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chanx_right_in[5]
port 11 nsew default input
rlabel metal2 s 8758 0 8814 480 6 chanx_right_in[6]
port 12 nsew default input
rlabel metal3 s 23520 9120 24000 9240 6 chanx_right_in[7]
port 13 nsew default input
rlabel metal3 s 23520 10480 24000 10600 6 chanx_right_in[8]
port 14 nsew default input
rlabel metal2 s 10322 0 10378 480 6 chanx_right_out[0]
port 15 nsew default tristate
rlabel metal2 s 1214 23520 1270 24000 6 chanx_right_out[1]
port 16 nsew default tristate
rlabel metal3 s 0 4088 480 4208 6 chanx_right_out[2]
port 17 nsew default tristate
rlabel metal2 s 11886 0 11942 480 6 chanx_right_out[3]
port 18 nsew default tristate
rlabel metal3 s 0 5312 480 5432 6 chanx_right_out[4]
port 19 nsew default tristate
rlabel metal3 s 0 6536 480 6656 6 chanx_right_out[5]
port 20 nsew default tristate
rlabel metal3 s 0 7624 480 7744 6 chanx_right_out[6]
port 21 nsew default tristate
rlabel metal3 s 0 8848 480 8968 6 chanx_right_out[7]
port 22 nsew default tristate
rlabel metal2 s 3606 23520 3662 24000 6 chanx_right_out[8]
port 23 nsew default tristate
rlabel metal3 s 23520 11840 24000 11960 6 chany_top_in[0]
port 24 nsew default input
rlabel metal3 s 23520 13336 24000 13456 6 chany_top_in[1]
port 25 nsew default input
rlabel metal3 s 23520 14696 24000 14816 6 chany_top_in[2]
port 26 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chany_top_in[3]
port 27 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chany_top_in[4]
port 28 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chany_top_in[5]
port 29 nsew default input
rlabel metal2 s 5998 23520 6054 24000 6 chany_top_in[6]
port 30 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chany_top_in[7]
port 31 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chany_top_in[8]
port 32 nsew default input
rlabel metal2 s 8390 23520 8446 24000 6 chany_top_out[0]
port 33 nsew default tristate
rlabel metal2 s 10782 23520 10838 24000 6 chany_top_out[1]
port 34 nsew default tristate
rlabel metal2 s 13174 23520 13230 24000 6 chany_top_out[2]
port 35 nsew default tristate
rlabel metal2 s 15566 23520 15622 24000 6 chany_top_out[3]
port 36 nsew default tristate
rlabel metal2 s 13542 0 13598 480 6 chany_top_out[4]
port 37 nsew default tristate
rlabel metal3 s 23520 16056 24000 16176 6 chany_top_out[5]
port 38 nsew default tristate
rlabel metal3 s 0 16056 480 16176 6 chany_top_out[6]
port 39 nsew default tristate
rlabel metal2 s 15106 0 15162 480 6 chany_top_out[7]
port 40 nsew default tristate
rlabel metal2 s 16762 0 16818 480 6 chany_top_out[8]
port 41 nsew default tristate
rlabel metal2 s 2318 0 2374 480 6 data_in
port 42 nsew default input
rlabel metal2 s 754 0 810 480 6 enable
port 43 nsew default input
rlabel metal3 s 0 17280 480 17400 6 right_bottom_grid_pin_11_
port 44 nsew default input
rlabel metal3 s 23520 20272 24000 20392 6 right_bottom_grid_pin_13_
port 45 nsew default input
rlabel metal2 s 21546 0 21602 480 6 right_bottom_grid_pin_15_
port 46 nsew default input
rlabel metal2 s 17958 23520 18014 24000 6 right_bottom_grid_pin_1_
port 47 nsew default input
rlabel metal2 s 18326 0 18382 480 6 right_bottom_grid_pin_3_
port 48 nsew default input
rlabel metal3 s 23520 17552 24000 17672 6 right_bottom_grid_pin_5_
port 49 nsew default input
rlabel metal2 s 19890 0 19946 480 6 right_bottom_grid_pin_7_
port 50 nsew default input
rlabel metal3 s 23520 18912 24000 19032 6 right_bottom_grid_pin_9_
port 51 nsew default input
rlabel metal3 s 0 18504 480 18624 6 right_top_grid_pin_10_
port 52 nsew default input
rlabel metal3 s 0 22040 480 22160 6 top_left_grid_pin_11_
port 53 nsew default input
rlabel metal3 s 0 23264 480 23384 6 top_left_grid_pin_13_
port 54 nsew default input
rlabel metal2 s 22742 23520 22798 24000 6 top_left_grid_pin_15_
port 55 nsew default input
rlabel metal3 s 0 19592 480 19712 6 top_left_grid_pin_1_
port 56 nsew default input
rlabel metal2 s 23110 0 23166 480 6 top_left_grid_pin_3_
port 57 nsew default input
rlabel metal3 s 0 20816 480 20936 6 top_left_grid_pin_5_
port 58 nsew default input
rlabel metal2 s 20350 23520 20406 24000 6 top_left_grid_pin_7_
port 59 nsew default input
rlabel metal3 s 23520 21768 24000 21888 6 top_left_grid_pin_9_
port 60 nsew default input
rlabel metal3 s 23520 23128 24000 23248 6 top_right_grid_pin_11_
port 61 nsew default input
rlabel metal4 s 4944 2128 5264 21808 6 vpwr
port 62 nsew default input
rlabel metal4 s 8944 2128 9264 21808 6 vgnd
port 63 nsew default input
<< end >>
