magic
tech EFS8A
magscale 1 2
timestamp 1602873179
<< locali >>
rect 24685 11679 24719 11781
rect 2651 11577 2789 11611
rect 20821 10523 20855 10761
rect 33885 9911 33919 10217
rect 5871 9673 6009 9707
rect 11431 9129 11437 9163
rect 34063 9129 34069 9163
rect 35811 9129 35817 9163
rect 11431 9061 11465 9129
rect 34063 9061 34097 9129
rect 35811 9061 35845 9129
rect 17819 8993 17946 9027
rect 2139 8041 2145 8075
rect 2139 7973 2173 8041
rect 10977 7191 11011 7293
rect 32505 7191 32539 7293
rect 19268 6885 19336 6919
rect 32413 6171 32447 6341
rect 23575 5865 23581 5899
rect 14933 5695 14967 5865
rect 23575 5797 23609 5865
rect 32079 5729 32206 5763
rect 35035 5321 35173 5355
rect 10333 5083 10367 5321
rect 16589 4471 16623 4777
rect 29687 4641 29722 4675
rect 6377 3927 6411 4165
rect 18981 4063 19015 4165
rect 16957 3587 16991 3689
rect 5123 3553 5158 3587
rect 20545 2907 20579 3009
rect 22845 2907 22879 3077
rect 22707 2873 22845 2907
rect 22937 2839 22971 3145
rect 21465 2431 21499 2533
rect 23857 2295 23891 2397
<< viali >>
rect 1593 13481 1627 13515
rect 1409 13345 1443 13379
rect 1593 12937 1627 12971
rect 1409 12733 1443 12767
rect 24292 12733 24326 12767
rect 24685 12665 24719 12699
rect 2053 12597 2087 12631
rect 2421 12597 2455 12631
rect 24363 12597 24397 12631
rect 35633 12393 35667 12427
rect 1720 12257 1754 12291
rect 2764 12257 2798 12291
rect 11044 12257 11078 12291
rect 19165 12257 19199 12291
rect 24108 12257 24142 12291
rect 25120 12257 25154 12291
rect 34412 12257 34446 12291
rect 35449 12257 35483 12291
rect 29561 12189 29595 12223
rect 1823 12053 1857 12087
rect 2835 12053 2869 12087
rect 10149 12053 10183 12087
rect 11115 12053 11149 12087
rect 19349 12053 19383 12087
rect 24179 12053 24213 12087
rect 25191 12053 25225 12087
rect 34483 12053 34517 12087
rect 1593 11849 1627 11883
rect 20867 11849 20901 11883
rect 31769 11849 31803 11883
rect 35357 11849 35391 11883
rect 35633 11849 35667 11883
rect 36691 11849 36725 11883
rect 18797 11781 18831 11815
rect 24685 11781 24719 11815
rect 24961 11781 24995 11815
rect 2421 11713 2455 11747
rect 24133 11713 24167 11747
rect 1409 11645 1443 11679
rect 2580 11645 2614 11679
rect 10333 11645 10367 11679
rect 10517 11645 10551 11679
rect 18613 11645 18647 11679
rect 19073 11645 19107 11679
rect 20796 11645 20830 11679
rect 24476 11645 24510 11679
rect 24685 11645 24719 11679
rect 25329 11645 25363 11679
rect 30056 11645 30090 11679
rect 30481 11645 30515 11679
rect 31284 11645 31318 11679
rect 33860 11645 33894 11679
rect 34253 11645 34287 11679
rect 35449 11645 35483 11679
rect 36001 11645 36035 11679
rect 36620 11645 36654 11679
rect 37013 11645 37047 11679
rect 2789 11577 2823 11611
rect 10793 11577 10827 11611
rect 34621 11577 34655 11611
rect 1961 11509 1995 11543
rect 3065 11509 3099 11543
rect 3433 11509 3467 11543
rect 9965 11509 9999 11543
rect 11161 11509 11195 11543
rect 15669 11509 15703 11543
rect 19441 11509 19475 11543
rect 19717 11509 19751 11543
rect 21281 11509 21315 11543
rect 24547 11509 24581 11543
rect 25421 11509 25455 11543
rect 30159 11509 30193 11543
rect 31355 11509 31389 11543
rect 33931 11509 33965 11543
rect 2697 11305 2731 11339
rect 10149 11305 10183 11339
rect 15761 11305 15795 11339
rect 26663 11305 26697 11339
rect 31493 11305 31527 11339
rect 35633 11305 35667 11339
rect 11621 11237 11655 11271
rect 21097 11237 21131 11271
rect 24409 11237 24443 11271
rect 24501 11237 24535 11271
rect 29837 11237 29871 11271
rect 29929 11237 29963 11271
rect 1409 11169 1443 11203
rect 2513 11169 2547 11203
rect 4144 11169 4178 11203
rect 8585 11169 8619 11203
rect 10057 11169 10091 11203
rect 10425 11169 10459 11203
rect 13001 11169 13035 11203
rect 15485 11169 15519 11203
rect 15945 11169 15979 11203
rect 18220 11169 18254 11203
rect 19165 11169 19199 11203
rect 19625 11169 19659 11203
rect 23340 11169 23374 11203
rect 26592 11169 26626 11203
rect 27813 11169 27847 11203
rect 28273 11169 28307 11203
rect 32137 11169 32171 11203
rect 32597 11169 32631 11203
rect 34345 11169 34379 11203
rect 35449 11169 35483 11203
rect 36553 11169 36587 11203
rect 11529 11101 11563 11135
rect 19901 11101 19935 11135
rect 21005 11101 21039 11135
rect 21649 11101 21683 11135
rect 25053 11101 25087 11135
rect 28549 11101 28583 11135
rect 32689 11101 32723 11135
rect 34989 11101 35023 11135
rect 12081 11033 12115 11067
rect 13185 11033 13219 11067
rect 30389 11033 30423 11067
rect 34529 11033 34563 11067
rect 1593 10965 1627 10999
rect 4215 10965 4249 10999
rect 8769 10965 8803 10999
rect 10885 10965 10919 10999
rect 12449 10965 12483 10999
rect 18291 10965 18325 10999
rect 20177 10965 20211 10999
rect 23443 10965 23477 10999
rect 27721 10965 27755 10999
rect 35265 10965 35299 10999
rect 36737 10965 36771 10999
rect 4721 10761 4755 10795
rect 8309 10761 8343 10795
rect 11529 10761 11563 10795
rect 16727 10761 16761 10795
rect 18337 10761 18371 10795
rect 20821 10761 20855 10795
rect 21465 10761 21499 10795
rect 24041 10761 24075 10795
rect 27077 10761 27111 10795
rect 29745 10761 29779 10795
rect 34345 10761 34379 10795
rect 36645 10761 36679 10795
rect 37013 10761 37047 10795
rect 10057 10693 10091 10727
rect 13461 10693 13495 10727
rect 19809 10693 19843 10727
rect 9275 10625 9309 10659
rect 11805 10625 11839 10659
rect 12265 10625 12299 10659
rect 15393 10625 15427 10659
rect 20085 10625 20119 10659
rect 20729 10625 20763 10659
rect 1409 10557 1443 10591
rect 2564 10557 2598 10591
rect 3960 10557 3994 10591
rect 8125 10557 8159 10591
rect 8585 10557 8619 10591
rect 9188 10557 9222 10591
rect 12449 10557 12483 10591
rect 13001 10557 13035 10591
rect 16624 10557 16658 10591
rect 17049 10557 17083 10591
rect 17877 10557 17911 10591
rect 18705 10557 18739 10591
rect 18981 10557 19015 10591
rect 29101 10693 29135 10727
rect 30573 10693 30607 10727
rect 36277 10693 36311 10727
rect 24593 10625 24627 10659
rect 25513 10625 25547 10659
rect 31585 10625 31619 10659
rect 35909 10625 35943 10659
rect 21557 10557 21591 10591
rect 22017 10557 22051 10591
rect 22620 10557 22654 10591
rect 23029 10557 23063 10591
rect 26157 10557 26191 10591
rect 26525 10557 26559 10591
rect 27537 10557 27571 10591
rect 27905 10557 27939 10591
rect 28089 10557 28123 10591
rect 32965 10557 32999 10591
rect 33057 10557 33091 10591
rect 33517 10557 33551 10591
rect 33793 10557 33827 10591
rect 36461 10557 36495 10591
rect 37616 10557 37650 10591
rect 2651 10489 2685 10523
rect 10241 10489 10275 10523
rect 10333 10489 10367 10523
rect 10885 10489 10919 10523
rect 15117 10489 15151 10523
rect 15209 10489 15243 10523
rect 16129 10489 16163 10523
rect 19165 10489 19199 10523
rect 20177 10489 20211 10523
rect 20821 10489 20855 10523
rect 22707 10489 22741 10523
rect 24685 10489 24719 10523
rect 25237 10489 25271 10523
rect 25973 10489 26007 10523
rect 28365 10489 28399 10523
rect 30021 10489 30055 10523
rect 30113 10489 30147 10523
rect 31309 10489 31343 10523
rect 31677 10489 31711 10523
rect 32229 10489 32263 10523
rect 34989 10489 35023 10523
rect 35081 10489 35115 10523
rect 35633 10489 35667 10523
rect 37703 10489 37737 10523
rect 1593 10421 1627 10455
rect 2053 10421 2087 10455
rect 3065 10421 3099 10455
rect 3341 10421 3375 10455
rect 4031 10421 4065 10455
rect 4353 10421 4387 10455
rect 6837 10421 6871 10455
rect 8953 10421 8987 10455
rect 9689 10421 9723 10455
rect 12541 10421 12575 10455
rect 14013 10421 14047 10455
rect 14933 10421 14967 10455
rect 19533 10421 19567 10455
rect 21005 10421 21039 10455
rect 21741 10421 21775 10455
rect 23397 10421 23431 10455
rect 24409 10421 24443 10455
rect 26157 10421 26191 10455
rect 28641 10421 28675 10455
rect 31033 10421 31067 10455
rect 32505 10421 32539 10455
rect 38025 10421 38059 10455
rect 2053 10217 2087 10251
rect 4951 10217 4985 10251
rect 10333 10217 10367 10251
rect 13737 10217 13771 10251
rect 19073 10217 19107 10251
rect 19257 10217 19291 10251
rect 20177 10217 20211 10251
rect 29469 10217 29503 10251
rect 29745 10217 29779 10251
rect 31585 10217 31619 10251
rect 32689 10217 32723 10251
rect 33885 10217 33919 10251
rect 36277 10217 36311 10251
rect 10609 10149 10643 10183
rect 12081 10149 12115 10183
rect 12173 10149 12207 10183
rect 15577 10149 15611 10183
rect 16037 10149 16071 10183
rect 21097 10149 21131 10183
rect 23305 10149 23339 10183
rect 24501 10149 24535 10183
rect 24777 10149 24811 10183
rect 24869 10149 24903 10183
rect 25421 10149 25455 10183
rect 26709 10149 26743 10183
rect 28870 10149 28904 10183
rect 30481 10149 30515 10183
rect 30573 10149 30607 10183
rect 33057 10149 33091 10183
rect 33149 10149 33183 10183
rect 33701 10149 33735 10183
rect 1961 10081 1995 10115
rect 2421 10081 2455 10115
rect 4880 10081 4914 10115
rect 7640 10081 7674 10115
rect 8620 10081 8654 10115
rect 13921 10081 13955 10115
rect 14197 10081 14231 10115
rect 17693 10081 17727 10115
rect 18153 10081 18187 10115
rect 19441 10081 19475 10115
rect 19717 10081 19751 10115
rect 21649 10081 21683 10115
rect 26157 10081 26191 10115
rect 6561 10013 6595 10047
rect 10517 10013 10551 10047
rect 12357 10013 12391 10047
rect 15025 10013 15059 10047
rect 15945 10013 15979 10047
rect 16221 10013 16255 10047
rect 18337 10013 18371 10047
rect 18705 10013 18739 10047
rect 21005 10013 21039 10047
rect 23213 10013 23247 10047
rect 23489 10013 23523 10047
rect 26617 10013 26651 10047
rect 26893 10013 26927 10047
rect 28549 10013 28583 10047
rect 31125 10013 31159 10047
rect 7711 9945 7745 9979
rect 11069 9945 11103 9979
rect 32321 9945 32355 9979
rect 34713 10149 34747 10183
rect 36645 10149 36679 10183
rect 36093 10081 36127 10115
rect 34621 10013 34655 10047
rect 34897 10013 34931 10047
rect 1685 9877 1719 9911
rect 8723 9877 8757 9911
rect 9045 9877 9079 9911
rect 9965 9877 9999 9911
rect 24133 9877 24167 9911
rect 27813 9877 27847 9911
rect 30113 9877 30147 9911
rect 33885 9877 33919 9911
rect 34069 9877 34103 9911
rect 2053 9673 2087 9707
rect 3985 9673 4019 9707
rect 5181 9673 5215 9707
rect 6009 9673 6043 9707
rect 9597 9673 9631 9707
rect 11437 9673 11471 9707
rect 11805 9673 11839 9707
rect 16589 9673 16623 9707
rect 17877 9673 17911 9707
rect 18797 9673 18831 9707
rect 20177 9673 20211 9707
rect 21925 9673 21959 9707
rect 22201 9673 22235 9707
rect 22753 9673 22787 9707
rect 23121 9673 23155 9707
rect 24593 9673 24627 9707
rect 24869 9673 24903 9707
rect 25237 9673 25271 9707
rect 26525 9673 26559 9707
rect 30849 9673 30883 9707
rect 31447 9673 31481 9707
rect 33241 9673 33275 9707
rect 33517 9673 33551 9707
rect 33977 9673 34011 9707
rect 6653 9605 6687 9639
rect 9229 9605 9263 9639
rect 13737 9605 13771 9639
rect 16221 9605 16255 9639
rect 27077 9605 27111 9639
rect 30205 9605 30239 9639
rect 30573 9605 30607 9639
rect 2329 9537 2363 9571
rect 3249 9537 3283 9571
rect 8677 9537 8711 9571
rect 10149 9537 10183 9571
rect 12541 9537 12575 9571
rect 12817 9537 12851 9571
rect 15025 9537 15059 9571
rect 19257 9537 19291 9571
rect 21005 9537 21039 9571
rect 23673 9537 23707 9571
rect 25513 9537 25547 9571
rect 25789 9537 25823 9571
rect 28365 9537 28399 9571
rect 29285 9537 29319 9571
rect 32321 9537 32355 9571
rect 34989 9537 35023 9571
rect 35265 9537 35299 9571
rect 36829 9537 36863 9571
rect 3709 9469 3743 9503
rect 4445 9469 4479 9503
rect 4629 9469 4663 9503
rect 5641 9469 5675 9503
rect 5768 9469 5802 9503
rect 6285 9469 6319 9503
rect 6837 9469 6871 9503
rect 7389 9469 7423 9503
rect 11069 9469 11103 9503
rect 12173 9469 12207 9503
rect 14080 9469 14114 9503
rect 14473 9469 14507 9503
rect 15945 9469 15979 9503
rect 17024 9469 17058 9503
rect 18312 9469 18346 9503
rect 27905 9469 27939 9503
rect 28089 9469 28123 9503
rect 31376 9469 31410 9503
rect 31769 9469 31803 9503
rect 2421 9401 2455 9435
rect 2973 9401 3007 9435
rect 8401 9401 8435 9435
rect 8769 9401 8803 9435
rect 10470 9401 10504 9435
rect 12633 9401 12667 9435
rect 14933 9401 14967 9435
rect 15387 9401 15421 9435
rect 19165 9401 19199 9435
rect 19619 9401 19653 9435
rect 20913 9401 20947 9435
rect 21367 9401 21401 9435
rect 23489 9401 23523 9435
rect 23994 9401 24028 9435
rect 25605 9401 25639 9435
rect 27537 9401 27571 9435
rect 29606 9401 29640 9435
rect 32642 9401 32676 9435
rect 34713 9401 34747 9435
rect 35081 9401 35115 9435
rect 36553 9401 36587 9435
rect 36645 9401 36679 9435
rect 1593 9333 1627 9367
rect 4261 9333 4295 9367
rect 6929 9333 6963 9367
rect 7849 9333 7883 9367
rect 9965 9333 9999 9367
rect 14151 9333 14185 9367
rect 17095 9333 17129 9367
rect 17509 9333 17543 9367
rect 18383 9333 18417 9367
rect 20545 9333 20579 9367
rect 28733 9333 28767 9367
rect 29009 9333 29043 9367
rect 32137 9333 32171 9367
rect 34345 9333 34379 9367
rect 36093 9333 36127 9367
rect 7573 9129 7607 9163
rect 8125 9129 8159 9163
rect 10149 9129 10183 9163
rect 10885 9129 10919 9163
rect 11437 9129 11471 9163
rect 11989 9129 12023 9163
rect 12449 9129 12483 9163
rect 15025 9129 15059 9163
rect 16681 9129 16715 9163
rect 17693 9129 17727 9163
rect 18705 9129 18739 9163
rect 20729 9129 20763 9163
rect 21833 9129 21867 9163
rect 25053 9129 25087 9163
rect 26617 9129 26651 9163
rect 28549 9129 28583 9163
rect 29561 9129 29595 9163
rect 34069 9129 34103 9163
rect 35265 9129 35299 9163
rect 35817 9129 35851 9163
rect 36369 9129 36403 9163
rect 36645 9129 36679 9163
rect 2605 9061 2639 9095
rect 5089 9061 5123 9095
rect 6561 9061 6595 9095
rect 6653 9061 6687 9095
rect 9827 9061 9861 9095
rect 13829 9061 13863 9095
rect 14381 9061 14415 9095
rect 16082 9061 16116 9095
rect 18981 9061 19015 9095
rect 19073 9061 19107 9095
rect 19993 9061 20027 9095
rect 23029 9061 23063 9095
rect 24178 9061 24212 9095
rect 25513 9061 25547 9095
rect 26341 9061 26375 9095
rect 28962 9061 28996 9095
rect 31217 9061 31251 9095
rect 33149 9061 33183 9095
rect 1476 8993 1510 9027
rect 8125 8993 8159 9027
rect 8493 8993 8527 9027
rect 9740 8993 9774 9027
rect 15761 8993 15795 9027
rect 17785 8993 17819 9027
rect 20948 8993 20982 9027
rect 22477 8993 22511 9027
rect 22845 8993 22879 9027
rect 24777 8993 24811 9027
rect 26525 8993 26559 9027
rect 27077 8993 27111 9027
rect 28641 8993 28675 9027
rect 30573 8993 30607 9027
rect 30941 8993 30975 9027
rect 32137 8993 32171 9027
rect 32597 8993 32631 9027
rect 34621 8993 34655 9027
rect 2513 8925 2547 8959
rect 3157 8925 3191 8959
rect 4721 8925 4755 8959
rect 4997 8925 5031 8959
rect 5273 8925 5307 8959
rect 6837 8925 6871 8959
rect 11069 8925 11103 8959
rect 13737 8925 13771 8959
rect 23857 8925 23891 8959
rect 32873 8925 32907 8959
rect 33517 8925 33551 8959
rect 33701 8925 33735 8959
rect 35449 8925 35483 8959
rect 19533 8857 19567 8891
rect 1547 8789 1581 8823
rect 1869 8789 1903 8823
rect 2329 8789 2363 8823
rect 9137 8789 9171 8823
rect 10609 8789 10643 8823
rect 12817 8789 12851 8823
rect 13461 8789 13495 8823
rect 18015 8789 18049 8823
rect 18429 8789 18463 8823
rect 21051 8789 21085 8823
rect 21557 8789 21591 8823
rect 23673 8789 23707 8823
rect 27721 8789 27755 8823
rect 30113 8789 30147 8823
rect 34989 8789 35023 8823
rect 1685 8585 1719 8619
rect 3249 8585 3283 8619
rect 3985 8585 4019 8619
rect 6285 8585 6319 8619
rect 8125 8585 8159 8619
rect 8493 8585 8527 8619
rect 9183 8585 9217 8619
rect 9965 8585 9999 8619
rect 10977 8585 11011 8619
rect 11713 8585 11747 8619
rect 13737 8585 13771 8619
rect 14013 8585 14047 8619
rect 17325 8585 17359 8619
rect 19257 8585 19291 8619
rect 20637 8585 20671 8619
rect 20913 8585 20947 8619
rect 21281 8585 21315 8619
rect 24593 8585 24627 8619
rect 24961 8585 24995 8619
rect 25513 8585 25547 8619
rect 27077 8585 27111 8619
rect 29009 8585 29043 8619
rect 31723 8585 31757 8619
rect 34069 8585 34103 8619
rect 35909 8585 35943 8619
rect 36277 8585 36311 8619
rect 36645 8585 36679 8619
rect 3617 8517 3651 8551
rect 15485 8517 15519 8551
rect 31033 8517 31067 8551
rect 2329 8449 2363 8483
rect 2973 8449 3007 8483
rect 5273 8449 5307 8483
rect 5549 8449 5583 8483
rect 6929 8449 6963 8483
rect 10057 8449 10091 8483
rect 16129 8449 16163 8483
rect 18245 8449 18279 8483
rect 18613 8449 18647 8483
rect 19717 8449 19751 8483
rect 25789 8449 25823 8483
rect 26433 8449 26467 8483
rect 30757 8449 30791 8483
rect 31493 8449 31527 8483
rect 35265 8449 35299 8483
rect 3801 8381 3835 8415
rect 4445 8381 4479 8415
rect 9080 8381 9114 8415
rect 9505 8381 9539 8415
rect 12817 8381 12851 8415
rect 14565 8381 14599 8415
rect 16313 8381 16347 8415
rect 16865 8381 16899 8415
rect 17877 8381 17911 8415
rect 21465 8381 21499 8415
rect 21925 8381 21959 8415
rect 23673 8381 23707 8415
rect 27629 8381 27663 8415
rect 28089 8381 28123 8415
rect 31652 8381 31686 8415
rect 32781 8381 32815 8415
rect 33701 8381 33735 8415
rect 34621 8381 34655 8415
rect 36461 8381 36495 8415
rect 37013 8381 37047 8415
rect 2145 8313 2179 8347
rect 2421 8313 2455 8347
rect 5089 8313 5123 8347
rect 5365 8313 5399 8347
rect 6653 8313 6687 8347
rect 7250 8313 7284 8347
rect 10378 8313 10412 8347
rect 11345 8313 11379 8347
rect 12633 8313 12667 8347
rect 13138 8313 13172 8347
rect 14927 8313 14961 8347
rect 17049 8313 17083 8347
rect 18337 8313 18371 8347
rect 19625 8313 19659 8347
rect 20079 8313 20113 8347
rect 24035 8313 24069 8347
rect 25881 8313 25915 8347
rect 28365 8313 28399 8347
rect 29929 8313 29963 8347
rect 30113 8313 30147 8347
rect 30205 8313 30239 8347
rect 32597 8313 32631 8347
rect 33143 8313 33177 8347
rect 34989 8313 35023 8347
rect 35081 8313 35115 8347
rect 7849 8245 7883 8279
rect 14473 8245 14507 8279
rect 15761 8245 15795 8279
rect 21557 8245 21591 8279
rect 22477 8245 22511 8279
rect 22937 8245 22971 8279
rect 23489 8245 23523 8279
rect 26709 8245 26743 8279
rect 27445 8245 27479 8279
rect 28733 8245 28767 8279
rect 32137 8245 32171 8279
rect 2145 8041 2179 8075
rect 2697 8041 2731 8075
rect 3893 8041 3927 8075
rect 5825 8041 5859 8075
rect 6561 8041 6595 8075
rect 7757 8041 7791 8075
rect 8723 8041 8757 8075
rect 13185 8041 13219 8075
rect 16957 8041 16991 8075
rect 18521 8041 18555 8075
rect 18981 8041 19015 8075
rect 20085 8041 20119 8075
rect 25421 8041 25455 8075
rect 25789 8041 25823 8075
rect 30665 8041 30699 8075
rect 32413 8041 32447 8075
rect 34437 8041 34471 8075
rect 3525 7973 3559 8007
rect 4169 7973 4203 8007
rect 4261 7973 4295 8007
rect 4813 7973 4847 8007
rect 5181 7973 5215 8007
rect 7199 7973 7233 8007
rect 11253 7973 11287 8007
rect 14381 7973 14415 8007
rect 14657 7973 14691 8007
rect 15663 7973 15697 8007
rect 17601 7973 17635 8007
rect 17693 7973 17727 8007
rect 19165 7973 19199 8007
rect 19257 7973 19291 8007
rect 21649 7973 21683 8007
rect 24822 7973 24856 8007
rect 26887 7973 26921 8007
rect 29238 7973 29272 8007
rect 33879 7973 33913 8007
rect 35449 7973 35483 8007
rect 1777 7905 1811 7939
rect 5641 7905 5675 7939
rect 8652 7905 8686 7939
rect 10793 7905 10827 7939
rect 11069 7905 11103 7939
rect 12081 7905 12115 7939
rect 12633 7905 12667 7939
rect 13645 7905 13679 7939
rect 14197 7905 14231 7939
rect 23029 7905 23063 7939
rect 23213 7905 23247 7939
rect 23949 7905 23983 7939
rect 29837 7905 29871 7939
rect 32572 7905 32606 7939
rect 6837 7837 6871 7871
rect 12817 7837 12851 7871
rect 15301 7837 15335 7871
rect 18245 7837 18279 7871
rect 19533 7837 19567 7871
rect 21281 7837 21315 7871
rect 21557 7837 21591 7871
rect 21833 7837 21867 7871
rect 23581 7837 23615 7871
rect 24501 7837 24535 7871
rect 26525 7837 26559 7871
rect 28917 7837 28951 7871
rect 30113 7837 30147 7871
rect 33517 7837 33551 7871
rect 35357 7837 35391 7871
rect 35633 7837 35667 7871
rect 16221 7769 16255 7803
rect 30481 7769 30515 7803
rect 3065 7701 3099 7735
rect 5457 7701 5491 7735
rect 10057 7701 10091 7735
rect 13553 7701 13587 7735
rect 16589 7701 16623 7735
rect 24225 7701 24259 7735
rect 27445 7701 27479 7735
rect 27721 7701 27755 7735
rect 32643 7701 32677 7735
rect 33241 7701 33275 7735
rect 34897 7701 34931 7735
rect 3157 7497 3191 7531
rect 8769 7497 8803 7531
rect 9597 7497 9631 7531
rect 11805 7497 11839 7531
rect 14565 7497 14599 7531
rect 15301 7497 15335 7531
rect 17601 7497 17635 7531
rect 19625 7497 19659 7531
rect 20085 7497 20119 7531
rect 22385 7497 22419 7531
rect 23489 7497 23523 7531
rect 32689 7497 32723 7531
rect 34253 7497 34287 7531
rect 35909 7497 35943 7531
rect 36645 7497 36679 7531
rect 11253 7429 11287 7463
rect 28273 7429 28307 7463
rect 32367 7429 32401 7463
rect 4169 7361 4203 7395
rect 5733 7361 5767 7395
rect 10241 7361 10275 7395
rect 13645 7361 13679 7395
rect 13921 7361 13955 7395
rect 16221 7361 16255 7395
rect 18705 7361 18739 7395
rect 19349 7361 19383 7395
rect 21465 7361 21499 7395
rect 24225 7361 24259 7395
rect 25881 7361 25915 7395
rect 27721 7361 27755 7395
rect 28917 7361 28951 7395
rect 29929 7361 29963 7395
rect 30113 7361 30147 7395
rect 34621 7361 34655 7395
rect 34989 7361 35023 7395
rect 35357 7361 35391 7395
rect 2237 7293 2271 7327
rect 6653 7293 6687 7327
rect 6837 7293 6871 7327
rect 7849 7293 7883 7327
rect 10057 7293 10091 7327
rect 10885 7293 10919 7327
rect 10977 7293 11011 7327
rect 12576 7293 12610 7327
rect 13001 7293 13035 7327
rect 15117 7293 15151 7327
rect 15669 7293 15703 7327
rect 16129 7293 16163 7327
rect 17141 7293 17175 7327
rect 18429 7293 18463 7327
rect 20228 7293 20262 7327
rect 20637 7293 20671 7327
rect 23949 7293 23983 7327
rect 24133 7293 24167 7327
rect 26801 7293 26835 7327
rect 27445 7293 27479 7327
rect 32264 7293 32298 7327
rect 32505 7293 32539 7327
rect 36461 7293 36495 7327
rect 1869 7225 1903 7259
rect 2599 7225 2633 7259
rect 4077 7225 4111 7259
rect 4531 7225 4565 7259
rect 7389 7225 7423 7259
rect 7757 7225 7791 7259
rect 8170 7225 8204 7259
rect 9321 7225 9355 7259
rect 10333 7225 10367 7259
rect 13369 7225 13403 7259
rect 13737 7225 13771 7259
rect 15025 7225 15059 7259
rect 16583 7225 16617 7259
rect 18797 7225 18831 7259
rect 20315 7225 20349 7259
rect 21373 7225 21407 7259
rect 21827 7225 21861 7259
rect 25697 7225 25731 7259
rect 26202 7225 26236 7259
rect 27077 7225 27111 7259
rect 27813 7225 27847 7259
rect 30434 7225 30468 7259
rect 33333 7225 33367 7259
rect 33425 7225 33459 7259
rect 33977 7225 34011 7259
rect 35081 7225 35115 7259
rect 37013 7225 37047 7259
rect 3525 7157 3559 7191
rect 5089 7157 5123 7191
rect 6285 7157 6319 7191
rect 7021 7157 7055 7191
rect 10977 7157 11011 7191
rect 12173 7157 12207 7191
rect 12679 7157 12713 7191
rect 22661 7157 22695 7191
rect 23029 7157 23063 7191
rect 24685 7157 24719 7191
rect 25053 7157 25087 7191
rect 29469 7157 29503 7191
rect 31033 7157 31067 7191
rect 32505 7157 32539 7191
rect 33149 7157 33183 7191
rect 1777 6953 1811 6987
rect 3433 6953 3467 6987
rect 8769 6953 8803 6987
rect 14013 6953 14047 6987
rect 14381 6953 14415 6987
rect 17509 6953 17543 6987
rect 18521 6953 18555 6987
rect 19901 6953 19935 6987
rect 21925 6953 21959 6987
rect 25973 6953 26007 6987
rect 30297 6953 30331 6987
rect 33885 6953 33919 6987
rect 35449 6953 35483 6987
rect 2558 6885 2592 6919
rect 3893 6885 3927 6919
rect 4537 6885 4571 6919
rect 6923 6885 6957 6919
rect 10010 6885 10044 6919
rect 12310 6885 12344 6919
rect 13737 6885 13771 6919
rect 15853 6885 15887 6919
rect 16129 6885 16163 6919
rect 19234 6885 19268 6919
rect 21005 6885 21039 6919
rect 21097 6885 21131 6919
rect 22293 6885 22327 6919
rect 24501 6885 24535 6919
rect 27261 6885 27295 6919
rect 28825 6885 28859 6919
rect 32458 6885 32492 6919
rect 34621 6885 34655 6919
rect 35173 6885 35207 6919
rect 36185 6885 36219 6919
rect 6561 6817 6595 6851
rect 8585 6817 8619 6851
rect 10609 6817 10643 6851
rect 14197 6817 14231 6851
rect 17601 6817 17635 6851
rect 17785 6817 17819 6851
rect 20637 6817 20671 6851
rect 21649 6817 21683 6851
rect 22512 6817 22546 6851
rect 24041 6817 24075 6851
rect 24317 6817 24351 6851
rect 25329 6817 25363 6851
rect 30481 6817 30515 6851
rect 30941 6817 30975 6851
rect 2237 6749 2271 6783
rect 4445 6749 4479 6783
rect 4721 6749 4755 6783
rect 9689 6749 9723 6783
rect 11989 6749 12023 6783
rect 16037 6749 16071 6783
rect 16313 6749 16347 6783
rect 18153 6749 18187 6783
rect 18981 6749 19015 6783
rect 27169 6749 27203 6783
rect 27537 6749 27571 6783
rect 28549 6749 28583 6783
rect 28733 6749 28767 6783
rect 29377 6749 29411 6783
rect 31217 6749 31251 6783
rect 32137 6749 32171 6783
rect 34529 6749 34563 6783
rect 36093 6749 36127 6783
rect 36369 6749 36403 6783
rect 25513 6681 25547 6715
rect 3157 6613 3191 6647
rect 7481 6613 7515 6647
rect 7941 6613 7975 6647
rect 9045 6613 9079 6647
rect 12909 6613 12943 6647
rect 16957 6613 16991 6647
rect 18889 6613 18923 6647
rect 22615 6613 22649 6647
rect 26709 6613 26743 6647
rect 33057 6613 33091 6647
rect 33517 6613 33551 6647
rect 1593 6409 1627 6443
rect 2329 6409 2363 6443
rect 4169 6409 4203 6443
rect 5273 6409 5307 6443
rect 6653 6409 6687 6443
rect 8309 6409 8343 6443
rect 10057 6409 10091 6443
rect 13369 6409 13403 6443
rect 15301 6409 15335 6443
rect 16313 6409 16347 6443
rect 17693 6409 17727 6443
rect 21281 6409 21315 6443
rect 23121 6409 23155 6443
rect 24961 6409 24995 6443
rect 25329 6409 25363 6443
rect 27169 6409 27203 6443
rect 28733 6409 28767 6443
rect 31033 6409 31067 6443
rect 33885 6409 33919 6443
rect 36599 6409 36633 6443
rect 11989 6341 12023 6375
rect 14381 6341 14415 6375
rect 16957 6341 16991 6375
rect 18245 6341 18279 6375
rect 21833 6341 21867 6375
rect 30481 6341 30515 6375
rect 32229 6341 32263 6375
rect 32413 6341 32447 6375
rect 32505 6341 32539 6375
rect 34253 6341 34287 6375
rect 36001 6341 36035 6375
rect 2053 6273 2087 6307
rect 2789 6273 2823 6307
rect 3065 6273 3099 6307
rect 6285 6273 6319 6307
rect 7573 6273 7607 6307
rect 11069 6273 11103 6307
rect 14749 6273 14783 6307
rect 18521 6273 18555 6307
rect 18797 6273 18831 6307
rect 27721 6273 27755 6307
rect 27997 6273 28031 6307
rect 29653 6273 29687 6307
rect 1409 6205 1443 6239
rect 8677 6205 8711 6239
rect 8861 6205 8895 6239
rect 12449 6205 12483 6239
rect 13645 6205 13679 6239
rect 14105 6205 14139 6239
rect 14197 6205 14231 6239
rect 15393 6205 15427 6239
rect 19993 6205 20027 6239
rect 22017 6205 22051 6239
rect 22477 6205 22511 6239
rect 23673 6205 23707 6239
rect 25881 6205 25915 6239
rect 31125 6205 31159 6239
rect 31585 6205 31619 6239
rect 31861 6205 31895 6239
rect 35357 6273 35391 6307
rect 32689 6205 32723 6239
rect 33609 6205 33643 6239
rect 34621 6205 34655 6239
rect 36528 6205 36562 6239
rect 2881 6137 2915 6171
rect 4353 6137 4387 6171
rect 4445 6137 4479 6171
rect 4997 6137 5031 6171
rect 6929 6137 6963 6171
rect 7021 6137 7055 6171
rect 10793 6137 10827 6171
rect 10885 6137 10919 6171
rect 12770 6137 12804 6171
rect 15714 6137 15748 6171
rect 18613 6137 18647 6171
rect 19533 6137 19567 6171
rect 19901 6137 19935 6171
rect 20355 6137 20389 6171
rect 24035 6137 24069 6171
rect 25697 6137 25731 6171
rect 26202 6137 26236 6171
rect 27813 6137 27847 6171
rect 29377 6137 29411 6171
rect 29469 6137 29503 6171
rect 32413 6137 32447 6171
rect 33010 6137 33044 6171
rect 34989 6137 35023 6171
rect 35081 6137 35115 6171
rect 3709 6069 3743 6103
rect 7849 6069 7883 6103
rect 8493 6069 8527 6103
rect 9781 6069 9815 6103
rect 10609 6069 10643 6103
rect 16589 6069 16623 6103
rect 20913 6069 20947 6103
rect 22293 6069 22327 6103
rect 23489 6069 23523 6103
rect 24593 6069 24627 6103
rect 26801 6069 26835 6103
rect 27537 6069 27571 6103
rect 29009 6069 29043 6103
rect 36921 6069 36955 6103
rect 1685 5865 1719 5899
rect 2973 5865 3007 5899
rect 3249 5865 3283 5899
rect 5089 5865 5123 5899
rect 6745 5865 6779 5899
rect 7297 5865 7331 5899
rect 8493 5865 8527 5899
rect 10609 5865 10643 5899
rect 13093 5865 13127 5899
rect 13553 5865 13587 5899
rect 14933 5865 14967 5899
rect 18521 5865 18555 5899
rect 22477 5865 22511 5899
rect 23581 5865 23615 5899
rect 24409 5865 24443 5899
rect 26341 5865 26375 5899
rect 31125 5865 31159 5899
rect 32689 5865 32723 5899
rect 33563 5865 33597 5899
rect 34253 5865 34287 5899
rect 35449 5865 35483 5899
rect 36461 5865 36495 5899
rect 2053 5797 2087 5831
rect 4261 5797 4295 5831
rect 5825 5797 5859 5831
rect 10010 5797 10044 5831
rect 12265 5797 12299 5831
rect 13737 5797 13771 5831
rect 13829 5797 13863 5831
rect 3617 5729 3651 5763
rect 4813 5729 4847 5763
rect 7113 5729 7147 5763
rect 7481 5729 7515 5763
rect 7757 5729 7791 5763
rect 15485 5797 15519 5831
rect 16957 5797 16991 5831
rect 17049 5797 17083 5831
rect 18975 5797 19009 5831
rect 21097 5797 21131 5831
rect 21649 5797 21683 5831
rect 27169 5797 27203 5831
rect 27721 5797 27755 5831
rect 28733 5797 28767 5831
rect 30849 5797 30883 5831
rect 34621 5797 34655 5831
rect 35173 5797 35207 5831
rect 18613 5729 18647 5763
rect 24961 5729 24995 5763
rect 25145 5729 25179 5763
rect 30113 5729 30147 5763
rect 30665 5729 30699 5763
rect 32045 5729 32079 5763
rect 33492 5729 33526 5763
rect 36052 5729 36086 5763
rect 1961 5661 1995 5695
rect 4169 5661 4203 5695
rect 5733 5661 5767 5695
rect 6009 5661 6043 5695
rect 9689 5661 9723 5695
rect 12173 5661 12207 5695
rect 14381 5661 14415 5695
rect 14933 5661 14967 5695
rect 15393 5661 15427 5695
rect 15669 5661 15703 5695
rect 17233 5661 17267 5695
rect 21005 5661 21039 5695
rect 23213 5661 23247 5695
rect 25513 5661 25547 5695
rect 26893 5661 26927 5695
rect 27077 5661 27111 5695
rect 28641 5661 28675 5695
rect 29653 5661 29687 5695
rect 32275 5661 32309 5695
rect 34529 5661 34563 5695
rect 36139 5661 36173 5695
rect 2513 5593 2547 5627
rect 10885 5593 10919 5627
rect 12725 5593 12759 5627
rect 17969 5593 18003 5627
rect 19533 5593 19567 5627
rect 19901 5593 19935 5627
rect 29193 5593 29227 5627
rect 8861 5525 8895 5559
rect 11989 5525 12023 5559
rect 14749 5525 14783 5559
rect 15117 5525 15151 5559
rect 16497 5525 16531 5559
rect 20177 5525 20211 5559
rect 20729 5525 20763 5559
rect 22109 5525 22143 5559
rect 24133 5525 24167 5559
rect 25881 5525 25915 5559
rect 28089 5525 28123 5559
rect 2513 5321 2547 5355
rect 3617 5321 3651 5355
rect 4629 5321 4663 5355
rect 4997 5321 5031 5355
rect 5641 5321 5675 5355
rect 5917 5321 5951 5355
rect 10333 5321 10367 5355
rect 10425 5321 10459 5355
rect 12081 5321 12115 5355
rect 14197 5321 14231 5355
rect 14565 5321 14599 5355
rect 17325 5321 17359 5355
rect 18337 5321 18371 5355
rect 19349 5321 19383 5355
rect 20545 5321 20579 5355
rect 20913 5321 20947 5355
rect 22477 5321 22511 5355
rect 26893 5321 26927 5355
rect 28549 5321 28583 5355
rect 29423 5321 29457 5355
rect 29837 5321 29871 5355
rect 30113 5321 30147 5355
rect 30757 5321 30791 5355
rect 33517 5321 33551 5355
rect 34161 5321 34195 5355
rect 34529 5321 34563 5355
rect 35173 5321 35207 5355
rect 36093 5321 36127 5355
rect 6653 5253 6687 5287
rect 7297 5253 7331 5287
rect 9137 5253 9171 5287
rect 1593 5117 1627 5151
rect 2789 5117 2823 5151
rect 3709 5117 3743 5151
rect 5733 5117 5767 5151
rect 7113 5117 7147 5151
rect 7573 5117 7607 5151
rect 8217 5117 8251 5151
rect 25053 5253 25087 5287
rect 26249 5253 26283 5287
rect 30435 5253 30469 5287
rect 14749 5185 14783 5219
rect 15393 5185 15427 5219
rect 20177 5185 20211 5219
rect 25881 5185 25915 5219
rect 27813 5185 27847 5219
rect 29009 5185 29043 5219
rect 31447 5185 31481 5219
rect 31769 5185 31803 5219
rect 10609 5117 10643 5151
rect 13829 5117 13863 5151
rect 16221 5117 16255 5151
rect 16773 5117 16807 5151
rect 18245 5117 18279 5151
rect 18981 5117 19015 5151
rect 19625 5117 19659 5151
rect 19993 5117 20027 5151
rect 21373 5117 21407 5151
rect 23765 5117 23799 5151
rect 24225 5117 24259 5151
rect 25237 5117 25271 5151
rect 25789 5117 25823 5151
rect 29352 5117 29386 5151
rect 30364 5117 30398 5151
rect 31360 5117 31394 5151
rect 34964 5117 34998 5151
rect 1955 5049 1989 5083
rect 4071 5049 4105 5083
rect 8125 5049 8159 5083
rect 8579 5049 8613 5083
rect 9689 5049 9723 5083
rect 10333 5049 10367 5083
rect 10930 5049 10964 5083
rect 13185 5049 13219 5083
rect 13277 5049 13311 5083
rect 14841 5049 14875 5083
rect 16129 5049 16163 5083
rect 17877 5049 17911 5083
rect 18061 5049 18095 5083
rect 21281 5049 21315 5083
rect 22937 5049 22971 5083
rect 27169 5049 27203 5083
rect 27261 5049 27295 5083
rect 3249 4981 3283 5015
rect 6285 4981 6319 5015
rect 10057 4981 10091 5015
rect 11529 4981 11563 5015
rect 12909 4981 12943 5015
rect 15761 4981 15795 5015
rect 16313 4981 16347 5015
rect 23305 4981 23339 5015
rect 23765 4981 23799 5015
rect 24685 4981 24719 5015
rect 28181 4981 28215 5015
rect 32137 4981 32171 5015
rect 35449 4981 35483 5015
rect 1961 4777 1995 4811
rect 2237 4777 2271 4811
rect 3709 4777 3743 4811
rect 4169 4777 4203 4811
rect 5549 4777 5583 4811
rect 7665 4777 7699 4811
rect 9505 4777 9539 4811
rect 11989 4777 12023 4811
rect 12357 4777 12391 4811
rect 13185 4777 13219 4811
rect 13461 4777 13495 4811
rect 14749 4777 14783 4811
rect 16589 4777 16623 4811
rect 19257 4777 19291 4811
rect 20637 4777 20671 4811
rect 20913 4777 20947 4811
rect 23765 4777 23799 4811
rect 27537 4777 27571 4811
rect 29791 4777 29825 4811
rect 30205 4777 30239 4811
rect 2605 4709 2639 4743
rect 6377 4709 6411 4743
rect 13829 4709 13863 4743
rect 14381 4709 14415 4743
rect 15301 4709 15335 4743
rect 16497 4709 16531 4743
rect 1476 4641 1510 4675
rect 4353 4641 4387 4675
rect 4629 4641 4663 4675
rect 5641 4641 5675 4675
rect 5917 4641 5951 4675
rect 7205 4641 7239 4675
rect 7481 4641 7515 4675
rect 9689 4641 9723 4675
rect 9965 4641 9999 4675
rect 12081 4641 12115 4675
rect 12541 4641 12575 4675
rect 15117 4641 15151 4675
rect 15485 4641 15519 4675
rect 2513 4573 2547 4607
rect 3157 4573 3191 4607
rect 10149 4573 10183 4607
rect 13737 4573 13771 4607
rect 15853 4573 15887 4607
rect 1547 4505 1581 4539
rect 5733 4505 5767 4539
rect 7021 4505 7055 4539
rect 7297 4505 7331 4539
rect 9781 4505 9815 4539
rect 10793 4505 10827 4539
rect 17785 4709 17819 4743
rect 18981 4709 19015 4743
rect 25513 4709 25547 4743
rect 28825 4709 28859 4743
rect 16681 4641 16715 4675
rect 18245 4641 18279 4675
rect 18797 4641 18831 4675
rect 19809 4641 19843 4675
rect 20269 4641 20303 4675
rect 22109 4641 22143 4675
rect 22937 4641 22971 4675
rect 24961 4641 24995 4675
rect 25329 4641 25363 4675
rect 27169 4641 27203 4675
rect 28273 4641 28307 4675
rect 28641 4641 28675 4675
rect 29653 4641 29687 4675
rect 16828 4573 16862 4607
rect 17049 4573 17083 4607
rect 18061 4573 18095 4607
rect 21741 4573 21775 4607
rect 22845 4573 22879 4607
rect 25789 4573 25823 4607
rect 26525 4573 26559 4607
rect 19993 4505 20027 4539
rect 23213 4505 23247 4539
rect 8401 4437 8435 4471
rect 8861 4437 8895 4471
rect 16589 4437 16623 4471
rect 16957 4437 16991 4471
rect 17141 4437 17175 4471
rect 19717 4437 19751 4471
rect 24501 4437 24535 4471
rect 1685 4233 1719 4267
rect 2881 4233 2915 4267
rect 4537 4233 4571 4267
rect 5273 4233 5307 4267
rect 7113 4233 7147 4267
rect 12265 4233 12299 4267
rect 13737 4233 13771 4267
rect 16313 4233 16347 4267
rect 19901 4233 19935 4267
rect 24041 4233 24075 4267
rect 25421 4233 25455 4267
rect 26157 4233 26191 4267
rect 27261 4233 27295 4267
rect 30205 4233 30239 4267
rect 5641 4165 5675 4199
rect 6377 4165 6411 4199
rect 9689 4165 9723 4199
rect 11897 4165 11931 4199
rect 16681 4165 16715 4199
rect 16865 4165 16899 4199
rect 17509 4165 17543 4199
rect 18981 4165 19015 4199
rect 19073 4165 19107 4199
rect 19441 4165 19475 4199
rect 19763 4165 19797 4199
rect 27721 4165 27755 4199
rect 27997 4165 28031 4199
rect 28273 4165 28307 4199
rect 2605 4097 2639 4131
rect 3341 4097 3375 4131
rect 3709 4029 3743 4063
rect 3893 4029 3927 4063
rect 4905 4029 4939 4063
rect 5733 4029 5767 4063
rect 1961 3961 1995 3995
rect 2053 3961 2087 3995
rect 10517 4097 10551 4131
rect 13001 4097 13035 4131
rect 14013 4097 14047 4131
rect 15577 4097 15611 4131
rect 16773 4097 16807 4131
rect 17877 4097 17911 4131
rect 19993 4097 20027 4131
rect 21557 4097 21591 4131
rect 23397 4097 23431 4131
rect 25697 4097 25731 4131
rect 29423 4097 29457 4131
rect 29837 4097 29871 4131
rect 6653 4029 6687 4063
rect 7481 4029 7515 4063
rect 8401 4029 8435 4063
rect 8493 4029 8527 4063
rect 8677 4029 8711 4063
rect 9965 4029 9999 4063
rect 10425 4029 10459 4063
rect 12449 4029 12483 4063
rect 12909 4029 12943 4063
rect 14749 4029 14783 4063
rect 15117 4029 15151 4063
rect 16552 4029 16586 4063
rect 18061 4029 18095 4063
rect 18153 4029 18187 4063
rect 18337 4029 18371 4063
rect 18981 4029 19015 4063
rect 21925 4029 21959 4063
rect 22109 4029 22143 4063
rect 22477 4029 22511 4063
rect 24501 4029 24535 4063
rect 27813 4029 27847 4063
rect 29336 4029 29370 4063
rect 30297 4029 30331 4063
rect 30757 4029 30791 4063
rect 11345 3961 11379 3995
rect 16405 3961 16439 3995
rect 19625 3961 19659 3995
rect 20637 3961 20671 3995
rect 23029 3961 23063 3995
rect 24409 3961 24443 3995
rect 24863 3961 24897 3995
rect 26341 3961 26375 3995
rect 26433 3961 26467 3995
rect 26985 3961 27019 3995
rect 28641 3961 28675 3995
rect 3525 3893 3559 3927
rect 5917 3893 5951 3927
rect 6193 3893 6227 3927
rect 6377 3893 6411 3927
rect 7849 3893 7883 3927
rect 8217 3893 8251 3927
rect 8861 3893 8895 3927
rect 11069 3893 11103 3927
rect 15853 3893 15887 3927
rect 18521 3893 18555 3927
rect 20269 3893 20303 3927
rect 21097 3893 21131 3927
rect 22753 3893 22787 3927
rect 30481 3893 30515 3927
rect 1777 3689 1811 3723
rect 2697 3689 2731 3723
rect 3065 3689 3099 3723
rect 4215 3689 4249 3723
rect 5825 3689 5859 3723
rect 6561 3689 6595 3723
rect 9229 3689 9263 3723
rect 9781 3689 9815 3723
rect 10701 3689 10735 3723
rect 12633 3689 12667 3723
rect 15945 3689 15979 3723
rect 16957 3689 16991 3723
rect 17601 3689 17635 3723
rect 20637 3689 20671 3723
rect 22661 3689 22695 3723
rect 23949 3689 23983 3723
rect 28641 3689 28675 3723
rect 5227 3621 5261 3655
rect 15577 3621 15611 3655
rect 17785 3621 17819 3655
rect 18521 3621 18555 3655
rect 19349 3621 19383 3655
rect 22293 3621 22327 3655
rect 24225 3621 24259 3655
rect 28083 3621 28117 3655
rect 29653 3621 29687 3655
rect 1961 3553 1995 3587
rect 2237 3553 2271 3587
rect 4144 3553 4178 3587
rect 5089 3553 5123 3587
rect 6377 3553 6411 3587
rect 7389 3553 7423 3587
rect 7665 3553 7699 3587
rect 9965 3553 9999 3587
rect 10241 3553 10275 3587
rect 11989 3553 12023 3587
rect 12909 3553 12943 3587
rect 13829 3553 13863 3587
rect 14013 3553 14047 3587
rect 14381 3553 14415 3587
rect 16405 3553 16439 3587
rect 16957 3553 16991 3587
rect 18797 3553 18831 3587
rect 19533 3553 19567 3587
rect 21189 3553 21223 3587
rect 21373 3553 21407 3587
rect 21741 3553 21775 3587
rect 22845 3553 22879 3587
rect 23673 3553 23707 3587
rect 24869 3553 24903 3587
rect 26560 3553 26594 3587
rect 27721 3553 27755 3587
rect 3525 3485 3559 3519
rect 7481 3485 7515 3519
rect 8125 3485 8159 3519
rect 8493 3485 8527 3519
rect 12265 3485 12299 3519
rect 16773 3485 16807 3519
rect 17049 3485 17083 3519
rect 17932 3485 17966 3519
rect 18153 3485 18187 3519
rect 19901 3485 19935 3519
rect 22017 3485 22051 3519
rect 23765 3485 23799 3519
rect 29561 3485 29595 3519
rect 18061 3417 18095 3451
rect 20177 3417 20211 3451
rect 30113 3417 30147 3451
rect 7205 3349 7239 3383
rect 14933 3349 14967 3383
rect 19165 3349 19199 3383
rect 24593 3349 24627 3383
rect 25237 3349 25271 3383
rect 26249 3349 26283 3383
rect 26663 3349 26697 3383
rect 26985 3349 27019 3383
rect 1777 3145 1811 3179
rect 3847 3145 3881 3179
rect 4629 3145 4663 3179
rect 5089 3145 5123 3179
rect 5641 3145 5675 3179
rect 5917 3145 5951 3179
rect 7389 3145 7423 3179
rect 8769 3145 8803 3179
rect 10609 3145 10643 3179
rect 11483 3145 11517 3179
rect 13415 3145 13449 3179
rect 15485 3145 15519 3179
rect 17509 3145 17543 3179
rect 18245 3145 18279 3179
rect 22937 3145 22971 3179
rect 27261 3145 27295 3179
rect 27629 3145 27663 3179
rect 27997 3145 28031 3179
rect 30757 3145 30791 3179
rect 3433 3077 3467 3111
rect 6653 3077 6687 3111
rect 7757 3077 7791 3111
rect 10241 3077 10275 3111
rect 15117 3077 15151 3111
rect 16497 3077 16531 3111
rect 18521 3077 18555 3111
rect 22845 3077 22879 3111
rect 2697 3009 2731 3043
rect 8125 3009 8159 3043
rect 9137 3009 9171 3043
rect 13185 3009 13219 3043
rect 15209 3009 15243 3043
rect 17785 3009 17819 3043
rect 19349 3009 19383 3043
rect 20545 3009 20579 3043
rect 20821 3009 20855 3043
rect 22385 3009 22419 3043
rect 2145 2941 2179 2975
rect 2421 2941 2455 2975
rect 2973 2941 3007 2975
rect 3776 2941 3810 2975
rect 5733 2941 5767 2975
rect 6285 2941 6319 2975
rect 7665 2941 7699 2975
rect 7941 2941 7975 2975
rect 9229 2941 9263 2975
rect 9781 2941 9815 2975
rect 11412 2941 11446 2975
rect 13312 2941 13346 2975
rect 14105 2941 14139 2975
rect 14749 2941 14783 2975
rect 14988 2941 15022 2975
rect 16037 2941 16071 2975
rect 16405 2941 16439 2975
rect 16681 2941 16715 2975
rect 17141 2941 17175 2975
rect 18061 2941 18095 2975
rect 22636 2941 22670 2975
rect 12265 2873 12299 2907
rect 13829 2873 13863 2907
rect 14841 2873 14875 2907
rect 19441 2873 19475 2907
rect 19993 2873 20027 2907
rect 20269 2873 20303 2907
rect 20545 2873 20579 2907
rect 21142 2873 21176 2907
rect 22845 2873 22879 2907
rect 23489 3077 23523 3111
rect 23673 3009 23707 3043
rect 26341 3009 26375 3043
rect 28641 3009 28675 3043
rect 29469 3009 29503 3043
rect 30113 3009 30147 3043
rect 30941 3009 30975 3043
rect 25605 2941 25639 2975
rect 27813 2941 27847 2975
rect 23994 2873 24028 2907
rect 26157 2873 26191 2907
rect 26433 2873 26467 2907
rect 26985 2873 27019 2907
rect 29561 2873 29595 2907
rect 4261 2805 4295 2839
rect 7113 2805 7147 2839
rect 9321 2805 9355 2839
rect 11897 2805 11931 2839
rect 19165 2805 19199 2839
rect 20637 2805 20671 2839
rect 21741 2805 21775 2839
rect 22109 2805 22143 2839
rect 22937 2805 22971 2839
rect 23029 2805 23063 2839
rect 24593 2805 24627 2839
rect 24869 2805 24903 2839
rect 25237 2805 25271 2839
rect 28365 2805 28399 2839
rect 29101 2805 29135 2839
rect 30389 2805 30423 2839
rect 2053 2601 2087 2635
rect 2375 2601 2409 2635
rect 8125 2601 8159 2635
rect 10057 2601 10091 2635
rect 11667 2601 11701 2635
rect 12955 2601 12989 2635
rect 14933 2601 14967 2635
rect 16589 2601 16623 2635
rect 17325 2601 17359 2635
rect 18061 2601 18095 2635
rect 18705 2601 18739 2635
rect 19073 2601 19107 2635
rect 20913 2601 20947 2635
rect 21649 2601 21683 2635
rect 22017 2601 22051 2635
rect 23765 2601 23799 2635
rect 25237 2601 25271 2635
rect 27031 2601 27065 2635
rect 29101 2601 29135 2635
rect 29469 2601 29503 2635
rect 7849 2533 7883 2567
rect 9597 2533 9631 2567
rect 14565 2533 14599 2567
rect 19441 2533 19475 2567
rect 19717 2533 19751 2567
rect 20269 2533 20303 2567
rect 21465 2533 21499 2567
rect 22569 2533 22603 2567
rect 24326 2533 24360 2567
rect 26525 2533 26559 2567
rect 29745 2533 29779 2567
rect 2272 2465 2306 2499
rect 2697 2465 2731 2499
rect 6745 2465 6779 2499
rect 7757 2465 7791 2499
rect 8677 2465 8711 2499
rect 9137 2465 9171 2499
rect 10057 2465 10091 2499
rect 10241 2465 10275 2499
rect 11596 2465 11630 2499
rect 11989 2465 12023 2499
rect 12884 2465 12918 2499
rect 13737 2465 13771 2499
rect 14473 2465 14507 2499
rect 15669 2465 15703 2499
rect 16313 2465 16347 2499
rect 16957 2465 16991 2499
rect 17141 2465 17175 2499
rect 17601 2465 17635 2499
rect 18521 2465 18555 2499
rect 21256 2465 21290 2499
rect 23121 2465 23155 2499
rect 24869 2465 24903 2499
rect 26960 2465 26994 2499
rect 27940 2465 27974 2499
rect 28365 2465 28399 2499
rect 29837 2465 29871 2499
rect 31344 2465 31378 2499
rect 31769 2465 31803 2499
rect 19625 2397 19659 2431
rect 21465 2397 21499 2431
rect 22477 2397 22511 2431
rect 23857 2397 23891 2431
rect 24225 2397 24259 2431
rect 25513 2397 25547 2431
rect 25697 2397 25731 2431
rect 8861 2329 8895 2363
rect 10793 2329 10827 2363
rect 21327 2329 21361 2363
rect 26157 2329 26191 2363
rect 31447 2329 31481 2363
rect 8585 2261 8619 2295
rect 13369 2261 13403 2295
rect 15209 2261 15243 2295
rect 23857 2261 23891 2295
rect 27445 2261 27479 2295
rect 28043 2261 28077 2295
<< metal1 >>
rect 5902 15512 5908 15564
rect 5960 15552 5966 15564
rect 7466 15552 7472 15564
rect 5960 15524 7472 15552
rect 5960 15512 5966 15524
rect 7466 15512 7472 15524
rect 7524 15512 7530 15564
rect 31202 15512 31208 15564
rect 31260 15552 31266 15564
rect 32490 15552 32496 15564
rect 31260 15524 32496 15552
rect 31260 15512 31266 15524
rect 32490 15512 32496 15524
rect 32548 15512 32554 15564
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 2406 13376 2412 13388
rect 1443 13348 2412 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 2406 13336 2412 13348
rect 2464 13336 2470 13388
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 106 12928 112 12980
rect 164 12968 170 12980
rect 1581 12971 1639 12977
rect 1581 12968 1593 12971
rect 164 12940 1593 12968
rect 164 12928 170 12940
rect 1581 12937 1593 12940
rect 1627 12937 1639 12971
rect 1581 12931 1639 12937
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 24280 12767 24338 12773
rect 1443 12736 2084 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 2056 12637 2084 12736
rect 24280 12733 24292 12767
rect 24326 12764 24338 12767
rect 24326 12733 24348 12764
rect 24280 12727 24348 12733
rect 24118 12656 24124 12708
rect 24176 12696 24182 12708
rect 24320 12696 24348 12727
rect 24673 12699 24731 12705
rect 24673 12696 24685 12699
rect 24176 12668 24685 12696
rect 24176 12656 24182 12668
rect 24673 12665 24685 12668
rect 24719 12665 24731 12699
rect 24673 12659 24731 12665
rect 2041 12631 2099 12637
rect 2041 12597 2053 12631
rect 2087 12628 2099 12631
rect 2130 12628 2136 12640
rect 2087 12600 2136 12628
rect 2087 12597 2099 12600
rect 2041 12591 2099 12597
rect 2130 12588 2136 12600
rect 2188 12588 2194 12640
rect 2406 12628 2412 12640
rect 2367 12600 2412 12628
rect 2406 12588 2412 12600
rect 2464 12588 2470 12640
rect 24351 12631 24409 12637
rect 24351 12597 24363 12631
rect 24397 12628 24409 12631
rect 24578 12628 24584 12640
rect 24397 12600 24584 12628
rect 24397 12597 24409 12600
rect 24351 12591 24409 12597
rect 24578 12588 24584 12600
rect 24636 12588 24642 12640
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 35621 12427 35679 12433
rect 35621 12393 35633 12427
rect 35667 12424 35679 12427
rect 39574 12424 39580 12436
rect 35667 12396 39580 12424
rect 35667 12393 35679 12396
rect 35621 12387 35679 12393
rect 39574 12384 39580 12396
rect 39632 12384 39638 12436
rect 1394 12248 1400 12300
rect 1452 12288 1458 12300
rect 1708 12291 1766 12297
rect 1708 12288 1720 12291
rect 1452 12260 1720 12288
rect 1452 12248 1458 12260
rect 1708 12257 1720 12260
rect 1754 12257 1766 12291
rect 1708 12251 1766 12257
rect 2752 12291 2810 12297
rect 2752 12257 2764 12291
rect 2798 12288 2810 12291
rect 3050 12288 3056 12300
rect 2798 12260 3056 12288
rect 2798 12257 2810 12260
rect 2752 12251 2810 12257
rect 3050 12248 3056 12260
rect 3108 12248 3114 12300
rect 11032 12291 11090 12297
rect 11032 12257 11044 12291
rect 11078 12288 11090 12291
rect 11146 12288 11152 12300
rect 11078 12260 11152 12288
rect 11078 12257 11090 12260
rect 11032 12251 11090 12257
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 19150 12288 19156 12300
rect 19111 12260 19156 12288
rect 19150 12248 19156 12260
rect 19208 12248 19214 12300
rect 24096 12291 24154 12297
rect 24096 12257 24108 12291
rect 24142 12288 24154 12291
rect 24210 12288 24216 12300
rect 24142 12260 24216 12288
rect 24142 12257 24154 12260
rect 24096 12251 24154 12257
rect 24210 12248 24216 12260
rect 24268 12248 24274 12300
rect 25108 12291 25166 12297
rect 25108 12257 25120 12291
rect 25154 12288 25166 12291
rect 25314 12288 25320 12300
rect 25154 12260 25320 12288
rect 25154 12257 25166 12260
rect 25108 12251 25166 12257
rect 25314 12248 25320 12260
rect 25372 12248 25378 12300
rect 34400 12291 34458 12297
rect 34400 12257 34412 12291
rect 34446 12288 34458 12291
rect 34606 12288 34612 12300
rect 34446 12260 34612 12288
rect 34446 12257 34458 12260
rect 34400 12251 34458 12257
rect 34606 12248 34612 12260
rect 34664 12248 34670 12300
rect 35434 12288 35440 12300
rect 35395 12260 35440 12288
rect 35434 12248 35440 12260
rect 35492 12248 35498 12300
rect 29546 12220 29552 12232
rect 29507 12192 29552 12220
rect 29546 12180 29552 12192
rect 29604 12180 29610 12232
rect 1811 12087 1869 12093
rect 1811 12053 1823 12087
rect 1857 12084 1869 12087
rect 2314 12084 2320 12096
rect 1857 12056 2320 12084
rect 1857 12053 1869 12056
rect 1811 12047 1869 12053
rect 2314 12044 2320 12056
rect 2372 12044 2378 12096
rect 2498 12044 2504 12096
rect 2556 12084 2562 12096
rect 2823 12087 2881 12093
rect 2823 12084 2835 12087
rect 2556 12056 2835 12084
rect 2556 12044 2562 12056
rect 2823 12053 2835 12056
rect 2869 12053 2881 12087
rect 10134 12084 10140 12096
rect 10095 12056 10140 12084
rect 2823 12047 2881 12053
rect 10134 12044 10140 12056
rect 10192 12044 10198 12096
rect 11103 12087 11161 12093
rect 11103 12053 11115 12087
rect 11149 12084 11161 12087
rect 11422 12084 11428 12096
rect 11149 12056 11428 12084
rect 11149 12053 11161 12056
rect 11103 12047 11161 12053
rect 11422 12044 11428 12056
rect 11480 12044 11486 12096
rect 18138 12044 18144 12096
rect 18196 12084 18202 12096
rect 19337 12087 19395 12093
rect 19337 12084 19349 12087
rect 18196 12056 19349 12084
rect 18196 12044 18202 12056
rect 19337 12053 19349 12056
rect 19383 12053 19395 12087
rect 19337 12047 19395 12053
rect 24167 12087 24225 12093
rect 24167 12053 24179 12087
rect 24213 12084 24225 12087
rect 24394 12084 24400 12096
rect 24213 12056 24400 12084
rect 24213 12053 24225 12056
rect 24167 12047 24225 12053
rect 24394 12044 24400 12056
rect 24452 12044 24458 12096
rect 24762 12044 24768 12096
rect 24820 12084 24826 12096
rect 25179 12087 25237 12093
rect 25179 12084 25191 12087
rect 24820 12056 25191 12084
rect 24820 12044 24826 12056
rect 25179 12053 25191 12056
rect 25225 12053 25237 12087
rect 25179 12047 25237 12053
rect 34471 12087 34529 12093
rect 34471 12053 34483 12087
rect 34517 12084 34529 12087
rect 34790 12084 34796 12096
rect 34517 12056 34796 12084
rect 34517 12053 34529 12056
rect 34471 12047 34529 12053
rect 34790 12044 34796 12056
rect 34848 12044 34854 12096
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 106 11840 112 11892
rect 164 11880 170 11892
rect 1581 11883 1639 11889
rect 1581 11880 1593 11883
rect 164 11852 1593 11880
rect 164 11840 170 11852
rect 1581 11849 1593 11852
rect 1627 11849 1639 11883
rect 1581 11843 1639 11849
rect 20855 11883 20913 11889
rect 20855 11849 20867 11883
rect 20901 11880 20913 11883
rect 22094 11880 22100 11892
rect 20901 11852 22100 11880
rect 20901 11849 20913 11852
rect 20855 11843 20913 11849
rect 22094 11840 22100 11852
rect 22152 11840 22158 11892
rect 31757 11883 31815 11889
rect 31757 11849 31769 11883
rect 31803 11880 31815 11883
rect 33594 11880 33600 11892
rect 31803 11852 33600 11880
rect 31803 11849 31815 11852
rect 31757 11843 31815 11849
rect 18785 11815 18843 11821
rect 18785 11781 18797 11815
rect 18831 11812 18843 11815
rect 19610 11812 19616 11824
rect 18831 11784 19616 11812
rect 18831 11781 18843 11784
rect 18785 11775 18843 11781
rect 19610 11772 19616 11784
rect 19668 11772 19674 11824
rect 24673 11815 24731 11821
rect 24673 11781 24685 11815
rect 24719 11812 24731 11815
rect 24949 11815 25007 11821
rect 24949 11812 24961 11815
rect 24719 11784 24961 11812
rect 24719 11781 24731 11784
rect 24673 11775 24731 11781
rect 24949 11781 24961 11784
rect 24995 11812 25007 11815
rect 29822 11812 29828 11824
rect 24995 11784 29828 11812
rect 24995 11781 25007 11784
rect 24949 11775 25007 11781
rect 29822 11772 29828 11784
rect 29880 11772 29886 11824
rect 2409 11747 2467 11753
rect 2409 11744 2421 11747
rect 1412 11716 2421 11744
rect 1412 11685 1440 11716
rect 2409 11713 2421 11716
rect 2455 11744 2467 11747
rect 2455 11716 4154 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11645 1455 11679
rect 1397 11639 1455 11645
rect 2568 11679 2626 11685
rect 2568 11645 2580 11679
rect 2614 11676 2626 11679
rect 4126 11676 4154 11716
rect 8294 11704 8300 11756
rect 8352 11744 8358 11756
rect 10134 11744 10140 11756
rect 8352 11716 10140 11744
rect 8352 11704 8358 11716
rect 10134 11704 10140 11716
rect 10192 11744 10198 11756
rect 11974 11744 11980 11756
rect 10192 11716 11980 11744
rect 10192 11704 10198 11716
rect 4706 11676 4712 11688
rect 2614 11648 3464 11676
rect 4126 11648 4712 11676
rect 2614 11645 2626 11648
rect 2568 11639 2626 11645
rect 2777 11611 2835 11617
rect 2777 11577 2789 11611
rect 2823 11608 2835 11611
rect 2866 11608 2872 11620
rect 2823 11580 2872 11608
rect 2823 11577 2835 11580
rect 2777 11571 2835 11577
rect 2866 11568 2872 11580
rect 2924 11568 2930 11620
rect 1394 11500 1400 11552
rect 1452 11540 1458 11552
rect 1949 11543 2007 11549
rect 1949 11540 1961 11543
rect 1452 11512 1961 11540
rect 1452 11500 1458 11512
rect 1949 11509 1961 11512
rect 1995 11509 2007 11543
rect 3050 11540 3056 11552
rect 3011 11512 3056 11540
rect 1949 11503 2007 11509
rect 3050 11500 3056 11512
rect 3108 11500 3114 11552
rect 3436 11549 3464 11648
rect 4706 11636 4712 11648
rect 4764 11676 4770 11688
rect 6638 11676 6644 11688
rect 4764 11648 6644 11676
rect 4764 11636 4770 11648
rect 6638 11636 6644 11648
rect 6696 11636 6702 11688
rect 10336 11685 10364 11716
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 24121 11747 24179 11753
rect 24121 11713 24133 11747
rect 24167 11744 24179 11747
rect 24210 11744 24216 11756
rect 24167 11716 24216 11744
rect 24167 11713 24179 11716
rect 24121 11707 24179 11713
rect 24210 11704 24216 11716
rect 24268 11744 24274 11756
rect 28442 11744 28448 11756
rect 24268 11716 28448 11744
rect 24268 11704 24274 11716
rect 28442 11704 28448 11716
rect 28500 11704 28506 11756
rect 10321 11679 10379 11685
rect 10321 11645 10333 11679
rect 10367 11645 10379 11679
rect 10505 11679 10563 11685
rect 10505 11676 10517 11679
rect 10321 11639 10379 11645
rect 10428 11648 10517 11676
rect 10428 11552 10456 11648
rect 10505 11645 10517 11648
rect 10551 11645 10563 11679
rect 10505 11639 10563 11645
rect 15654 11636 15660 11688
rect 15712 11676 15718 11688
rect 18601 11679 18659 11685
rect 18601 11676 18613 11679
rect 15712 11648 18613 11676
rect 15712 11636 15718 11648
rect 18601 11645 18613 11648
rect 18647 11676 18659 11679
rect 19061 11679 19119 11685
rect 19061 11676 19073 11679
rect 18647 11648 19073 11676
rect 18647 11645 18659 11648
rect 18601 11639 18659 11645
rect 19061 11645 19073 11648
rect 19107 11645 19119 11679
rect 19061 11639 19119 11645
rect 20784 11679 20842 11685
rect 20784 11645 20796 11679
rect 20830 11676 20842 11679
rect 20830 11648 21312 11676
rect 20830 11645 20842 11648
rect 20784 11639 20842 11645
rect 10778 11608 10784 11620
rect 10739 11580 10784 11608
rect 10778 11568 10784 11580
rect 10836 11568 10842 11620
rect 3421 11543 3479 11549
rect 3421 11509 3433 11543
rect 3467 11540 3479 11543
rect 3602 11540 3608 11552
rect 3467 11512 3608 11540
rect 3467 11509 3479 11512
rect 3421 11503 3479 11509
rect 3602 11500 3608 11512
rect 3660 11500 3666 11552
rect 9953 11543 10011 11549
rect 9953 11509 9965 11543
rect 9999 11540 10011 11543
rect 10410 11540 10416 11552
rect 9999 11512 10416 11540
rect 9999 11509 10011 11512
rect 9953 11503 10011 11509
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 11146 11540 11152 11552
rect 11107 11512 11152 11540
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 15657 11543 15715 11549
rect 15657 11509 15669 11543
rect 15703 11540 15715 11543
rect 15930 11540 15936 11552
rect 15703 11512 15936 11540
rect 15703 11509 15715 11512
rect 15657 11503 15715 11509
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 16574 11500 16580 11552
rect 16632 11540 16638 11552
rect 19150 11540 19156 11552
rect 16632 11512 19156 11540
rect 16632 11500 16638 11512
rect 19150 11500 19156 11512
rect 19208 11540 19214 11552
rect 19429 11543 19487 11549
rect 19429 11540 19441 11543
rect 19208 11512 19441 11540
rect 19208 11500 19214 11512
rect 19429 11509 19441 11512
rect 19475 11509 19487 11543
rect 19702 11540 19708 11552
rect 19663 11512 19708 11540
rect 19429 11503 19487 11509
rect 19702 11500 19708 11512
rect 19760 11500 19766 11552
rect 21284 11549 21312 11648
rect 21358 11636 21364 11688
rect 21416 11676 21422 11688
rect 24464 11679 24522 11685
rect 24464 11676 24476 11679
rect 21416 11648 24476 11676
rect 21416 11636 21422 11648
rect 24464 11645 24476 11648
rect 24510 11676 24522 11679
rect 24673 11679 24731 11685
rect 24673 11676 24685 11679
rect 24510 11648 24685 11676
rect 24510 11645 24522 11648
rect 24464 11639 24522 11645
rect 24673 11645 24685 11648
rect 24719 11645 24731 11679
rect 25314 11676 25320 11688
rect 25275 11648 25320 11676
rect 24673 11639 24731 11645
rect 25314 11636 25320 11648
rect 25372 11636 25378 11688
rect 30044 11679 30102 11685
rect 30044 11676 30056 11679
rect 29288 11648 30056 11676
rect 22002 11568 22008 11620
rect 22060 11608 22066 11620
rect 29288 11608 29316 11648
rect 30044 11645 30056 11648
rect 30090 11676 30102 11679
rect 30469 11679 30527 11685
rect 30469 11676 30481 11679
rect 30090 11648 30481 11676
rect 30090 11645 30102 11648
rect 30044 11639 30102 11645
rect 30469 11645 30481 11648
rect 30515 11645 30527 11679
rect 30469 11639 30527 11645
rect 31272 11679 31330 11685
rect 31272 11645 31284 11679
rect 31318 11676 31330 11679
rect 31772 11676 31800 11843
rect 33594 11840 33600 11852
rect 33652 11880 33658 11892
rect 35345 11883 35403 11889
rect 35345 11880 35357 11883
rect 33652 11852 35357 11880
rect 33652 11840 33658 11852
rect 35345 11849 35357 11852
rect 35391 11880 35403 11883
rect 35434 11880 35440 11892
rect 35391 11852 35440 11880
rect 35391 11849 35403 11852
rect 35345 11843 35403 11849
rect 35434 11840 35440 11852
rect 35492 11840 35498 11892
rect 35618 11880 35624 11892
rect 35579 11852 35624 11880
rect 35618 11840 35624 11852
rect 35676 11840 35682 11892
rect 36679 11883 36737 11889
rect 36679 11849 36691 11883
rect 36725 11880 36737 11883
rect 37182 11880 37188 11892
rect 36725 11852 37188 11880
rect 36725 11849 36737 11852
rect 36679 11843 36737 11849
rect 37182 11840 37188 11852
rect 37240 11840 37246 11892
rect 34422 11704 34428 11756
rect 34480 11744 34486 11756
rect 34480 11716 36651 11744
rect 34480 11704 34486 11716
rect 31318 11648 31800 11676
rect 31318 11645 31330 11648
rect 31272 11639 31330 11645
rect 22060 11580 29316 11608
rect 30484 11608 30512 11639
rect 32582 11636 32588 11688
rect 32640 11676 32646 11688
rect 33848 11679 33906 11685
rect 33848 11676 33860 11679
rect 32640 11648 33860 11676
rect 32640 11636 32646 11648
rect 33848 11645 33860 11648
rect 33894 11676 33906 11679
rect 34241 11679 34299 11685
rect 34241 11676 34253 11679
rect 33894 11648 34253 11676
rect 33894 11645 33906 11648
rect 33848 11639 33906 11645
rect 34241 11645 34253 11648
rect 34287 11645 34299 11679
rect 34241 11639 34299 11645
rect 35158 11636 35164 11688
rect 35216 11676 35222 11688
rect 36623 11685 36651 11716
rect 35437 11679 35495 11685
rect 35437 11676 35449 11679
rect 35216 11648 35449 11676
rect 35216 11636 35222 11648
rect 35437 11645 35449 11648
rect 35483 11676 35495 11679
rect 35989 11679 36047 11685
rect 35989 11676 36001 11679
rect 35483 11648 36001 11676
rect 35483 11645 35495 11648
rect 35437 11639 35495 11645
rect 35989 11645 36001 11648
rect 36035 11645 36047 11679
rect 35989 11639 36047 11645
rect 36608 11679 36666 11685
rect 36608 11645 36620 11679
rect 36654 11676 36666 11679
rect 37001 11679 37059 11685
rect 37001 11676 37013 11679
rect 36654 11648 37013 11676
rect 36654 11645 36666 11648
rect 36608 11639 36666 11645
rect 37001 11645 37013 11648
rect 37047 11645 37059 11679
rect 37001 11639 37059 11645
rect 33410 11608 33416 11620
rect 30484 11580 33416 11608
rect 22060 11568 22066 11580
rect 33410 11568 33416 11580
rect 33468 11568 33474 11620
rect 34606 11608 34612 11620
rect 33831 11580 34612 11608
rect 21269 11543 21327 11549
rect 21269 11509 21281 11543
rect 21315 11540 21327 11543
rect 21634 11540 21640 11552
rect 21315 11512 21640 11540
rect 21315 11509 21327 11512
rect 21269 11503 21327 11509
rect 21634 11500 21640 11512
rect 21692 11500 21698 11552
rect 24535 11543 24593 11549
rect 24535 11509 24547 11543
rect 24581 11540 24593 11543
rect 24670 11540 24676 11552
rect 24581 11512 24676 11540
rect 24581 11509 24593 11512
rect 24535 11503 24593 11509
rect 24670 11500 24676 11512
rect 24728 11500 24734 11552
rect 25406 11540 25412 11552
rect 25367 11512 25412 11540
rect 25406 11500 25412 11512
rect 25464 11500 25470 11552
rect 30147 11543 30205 11549
rect 30147 11509 30159 11543
rect 30193 11540 30205 11543
rect 30282 11540 30288 11552
rect 30193 11512 30288 11540
rect 30193 11509 30205 11512
rect 30147 11503 30205 11509
rect 30282 11500 30288 11512
rect 30340 11500 30346 11552
rect 31343 11543 31401 11549
rect 31343 11509 31355 11543
rect 31389 11540 31401 11543
rect 31478 11540 31484 11552
rect 31389 11512 31484 11540
rect 31389 11509 31401 11512
rect 31343 11503 31401 11509
rect 31478 11500 31484 11512
rect 31536 11500 31542 11552
rect 31846 11500 31852 11552
rect 31904 11540 31910 11552
rect 33831 11540 33859 11580
rect 34606 11568 34612 11580
rect 34664 11568 34670 11620
rect 31904 11512 33859 11540
rect 33919 11543 33977 11549
rect 31904 11500 31910 11512
rect 33919 11509 33931 11543
rect 33965 11540 33977 11543
rect 34882 11540 34888 11552
rect 33965 11512 34888 11540
rect 33965 11509 33977 11512
rect 33919 11503 33977 11509
rect 34882 11500 34888 11512
rect 34940 11500 34946 11552
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 2682 11336 2688 11348
rect 2643 11308 2688 11336
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 10134 11336 10140 11348
rect 10095 11308 10140 11336
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 15746 11336 15752 11348
rect 15707 11308 15752 11336
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 26651 11339 26709 11345
rect 26651 11305 26663 11339
rect 26697 11336 26709 11339
rect 27062 11336 27068 11348
rect 26697 11308 27068 11336
rect 26697 11305 26709 11308
rect 26651 11299 26709 11305
rect 27062 11296 27068 11308
rect 27120 11296 27126 11348
rect 31478 11336 31484 11348
rect 31439 11308 31484 11336
rect 31478 11296 31484 11308
rect 31536 11296 31542 11348
rect 35618 11336 35624 11348
rect 35579 11308 35624 11336
rect 35618 11296 35624 11308
rect 35676 11296 35682 11348
rect 11606 11268 11612 11280
rect 11567 11240 11612 11268
rect 11606 11228 11612 11240
rect 11664 11228 11670 11280
rect 20622 11228 20628 11280
rect 20680 11268 20686 11280
rect 21085 11271 21143 11277
rect 21085 11268 21097 11271
rect 20680 11240 21097 11268
rect 20680 11228 20686 11240
rect 21085 11237 21097 11240
rect 21131 11237 21143 11271
rect 24394 11268 24400 11280
rect 24355 11240 24400 11268
rect 21085 11231 21143 11237
rect 24394 11228 24400 11240
rect 24452 11228 24458 11280
rect 24486 11228 24492 11280
rect 24544 11268 24550 11280
rect 24544 11240 24589 11268
rect 24544 11228 24550 11240
rect 29546 11228 29552 11280
rect 29604 11268 29610 11280
rect 29825 11271 29883 11277
rect 29825 11268 29837 11271
rect 29604 11240 29837 11268
rect 29604 11228 29610 11240
rect 29825 11237 29837 11240
rect 29871 11237 29883 11271
rect 29825 11231 29883 11237
rect 29914 11228 29920 11280
rect 29972 11268 29978 11280
rect 29972 11240 30017 11268
rect 29972 11228 29978 11240
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 1670 11200 1676 11212
rect 1443 11172 1676 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 1670 11160 1676 11172
rect 1728 11160 1734 11212
rect 2501 11203 2559 11209
rect 2501 11169 2513 11203
rect 2547 11200 2559 11203
rect 3326 11200 3332 11212
rect 2547 11172 3332 11200
rect 2547 11169 2559 11172
rect 2501 11163 2559 11169
rect 3326 11160 3332 11172
rect 3384 11160 3390 11212
rect 4132 11203 4190 11209
rect 4132 11169 4144 11203
rect 4178 11200 4190 11203
rect 4706 11200 4712 11212
rect 4178 11172 4712 11200
rect 4178 11169 4190 11172
rect 4132 11163 4190 11169
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 8570 11200 8576 11212
rect 8531 11172 8576 11200
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 10042 11200 10048 11212
rect 10003 11172 10048 11200
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 10410 11200 10416 11212
rect 10371 11172 10416 11200
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 12986 11200 12992 11212
rect 12947 11172 12992 11200
rect 12986 11160 12992 11172
rect 13044 11160 13050 11212
rect 15470 11200 15476 11212
rect 15431 11172 15476 11200
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 15562 11160 15568 11212
rect 15620 11200 15626 11212
rect 15933 11203 15991 11209
rect 15933 11200 15945 11203
rect 15620 11172 15945 11200
rect 15620 11160 15626 11172
rect 15933 11169 15945 11172
rect 15979 11169 15991 11203
rect 15933 11163 15991 11169
rect 16482 11160 16488 11212
rect 16540 11200 16546 11212
rect 18208 11203 18266 11209
rect 18208 11200 18220 11203
rect 16540 11172 18220 11200
rect 16540 11160 16546 11172
rect 18208 11169 18220 11172
rect 18254 11200 18266 11203
rect 18322 11200 18328 11212
rect 18254 11172 18328 11200
rect 18254 11169 18266 11172
rect 18208 11163 18266 11169
rect 18322 11160 18328 11172
rect 18380 11160 18386 11212
rect 19150 11200 19156 11212
rect 19111 11172 19156 11200
rect 19150 11160 19156 11172
rect 19208 11160 19214 11212
rect 19610 11200 19616 11212
rect 19571 11172 19616 11200
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 23106 11160 23112 11212
rect 23164 11200 23170 11212
rect 23328 11203 23386 11209
rect 23328 11200 23340 11203
rect 23164 11172 23340 11200
rect 23164 11160 23170 11172
rect 23328 11169 23340 11172
rect 23374 11169 23386 11203
rect 23328 11163 23386 11169
rect 26580 11203 26638 11209
rect 26580 11169 26592 11203
rect 26626 11200 26638 11203
rect 27062 11200 27068 11212
rect 26626 11172 27068 11200
rect 26626 11169 26638 11172
rect 26580 11163 26638 11169
rect 27062 11160 27068 11172
rect 27120 11160 27126 11212
rect 27522 11160 27528 11212
rect 27580 11200 27586 11212
rect 27801 11203 27859 11209
rect 27801 11200 27813 11203
rect 27580 11172 27813 11200
rect 27580 11160 27586 11172
rect 27801 11169 27813 11172
rect 27847 11169 27859 11203
rect 27801 11163 27859 11169
rect 28074 11160 28080 11212
rect 28132 11200 28138 11212
rect 28261 11203 28319 11209
rect 28261 11200 28273 11203
rect 28132 11172 28273 11200
rect 28132 11160 28138 11172
rect 28261 11169 28273 11172
rect 28307 11169 28319 11203
rect 28261 11163 28319 11169
rect 31386 11160 31392 11212
rect 31444 11200 31450 11212
rect 32125 11203 32183 11209
rect 32125 11200 32137 11203
rect 31444 11172 32137 11200
rect 31444 11160 31450 11172
rect 32125 11169 32137 11172
rect 32171 11169 32183 11203
rect 32125 11163 32183 11169
rect 32490 11160 32496 11212
rect 32548 11200 32554 11212
rect 32585 11203 32643 11209
rect 32585 11200 32597 11203
rect 32548 11172 32597 11200
rect 32548 11160 32554 11172
rect 32585 11169 32597 11172
rect 32631 11169 32643 11203
rect 32585 11163 32643 11169
rect 34146 11160 34152 11212
rect 34204 11200 34210 11212
rect 34333 11203 34391 11209
rect 34333 11200 34345 11203
rect 34204 11172 34345 11200
rect 34204 11160 34210 11172
rect 34333 11169 34345 11172
rect 34379 11169 34391 11203
rect 35434 11200 35440 11212
rect 35395 11172 35440 11200
rect 34333 11163 34391 11169
rect 35434 11160 35440 11172
rect 35492 11160 35498 11212
rect 36541 11203 36599 11209
rect 36541 11169 36553 11203
rect 36587 11200 36599 11203
rect 36998 11200 37004 11212
rect 36587 11172 37004 11200
rect 36587 11169 36599 11172
rect 36541 11163 36599 11169
rect 36998 11160 37004 11172
rect 37056 11160 37062 11212
rect 11514 11132 11520 11144
rect 11475 11104 11520 11132
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 19886 11132 19892 11144
rect 11624 11104 13216 11132
rect 19847 11104 19892 11132
rect 8110 11024 8116 11076
rect 8168 11064 8174 11076
rect 11624 11064 11652 11104
rect 13188 11076 13216 11104
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 20993 11135 21051 11141
rect 20993 11101 21005 11135
rect 21039 11132 21051 11135
rect 21450 11132 21456 11144
rect 21039 11104 21456 11132
rect 21039 11101 21051 11104
rect 20993 11095 21051 11101
rect 21450 11092 21456 11104
rect 21508 11092 21514 11144
rect 21634 11132 21640 11144
rect 21595 11104 21640 11132
rect 21634 11092 21640 11104
rect 21692 11092 21698 11144
rect 25041 11135 25099 11141
rect 25041 11101 25053 11135
rect 25087 11132 25099 11135
rect 25222 11132 25228 11144
rect 25087 11104 25228 11132
rect 25087 11101 25099 11104
rect 25041 11095 25099 11101
rect 25222 11092 25228 11104
rect 25280 11092 25286 11144
rect 28537 11135 28595 11141
rect 28537 11101 28549 11135
rect 28583 11132 28595 11135
rect 29638 11132 29644 11144
rect 28583 11104 29644 11132
rect 28583 11101 28595 11104
rect 28537 11095 28595 11101
rect 29638 11092 29644 11104
rect 29696 11092 29702 11144
rect 32674 11132 32680 11144
rect 32635 11104 32680 11132
rect 32674 11092 32680 11104
rect 32732 11092 32738 11144
rect 34977 11135 35035 11141
rect 34977 11101 34989 11135
rect 35023 11132 35035 11135
rect 35066 11132 35072 11144
rect 35023 11104 35072 11132
rect 35023 11101 35035 11104
rect 34977 11095 35035 11101
rect 35066 11092 35072 11104
rect 35124 11092 35130 11144
rect 12066 11064 12072 11076
rect 8168 11036 11652 11064
rect 12027 11036 12072 11064
rect 8168 11024 8174 11036
rect 12066 11024 12072 11036
rect 12124 11024 12130 11076
rect 13170 11064 13176 11076
rect 13083 11036 13176 11064
rect 13170 11024 13176 11036
rect 13228 11024 13234 11076
rect 30377 11067 30435 11073
rect 30377 11033 30389 11067
rect 30423 11064 30435 11067
rect 30558 11064 30564 11076
rect 30423 11036 30564 11064
rect 30423 11033 30435 11036
rect 30377 11027 30435 11033
rect 30558 11024 30564 11036
rect 30616 11064 30622 11076
rect 33686 11064 33692 11076
rect 30616 11036 33692 11064
rect 30616 11024 30622 11036
rect 33686 11024 33692 11036
rect 33744 11064 33750 11076
rect 34422 11064 34428 11076
rect 33744 11036 34428 11064
rect 33744 11024 33750 11036
rect 34422 11024 34428 11036
rect 34480 11024 34486 11076
rect 34517 11067 34575 11073
rect 34517 11033 34529 11067
rect 34563 11064 34575 11067
rect 39574 11064 39580 11076
rect 34563 11036 39580 11064
rect 34563 11033 34575 11036
rect 34517 11027 34575 11033
rect 39574 11024 39580 11036
rect 39632 11024 39638 11076
rect 1578 10996 1584 11008
rect 1539 10968 1584 10996
rect 1578 10956 1584 10968
rect 1636 10956 1642 11008
rect 3786 10956 3792 11008
rect 3844 10996 3850 11008
rect 4203 10999 4261 11005
rect 4203 10996 4215 10999
rect 3844 10968 4215 10996
rect 3844 10956 3850 10968
rect 4203 10965 4215 10968
rect 4249 10965 4261 10999
rect 4203 10959 4261 10965
rect 8757 10999 8815 11005
rect 8757 10965 8769 10999
rect 8803 10996 8815 10999
rect 10042 10996 10048 11008
rect 8803 10968 10048 10996
rect 8803 10965 8815 10968
rect 8757 10959 8815 10965
rect 10042 10956 10048 10968
rect 10100 10956 10106 11008
rect 10226 10956 10232 11008
rect 10284 10996 10290 11008
rect 10873 10999 10931 11005
rect 10873 10996 10885 10999
rect 10284 10968 10885 10996
rect 10284 10956 10290 10968
rect 10873 10965 10885 10968
rect 10919 10965 10931 10999
rect 12434 10996 12440 11008
rect 12395 10968 12440 10996
rect 10873 10959 10931 10965
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 17586 10956 17592 11008
rect 17644 10996 17650 11008
rect 18279 10999 18337 11005
rect 18279 10996 18291 10999
rect 17644 10968 18291 10996
rect 17644 10956 17650 10968
rect 18279 10965 18291 10968
rect 18325 10965 18337 10999
rect 20162 10996 20168 11008
rect 20123 10968 20168 10996
rect 18279 10959 18337 10965
rect 20162 10956 20168 10968
rect 20220 10956 20226 11008
rect 23014 10956 23020 11008
rect 23072 10996 23078 11008
rect 23431 10999 23489 11005
rect 23431 10996 23443 10999
rect 23072 10968 23443 10996
rect 23072 10956 23078 10968
rect 23431 10965 23443 10968
rect 23477 10965 23489 10999
rect 23431 10959 23489 10965
rect 27709 10999 27767 11005
rect 27709 10965 27721 10999
rect 27755 10996 27767 10999
rect 28074 10996 28080 11008
rect 27755 10968 28080 10996
rect 27755 10965 27767 10968
rect 27709 10959 27767 10965
rect 28074 10956 28080 10968
rect 28132 10956 28138 11008
rect 34974 10956 34980 11008
rect 35032 10996 35038 11008
rect 35253 10999 35311 11005
rect 35253 10996 35265 10999
rect 35032 10968 35265 10996
rect 35032 10956 35038 10968
rect 35253 10965 35265 10968
rect 35299 10965 35311 10999
rect 36722 10996 36728 11008
rect 36683 10968 36728 10996
rect 35253 10959 35311 10965
rect 36722 10956 36728 10968
rect 36780 10956 36786 11008
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 4706 10792 4712 10804
rect 4667 10764 4712 10792
rect 4706 10752 4712 10764
rect 4764 10752 4770 10804
rect 8294 10792 8300 10804
rect 8255 10764 8300 10792
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 11517 10795 11575 10801
rect 11517 10761 11529 10795
rect 11563 10792 11575 10795
rect 11606 10792 11612 10804
rect 11563 10764 11612 10792
rect 11563 10761 11575 10764
rect 11517 10755 11575 10761
rect 11606 10752 11612 10764
rect 11664 10752 11670 10804
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 16482 10792 16488 10804
rect 11756 10764 16488 10792
rect 11756 10752 11762 10764
rect 16482 10752 16488 10764
rect 16540 10752 16546 10804
rect 16715 10795 16773 10801
rect 16715 10761 16727 10795
rect 16761 10792 16773 10795
rect 17126 10792 17132 10804
rect 16761 10764 17132 10792
rect 16761 10761 16773 10764
rect 16715 10755 16773 10761
rect 17126 10752 17132 10764
rect 17184 10752 17190 10804
rect 18322 10792 18328 10804
rect 18235 10764 18328 10792
rect 18322 10752 18328 10764
rect 18380 10792 18386 10804
rect 20809 10795 20867 10801
rect 20809 10792 20821 10795
rect 18380 10764 20821 10792
rect 18380 10752 18386 10764
rect 20809 10761 20821 10764
rect 20855 10761 20867 10795
rect 21450 10792 21456 10804
rect 21411 10764 21456 10792
rect 20809 10755 20867 10761
rect 21450 10752 21456 10764
rect 21508 10792 21514 10804
rect 23474 10792 23480 10804
rect 21508 10764 23480 10792
rect 21508 10752 21514 10764
rect 23474 10752 23480 10764
rect 23532 10752 23538 10804
rect 24029 10795 24087 10801
rect 24029 10761 24041 10795
rect 24075 10792 24087 10795
rect 24394 10792 24400 10804
rect 24075 10764 24400 10792
rect 24075 10761 24087 10764
rect 24029 10755 24087 10761
rect 24394 10752 24400 10764
rect 24452 10752 24458 10804
rect 27062 10792 27068 10804
rect 27023 10764 27068 10792
rect 27062 10752 27068 10764
rect 27120 10752 27126 10804
rect 29546 10752 29552 10804
rect 29604 10792 29610 10804
rect 29733 10795 29791 10801
rect 29733 10792 29745 10795
rect 29604 10764 29745 10792
rect 29604 10752 29610 10764
rect 29733 10761 29745 10764
rect 29779 10761 29791 10795
rect 29733 10755 29791 10761
rect 31754 10752 31760 10804
rect 31812 10792 31818 10804
rect 34146 10792 34152 10804
rect 31812 10764 34152 10792
rect 31812 10752 31818 10764
rect 34146 10752 34152 10764
rect 34204 10792 34210 10804
rect 34333 10795 34391 10801
rect 34333 10792 34345 10795
rect 34204 10764 34345 10792
rect 34204 10752 34210 10764
rect 34333 10761 34345 10764
rect 34379 10761 34391 10795
rect 36630 10792 36636 10804
rect 36591 10764 36636 10792
rect 34333 10755 34391 10761
rect 36630 10752 36636 10764
rect 36688 10752 36694 10804
rect 36998 10792 37004 10804
rect 36959 10764 37004 10792
rect 36998 10752 37004 10764
rect 37056 10752 37062 10804
rect 2406 10684 2412 10736
rect 2464 10724 2470 10736
rect 10045 10727 10103 10733
rect 2464 10696 9214 10724
rect 2464 10684 2470 10696
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1443 10560 2084 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 2056 10464 2084 10560
rect 2130 10548 2136 10600
rect 2188 10588 2194 10600
rect 2552 10591 2610 10597
rect 2552 10588 2564 10591
rect 2188 10560 2564 10588
rect 2188 10548 2194 10560
rect 2552 10557 2564 10560
rect 2598 10588 2610 10591
rect 3948 10591 4006 10597
rect 2598 10557 2611 10588
rect 2552 10551 2611 10557
rect 3948 10557 3960 10591
rect 3994 10588 4006 10591
rect 8113 10591 8171 10597
rect 3994 10560 4154 10588
rect 3994 10557 4006 10560
rect 3948 10551 4006 10557
rect 106 10412 112 10464
rect 164 10452 170 10464
rect 1581 10455 1639 10461
rect 1581 10452 1593 10455
rect 164 10424 1593 10452
rect 164 10412 170 10424
rect 1581 10421 1593 10424
rect 1627 10421 1639 10455
rect 2038 10452 2044 10464
rect 1999 10424 2044 10452
rect 1581 10415 1639 10421
rect 2038 10412 2044 10424
rect 2096 10412 2102 10464
rect 2583 10452 2611 10551
rect 2639 10523 2697 10529
rect 2639 10489 2651 10523
rect 2685 10520 2697 10523
rect 3418 10520 3424 10532
rect 2685 10492 3424 10520
rect 2685 10489 2697 10492
rect 2639 10483 2697 10489
rect 3418 10480 3424 10492
rect 3476 10480 3482 10532
rect 3053 10455 3111 10461
rect 3053 10452 3065 10455
rect 2583 10424 3065 10452
rect 3053 10421 3065 10424
rect 3099 10452 3111 10455
rect 3142 10452 3148 10464
rect 3099 10424 3148 10452
rect 3099 10421 3111 10424
rect 3053 10415 3111 10421
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 3326 10452 3332 10464
rect 3287 10424 3332 10452
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 3878 10412 3884 10464
rect 3936 10452 3942 10464
rect 4019 10455 4077 10461
rect 4019 10452 4031 10455
rect 3936 10424 4031 10452
rect 3936 10412 3942 10424
rect 4019 10421 4031 10424
rect 4065 10421 4077 10455
rect 4126 10452 4154 10560
rect 8113 10557 8125 10591
rect 8159 10588 8171 10591
rect 8202 10588 8208 10600
rect 8159 10560 8208 10588
rect 8159 10557 8171 10560
rect 8113 10551 8171 10557
rect 8202 10548 8208 10560
rect 8260 10588 8266 10600
rect 9186 10597 9214 10696
rect 10045 10693 10057 10727
rect 10091 10724 10103 10727
rect 10410 10724 10416 10736
rect 10091 10696 10416 10724
rect 10091 10693 10103 10696
rect 10045 10687 10103 10693
rect 10410 10684 10416 10696
rect 10468 10724 10474 10736
rect 10468 10696 12296 10724
rect 10468 10684 10474 10696
rect 9263 10659 9321 10665
rect 9263 10625 9275 10659
rect 9309 10656 9321 10659
rect 11514 10656 11520 10668
rect 9309 10628 11520 10656
rect 9309 10625 9321 10628
rect 9263 10619 9321 10625
rect 11514 10616 11520 10628
rect 11572 10656 11578 10668
rect 12268 10665 12296 10696
rect 12986 10684 12992 10736
rect 13044 10724 13050 10736
rect 13449 10727 13507 10733
rect 13449 10724 13461 10727
rect 13044 10696 13461 10724
rect 13044 10684 13050 10696
rect 13449 10693 13461 10696
rect 13495 10693 13507 10727
rect 19150 10724 19156 10736
rect 13449 10687 13507 10693
rect 13786 10696 19156 10724
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 11572 10628 11805 10656
rect 11572 10616 11578 10628
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 11793 10619 11851 10625
rect 12253 10659 12311 10665
rect 12253 10625 12265 10659
rect 12299 10656 12311 10659
rect 12299 10628 13032 10656
rect 12299 10625 12311 10628
rect 12253 10619 12311 10625
rect 8573 10591 8631 10597
rect 8573 10588 8585 10591
rect 8260 10560 8585 10588
rect 8260 10548 8266 10560
rect 8573 10557 8585 10560
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 9176 10591 9234 10597
rect 9176 10557 9188 10591
rect 9222 10588 9234 10591
rect 12434 10588 12440 10600
rect 9222 10560 9720 10588
rect 12395 10560 12440 10588
rect 9222 10557 9234 10560
rect 9176 10551 9234 10557
rect 9692 10464 9720 10560
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 13004 10597 13032 10628
rect 13170 10616 13176 10668
rect 13228 10656 13234 10668
rect 13786 10656 13814 10696
rect 19150 10684 19156 10696
rect 19208 10724 19214 10736
rect 19797 10727 19855 10733
rect 19797 10724 19809 10727
rect 19208 10696 19809 10724
rect 19208 10684 19214 10696
rect 19797 10693 19809 10696
rect 19843 10724 19855 10727
rect 21266 10724 21272 10736
rect 19843 10696 21272 10724
rect 19843 10693 19855 10696
rect 19797 10687 19855 10693
rect 21266 10684 21272 10696
rect 21324 10724 21330 10736
rect 29089 10727 29147 10733
rect 21324 10696 26188 10724
rect 21324 10684 21330 10696
rect 15378 10656 15384 10668
rect 13228 10628 13814 10656
rect 15339 10628 15384 10656
rect 13228 10616 13234 10628
rect 15378 10616 15384 10628
rect 15436 10656 15442 10668
rect 19518 10656 19524 10668
rect 15436 10628 16655 10656
rect 15436 10616 15442 10628
rect 12989 10591 13047 10597
rect 12989 10557 13001 10591
rect 13035 10588 13047 10591
rect 14182 10588 14188 10600
rect 13035 10560 14188 10588
rect 13035 10557 13047 10560
rect 12989 10551 13047 10557
rect 14182 10548 14188 10560
rect 14240 10548 14246 10600
rect 16627 10597 16655 10628
rect 18708 10628 19524 10656
rect 18708 10597 18736 10628
rect 19518 10616 19524 10628
rect 19576 10616 19582 10668
rect 19702 10616 19708 10668
rect 19760 10656 19766 10668
rect 20070 10656 20076 10668
rect 19760 10628 20076 10656
rect 19760 10616 19766 10628
rect 20070 10616 20076 10628
rect 20128 10616 20134 10668
rect 20717 10659 20775 10665
rect 20717 10625 20729 10659
rect 20763 10656 20775 10659
rect 21634 10656 21640 10668
rect 20763 10628 21640 10656
rect 20763 10625 20775 10628
rect 20717 10619 20775 10625
rect 21634 10616 21640 10628
rect 21692 10616 21698 10668
rect 24578 10656 24584 10668
rect 24539 10628 24584 10656
rect 24578 10616 24584 10628
rect 24636 10656 24642 10668
rect 25501 10659 25559 10665
rect 25501 10656 25513 10659
rect 24636 10628 25513 10656
rect 24636 10616 24642 10628
rect 25501 10625 25513 10628
rect 25547 10625 25559 10659
rect 25501 10619 25559 10625
rect 16612 10591 16670 10597
rect 16612 10557 16624 10591
rect 16658 10588 16670 10591
rect 17037 10591 17095 10597
rect 17037 10588 17049 10591
rect 16658 10560 17049 10588
rect 16658 10557 16670 10560
rect 16612 10551 16670 10557
rect 17037 10557 17049 10560
rect 17083 10557 17095 10591
rect 17037 10551 17095 10557
rect 17865 10591 17923 10597
rect 17865 10557 17877 10591
rect 17911 10588 17923 10591
rect 18693 10591 18751 10597
rect 18693 10588 18705 10591
rect 17911 10560 18705 10588
rect 17911 10557 17923 10560
rect 17865 10551 17923 10557
rect 18693 10557 18705 10560
rect 18739 10557 18751 10591
rect 18693 10551 18751 10557
rect 18969 10591 19027 10597
rect 18969 10557 18981 10591
rect 19015 10588 19027 10591
rect 19015 10560 19564 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 10226 10520 10232 10532
rect 10187 10492 10232 10520
rect 10226 10480 10232 10492
rect 10284 10480 10290 10532
rect 10318 10480 10324 10532
rect 10376 10520 10382 10532
rect 10873 10523 10931 10529
rect 10376 10492 10421 10520
rect 10376 10480 10382 10492
rect 10873 10489 10885 10523
rect 10919 10520 10931 10523
rect 11054 10520 11060 10532
rect 10919 10492 11060 10520
rect 10919 10489 10931 10492
rect 10873 10483 10931 10489
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 15102 10520 15108 10532
rect 15063 10492 15108 10520
rect 15102 10480 15108 10492
rect 15160 10480 15166 10532
rect 15194 10480 15200 10532
rect 15252 10520 15258 10532
rect 15252 10492 15297 10520
rect 15252 10480 15258 10492
rect 15470 10480 15476 10532
rect 15528 10520 15534 10532
rect 16117 10523 16175 10529
rect 16117 10520 16129 10523
rect 15528 10492 16129 10520
rect 15528 10480 15534 10492
rect 16117 10489 16129 10492
rect 16163 10520 16175 10523
rect 17880 10520 17908 10551
rect 19150 10520 19156 10532
rect 16163 10492 17908 10520
rect 19111 10492 19156 10520
rect 16163 10489 16175 10492
rect 16117 10483 16175 10489
rect 19150 10480 19156 10492
rect 19208 10480 19214 10532
rect 4338 10452 4344 10464
rect 4126 10424 4344 10452
rect 4019 10415 4077 10421
rect 4338 10412 4344 10424
rect 4396 10412 4402 10464
rect 6546 10412 6552 10464
rect 6604 10452 6610 10464
rect 6825 10455 6883 10461
rect 6825 10452 6837 10455
rect 6604 10424 6837 10452
rect 6604 10412 6610 10424
rect 6825 10421 6837 10424
rect 6871 10421 6883 10455
rect 6825 10415 6883 10421
rect 7282 10412 7288 10464
rect 7340 10452 7346 10464
rect 8570 10452 8576 10464
rect 7340 10424 8576 10452
rect 7340 10412 7346 10424
rect 8570 10412 8576 10424
rect 8628 10452 8634 10464
rect 8941 10455 8999 10461
rect 8941 10452 8953 10455
rect 8628 10424 8953 10452
rect 8628 10412 8634 10424
rect 8941 10421 8953 10424
rect 8987 10421 8999 10455
rect 9674 10452 9680 10464
rect 9635 10424 9680 10452
rect 8941 10415 8999 10421
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 12526 10452 12532 10464
rect 12487 10424 12532 10452
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 14001 10455 14059 10461
rect 14001 10421 14013 10455
rect 14047 10452 14059 10455
rect 14826 10452 14832 10464
rect 14047 10424 14832 10452
rect 14047 10421 14059 10424
rect 14001 10415 14059 10421
rect 14826 10412 14832 10424
rect 14884 10412 14890 10464
rect 14921 10455 14979 10461
rect 14921 10421 14933 10455
rect 14967 10452 14979 10455
rect 15212 10452 15240 10480
rect 19536 10461 19564 10560
rect 21450 10548 21456 10600
rect 21508 10588 21514 10600
rect 21545 10591 21603 10597
rect 21545 10588 21557 10591
rect 21508 10560 21557 10588
rect 21508 10548 21514 10560
rect 21545 10557 21557 10560
rect 21591 10588 21603 10591
rect 22005 10591 22063 10597
rect 22005 10588 22017 10591
rect 21591 10560 22017 10588
rect 21591 10557 21603 10560
rect 21545 10551 21603 10557
rect 22005 10557 22017 10560
rect 22051 10557 22063 10591
rect 22005 10551 22063 10557
rect 22608 10591 22666 10597
rect 22608 10557 22620 10591
rect 22654 10588 22666 10591
rect 22830 10588 22836 10600
rect 22654 10560 22836 10588
rect 22654 10557 22666 10560
rect 22608 10551 22666 10557
rect 22830 10548 22836 10560
rect 22888 10588 22894 10600
rect 26160 10597 26188 10696
rect 29089 10693 29101 10727
rect 29135 10724 29147 10727
rect 29454 10724 29460 10736
rect 29135 10696 29460 10724
rect 29135 10693 29147 10696
rect 29089 10687 29147 10693
rect 29454 10684 29460 10696
rect 29512 10724 29518 10736
rect 29914 10724 29920 10736
rect 29512 10696 29920 10724
rect 29512 10684 29518 10696
rect 29914 10684 29920 10696
rect 29972 10684 29978 10736
rect 30558 10724 30564 10736
rect 30519 10696 30564 10724
rect 30558 10684 30564 10696
rect 30616 10684 30622 10736
rect 31478 10684 31484 10736
rect 31536 10724 31542 10736
rect 31536 10696 31616 10724
rect 31536 10684 31542 10696
rect 30006 10656 30012 10668
rect 27908 10628 30012 10656
rect 23017 10591 23075 10597
rect 23017 10588 23029 10591
rect 22888 10560 23029 10588
rect 22888 10548 22894 10560
rect 23017 10557 23029 10560
rect 23063 10557 23075 10591
rect 23017 10551 23075 10557
rect 26145 10591 26203 10597
rect 26145 10557 26157 10591
rect 26191 10557 26203 10591
rect 26145 10551 26203 10557
rect 20162 10480 20168 10532
rect 20220 10520 20226 10532
rect 20809 10523 20867 10529
rect 20220 10492 20265 10520
rect 20220 10480 20226 10492
rect 20809 10489 20821 10523
rect 20855 10520 20867 10523
rect 22695 10523 22753 10529
rect 20855 10492 21858 10520
rect 20855 10489 20867 10492
rect 20809 10483 20867 10489
rect 14967 10424 15240 10452
rect 19521 10455 19579 10461
rect 14967 10421 14979 10424
rect 14921 10415 14979 10421
rect 19521 10421 19533 10455
rect 19567 10452 19579 10455
rect 19702 10452 19708 10464
rect 19567 10424 19708 10452
rect 19567 10421 19579 10424
rect 19521 10415 19579 10421
rect 19702 10412 19708 10424
rect 19760 10412 19766 10464
rect 20622 10412 20628 10464
rect 20680 10452 20686 10464
rect 20993 10455 21051 10461
rect 20993 10452 21005 10455
rect 20680 10424 21005 10452
rect 20680 10412 20686 10424
rect 20993 10421 21005 10424
rect 21039 10421 21051 10455
rect 21726 10452 21732 10464
rect 21687 10424 21732 10452
rect 20993 10415 21051 10421
rect 21726 10412 21732 10424
rect 21784 10412 21790 10464
rect 21830 10452 21858 10492
rect 22695 10489 22707 10523
rect 22741 10520 22753 10523
rect 23290 10520 23296 10532
rect 22741 10492 23296 10520
rect 22741 10489 22753 10492
rect 22695 10483 22753 10489
rect 23290 10480 23296 10492
rect 23348 10480 23354 10532
rect 24578 10480 24584 10532
rect 24636 10520 24642 10532
rect 24673 10523 24731 10529
rect 24673 10520 24685 10523
rect 24636 10492 24685 10520
rect 24636 10480 24642 10492
rect 24673 10489 24685 10492
rect 24719 10489 24731 10523
rect 25222 10520 25228 10532
rect 25183 10492 25228 10520
rect 24673 10483 24731 10489
rect 25222 10480 25228 10492
rect 25280 10480 25286 10532
rect 25961 10523 26019 10529
rect 25961 10489 25973 10523
rect 26007 10520 26019 10523
rect 26160 10520 26188 10551
rect 26234 10548 26240 10600
rect 26292 10588 26298 10600
rect 27908 10597 27936 10628
rect 30006 10616 30012 10628
rect 30064 10616 30070 10668
rect 31588 10665 31616 10696
rect 34054 10684 34060 10736
rect 34112 10724 34118 10736
rect 36265 10727 36323 10733
rect 36265 10724 36277 10727
rect 34112 10696 36277 10724
rect 34112 10684 34118 10696
rect 36265 10693 36277 10696
rect 36311 10693 36323 10727
rect 36265 10687 36323 10693
rect 31573 10659 31631 10665
rect 31573 10625 31585 10659
rect 31619 10625 31631 10659
rect 31573 10619 31631 10625
rect 32490 10616 32496 10668
rect 32548 10656 32554 10668
rect 33318 10656 33324 10668
rect 32548 10628 33324 10656
rect 32548 10616 32554 10628
rect 33318 10616 33324 10628
rect 33376 10656 33382 10668
rect 33376 10628 33548 10656
rect 33376 10616 33382 10628
rect 26513 10591 26571 10597
rect 26513 10588 26525 10591
rect 26292 10560 26525 10588
rect 26292 10548 26298 10560
rect 26513 10557 26525 10560
rect 26559 10557 26571 10591
rect 26513 10551 26571 10557
rect 27525 10591 27583 10597
rect 27525 10557 27537 10591
rect 27571 10588 27583 10591
rect 27893 10591 27951 10597
rect 27893 10588 27905 10591
rect 27571 10560 27905 10588
rect 27571 10557 27583 10560
rect 27525 10551 27583 10557
rect 27893 10557 27905 10560
rect 27939 10557 27951 10591
rect 28074 10588 28080 10600
rect 28035 10560 28080 10588
rect 27893 10551 27951 10557
rect 27540 10520 27568 10551
rect 28074 10548 28080 10560
rect 28132 10548 28138 10600
rect 32950 10588 32956 10600
rect 32863 10560 32956 10588
rect 32950 10548 32956 10560
rect 33008 10588 33014 10600
rect 33520 10597 33548 10628
rect 34146 10616 34152 10668
rect 34204 10656 34210 10668
rect 35434 10656 35440 10668
rect 34204 10628 35440 10656
rect 34204 10616 34210 10628
rect 35434 10616 35440 10628
rect 35492 10656 35498 10668
rect 35897 10659 35955 10665
rect 35897 10656 35909 10659
rect 35492 10628 35909 10656
rect 35492 10616 35498 10628
rect 35897 10625 35909 10628
rect 35943 10625 35955 10659
rect 35897 10619 35955 10625
rect 33045 10591 33103 10597
rect 33045 10588 33057 10591
rect 33008 10560 33057 10588
rect 33008 10548 33014 10560
rect 33045 10557 33057 10560
rect 33091 10557 33103 10591
rect 33045 10551 33103 10557
rect 33505 10591 33563 10597
rect 33505 10557 33517 10591
rect 33551 10557 33563 10591
rect 33778 10588 33784 10600
rect 33739 10560 33784 10588
rect 33505 10551 33563 10557
rect 33778 10548 33784 10560
rect 33836 10548 33842 10600
rect 36280 10588 36308 10687
rect 36449 10591 36507 10597
rect 36449 10588 36461 10591
rect 36280 10560 36461 10588
rect 36449 10557 36461 10560
rect 36495 10557 36507 10591
rect 36449 10551 36507 10557
rect 37604 10591 37662 10597
rect 37604 10557 37616 10591
rect 37650 10588 37662 10591
rect 37650 10560 37872 10588
rect 37650 10557 37662 10560
rect 37604 10551 37662 10557
rect 28350 10520 28356 10532
rect 26007 10492 27568 10520
rect 28311 10492 28356 10520
rect 26007 10489 26019 10492
rect 25961 10483 26019 10489
rect 28350 10480 28356 10492
rect 28408 10480 28414 10532
rect 30009 10523 30067 10529
rect 30009 10489 30021 10523
rect 30055 10489 30067 10523
rect 30009 10483 30067 10489
rect 23106 10452 23112 10464
rect 21830 10424 23112 10452
rect 23106 10412 23112 10424
rect 23164 10452 23170 10464
rect 23385 10455 23443 10461
rect 23385 10452 23397 10455
rect 23164 10424 23397 10452
rect 23164 10412 23170 10424
rect 23385 10421 23397 10424
rect 23431 10421 23443 10455
rect 24394 10452 24400 10464
rect 24355 10424 24400 10452
rect 23385 10415 23443 10421
rect 24394 10412 24400 10424
rect 24452 10412 24458 10464
rect 26142 10452 26148 10464
rect 26103 10424 26148 10452
rect 26142 10412 26148 10424
rect 26200 10412 26206 10464
rect 27522 10412 27528 10464
rect 27580 10452 27586 10464
rect 28629 10455 28687 10461
rect 28629 10452 28641 10455
rect 27580 10424 28641 10452
rect 27580 10412 27586 10424
rect 28629 10421 28641 10424
rect 28675 10421 28687 10455
rect 30024 10452 30052 10483
rect 30098 10480 30104 10532
rect 30156 10520 30162 10532
rect 30156 10492 30201 10520
rect 30156 10480 30162 10492
rect 30650 10480 30656 10532
rect 30708 10520 30714 10532
rect 31297 10523 31355 10529
rect 31297 10520 31309 10523
rect 30708 10492 31309 10520
rect 30708 10480 30714 10492
rect 31297 10489 31309 10492
rect 31343 10520 31355 10523
rect 31386 10520 31392 10532
rect 31343 10492 31392 10520
rect 31343 10489 31355 10492
rect 31297 10483 31355 10489
rect 31386 10480 31392 10492
rect 31444 10480 31450 10532
rect 31662 10520 31668 10532
rect 31623 10492 31668 10520
rect 31662 10480 31668 10492
rect 31720 10480 31726 10532
rect 32214 10520 32220 10532
rect 32175 10492 32220 10520
rect 32214 10480 32220 10492
rect 32272 10480 32278 10532
rect 32306 10480 32312 10532
rect 32364 10520 32370 10532
rect 34974 10520 34980 10532
rect 32364 10492 34980 10520
rect 32364 10480 32370 10492
rect 34974 10480 34980 10492
rect 35032 10480 35038 10532
rect 35066 10480 35072 10532
rect 35124 10520 35130 10532
rect 35618 10520 35624 10532
rect 35124 10492 35169 10520
rect 35579 10492 35624 10520
rect 35124 10480 35130 10492
rect 35618 10480 35624 10492
rect 35676 10480 35682 10532
rect 37691 10523 37749 10529
rect 37691 10520 37703 10523
rect 35820 10492 37703 10520
rect 31021 10455 31079 10461
rect 31021 10452 31033 10455
rect 30024 10424 31033 10452
rect 28629 10415 28687 10421
rect 31021 10421 31033 10424
rect 31067 10452 31079 10455
rect 31110 10452 31116 10464
rect 31067 10424 31116 10452
rect 31067 10421 31079 10424
rect 31021 10415 31079 10421
rect 31110 10412 31116 10424
rect 31168 10412 31174 10464
rect 32490 10452 32496 10464
rect 32451 10424 32496 10452
rect 32490 10412 32496 10424
rect 32548 10412 32554 10464
rect 34606 10412 34612 10464
rect 34664 10452 34670 10464
rect 35820 10452 35848 10492
rect 37691 10489 37703 10492
rect 37737 10489 37749 10523
rect 37691 10483 37749 10489
rect 34664 10424 35848 10452
rect 34664 10412 34670 10424
rect 36078 10412 36084 10464
rect 36136 10452 36142 10464
rect 37844 10452 37872 10560
rect 38013 10455 38071 10461
rect 38013 10452 38025 10455
rect 36136 10424 38025 10452
rect 36136 10412 36142 10424
rect 38013 10421 38025 10424
rect 38059 10421 38071 10455
rect 38013 10415 38071 10421
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 1762 10208 1768 10260
rect 1820 10248 1826 10260
rect 2041 10251 2099 10257
rect 2041 10248 2053 10251
rect 1820 10220 2053 10248
rect 1820 10208 1826 10220
rect 2041 10217 2053 10220
rect 2087 10217 2099 10251
rect 2041 10211 2099 10217
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 4939 10251 4997 10257
rect 4939 10248 4951 10251
rect 2832 10220 4951 10248
rect 2832 10208 2838 10220
rect 4939 10217 4951 10220
rect 4985 10217 4997 10251
rect 10318 10248 10324 10260
rect 10279 10220 10324 10248
rect 4939 10211 4997 10217
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 11606 10208 11612 10260
rect 11664 10248 11670 10260
rect 11664 10220 12204 10248
rect 11664 10208 11670 10220
rect 10594 10180 10600 10192
rect 10555 10152 10600 10180
rect 10594 10140 10600 10152
rect 10652 10140 10658 10192
rect 11422 10140 11428 10192
rect 11480 10180 11486 10192
rect 12176 10189 12204 10220
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 13725 10251 13783 10257
rect 13725 10248 13737 10251
rect 13688 10220 13737 10248
rect 13688 10208 13694 10220
rect 13725 10217 13737 10220
rect 13771 10217 13783 10251
rect 19061 10251 19119 10257
rect 13725 10211 13783 10217
rect 14016 10220 16160 10248
rect 12069 10183 12127 10189
rect 12069 10180 12081 10183
rect 11480 10152 12081 10180
rect 11480 10140 11486 10152
rect 12069 10149 12081 10152
rect 12115 10149 12127 10183
rect 12069 10143 12127 10149
rect 12161 10183 12219 10189
rect 12161 10149 12173 10183
rect 12207 10149 12219 10183
rect 12161 10143 12219 10149
rect 1486 10072 1492 10124
rect 1544 10112 1550 10124
rect 1949 10115 2007 10121
rect 1949 10112 1961 10115
rect 1544 10084 1961 10112
rect 1544 10072 1550 10084
rect 1949 10081 1961 10084
rect 1995 10081 2007 10115
rect 2406 10112 2412 10124
rect 2367 10084 2412 10112
rect 1949 10075 2007 10081
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 4868 10115 4926 10121
rect 4868 10081 4880 10115
rect 4914 10112 4926 10115
rect 5166 10112 5172 10124
rect 4914 10084 5172 10112
rect 4914 10081 4926 10084
rect 4868 10075 4926 10081
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 7628 10115 7686 10121
rect 7628 10081 7640 10115
rect 7674 10112 7686 10115
rect 8018 10112 8024 10124
rect 7674 10084 8024 10112
rect 7674 10081 7686 10084
rect 7628 10075 7686 10081
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 8608 10115 8666 10121
rect 8608 10112 8620 10115
rect 8444 10084 8620 10112
rect 8444 10072 8450 10084
rect 8608 10081 8620 10084
rect 8654 10081 8666 10115
rect 8608 10075 8666 10081
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 13909 10115 13967 10121
rect 13909 10112 13921 10115
rect 13872 10084 13921 10112
rect 13872 10072 13878 10084
rect 13909 10081 13921 10084
rect 13955 10112 13967 10115
rect 14016 10112 14044 10220
rect 15562 10140 15568 10192
rect 15620 10180 15626 10192
rect 16022 10180 16028 10192
rect 15620 10152 15700 10180
rect 15983 10152 16028 10180
rect 15620 10140 15626 10152
rect 14182 10112 14188 10124
rect 13955 10084 14044 10112
rect 14095 10084 14188 10112
rect 13955 10081 13967 10084
rect 13909 10075 13967 10081
rect 14182 10072 14188 10084
rect 14240 10112 14246 10124
rect 15672 10112 15700 10152
rect 16022 10140 16028 10152
rect 16080 10140 16086 10192
rect 16132 10180 16160 10220
rect 19061 10217 19073 10251
rect 19107 10248 19119 10251
rect 19150 10248 19156 10260
rect 19107 10220 19156 10248
rect 19107 10217 19119 10220
rect 19061 10211 19119 10217
rect 19150 10208 19156 10220
rect 19208 10208 19214 10260
rect 19242 10208 19248 10260
rect 19300 10248 19306 10260
rect 19300 10220 19345 10248
rect 19300 10208 19306 10220
rect 20070 10208 20076 10260
rect 20128 10248 20134 10260
rect 20165 10251 20223 10257
rect 20165 10248 20177 10251
rect 20128 10220 20177 10248
rect 20128 10208 20134 10220
rect 20165 10217 20177 10220
rect 20211 10217 20223 10251
rect 25222 10248 25228 10260
rect 20165 10211 20223 10217
rect 22940 10220 25228 10248
rect 21085 10183 21143 10189
rect 16132 10152 19472 10180
rect 17678 10112 17684 10124
rect 14240 10084 15700 10112
rect 17639 10084 17684 10112
rect 14240 10072 14246 10084
rect 17678 10072 17684 10084
rect 17736 10072 17742 10124
rect 18138 10112 18144 10124
rect 18099 10084 18144 10112
rect 18138 10072 18144 10084
rect 18196 10072 18202 10124
rect 19444 10121 19472 10152
rect 21085 10149 21097 10183
rect 21131 10180 21143 10183
rect 21910 10180 21916 10192
rect 21131 10152 21916 10180
rect 21131 10149 21143 10152
rect 21085 10143 21143 10149
rect 21910 10140 21916 10152
rect 21968 10140 21974 10192
rect 19429 10115 19487 10121
rect 19429 10081 19441 10115
rect 19475 10112 19487 10115
rect 19518 10112 19524 10124
rect 19475 10084 19524 10112
rect 19475 10081 19487 10084
rect 19429 10075 19487 10081
rect 19518 10072 19524 10084
rect 19576 10072 19582 10124
rect 19702 10112 19708 10124
rect 19663 10084 19708 10112
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 21634 10072 21640 10124
rect 21692 10112 21698 10124
rect 21692 10084 21737 10112
rect 21692 10072 21698 10084
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 9582 10044 9588 10056
rect 6595 10016 9588 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 9582 10004 9588 10016
rect 9640 10004 9646 10056
rect 10502 10044 10508 10056
rect 10463 10016 10508 10044
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 12342 10044 12348 10056
rect 12303 10016 12348 10044
rect 12342 10004 12348 10016
rect 12400 10044 12406 10056
rect 15013 10047 15071 10053
rect 15013 10044 15025 10047
rect 12400 10016 15025 10044
rect 12400 10004 12406 10016
rect 15013 10013 15025 10016
rect 15059 10044 15071 10047
rect 15102 10044 15108 10056
rect 15059 10016 15108 10044
rect 15059 10013 15071 10016
rect 15013 10007 15071 10013
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 15930 10044 15936 10056
rect 15891 10016 15936 10044
rect 15930 10004 15936 10016
rect 15988 10004 15994 10056
rect 16209 10047 16267 10053
rect 16209 10013 16221 10047
rect 16255 10013 16267 10047
rect 18322 10044 18328 10056
rect 18283 10016 18328 10044
rect 16209 10007 16267 10013
rect 7699 9979 7757 9985
rect 7699 9945 7711 9979
rect 7745 9976 7757 9979
rect 10962 9976 10968 9988
rect 7745 9948 10968 9976
rect 7745 9945 7757 9948
rect 7699 9939 7757 9945
rect 10962 9936 10968 9948
rect 11020 9936 11026 9988
rect 11054 9936 11060 9988
rect 11112 9976 11118 9988
rect 12066 9976 12072 9988
rect 11112 9948 12072 9976
rect 11112 9936 11118 9948
rect 12066 9936 12072 9948
rect 12124 9976 12130 9988
rect 13170 9976 13176 9988
rect 12124 9948 13176 9976
rect 12124 9936 12130 9948
rect 13170 9936 13176 9948
rect 13228 9936 13234 9988
rect 15378 9936 15384 9988
rect 15436 9976 15442 9988
rect 16224 9976 16252 10007
rect 18322 10004 18328 10016
rect 18380 10004 18386 10056
rect 18693 10047 18751 10053
rect 18693 10013 18705 10047
rect 18739 10044 18751 10047
rect 19720 10044 19748 10072
rect 18739 10016 19748 10044
rect 18739 10013 18751 10016
rect 18693 10007 18751 10013
rect 20714 10004 20720 10056
rect 20772 10044 20778 10056
rect 20993 10047 21051 10053
rect 20993 10044 21005 10047
rect 20772 10016 21005 10044
rect 20772 10004 20778 10016
rect 20993 10013 21005 10016
rect 21039 10044 21051 10047
rect 22940 10044 22968 10220
rect 25222 10208 25228 10220
rect 25280 10248 25286 10260
rect 29454 10248 29460 10260
rect 25280 10220 25452 10248
rect 29415 10220 29460 10248
rect 25280 10208 25286 10220
rect 23198 10140 23204 10192
rect 23256 10180 23262 10192
rect 23293 10183 23351 10189
rect 23293 10180 23305 10183
rect 23256 10152 23305 10180
rect 23256 10140 23262 10152
rect 23293 10149 23305 10152
rect 23339 10180 23351 10183
rect 24489 10183 24547 10189
rect 24489 10180 24501 10183
rect 23339 10152 24501 10180
rect 23339 10149 23351 10152
rect 23293 10143 23351 10149
rect 24489 10149 24501 10152
rect 24535 10180 24547 10183
rect 24578 10180 24584 10192
rect 24535 10152 24584 10180
rect 24535 10149 24547 10152
rect 24489 10143 24547 10149
rect 24578 10140 24584 10152
rect 24636 10140 24642 10192
rect 24762 10180 24768 10192
rect 24723 10152 24768 10180
rect 24762 10140 24768 10152
rect 24820 10140 24826 10192
rect 24854 10140 24860 10192
rect 24912 10180 24918 10192
rect 25424 10189 25452 10220
rect 29454 10208 29460 10220
rect 29512 10208 29518 10260
rect 29638 10208 29644 10260
rect 29696 10248 29702 10260
rect 29733 10251 29791 10257
rect 29733 10248 29745 10251
rect 29696 10220 29745 10248
rect 29696 10208 29702 10220
rect 29733 10217 29745 10220
rect 29779 10217 29791 10251
rect 31573 10251 31631 10257
rect 31573 10248 31585 10251
rect 29733 10211 29791 10217
rect 30576 10220 31585 10248
rect 30576 10192 30604 10220
rect 31573 10217 31585 10220
rect 31619 10248 31631 10251
rect 31662 10248 31668 10260
rect 31619 10220 31668 10248
rect 31619 10217 31631 10220
rect 31573 10211 31631 10217
rect 31662 10208 31668 10220
rect 31720 10208 31726 10260
rect 32674 10248 32680 10260
rect 32635 10220 32680 10248
rect 32674 10208 32680 10220
rect 32732 10208 32738 10260
rect 33873 10251 33931 10257
rect 33873 10248 33885 10251
rect 33060 10220 33885 10248
rect 25409 10183 25467 10189
rect 24912 10152 24957 10180
rect 24912 10140 24918 10152
rect 25409 10149 25421 10183
rect 25455 10149 25467 10183
rect 25409 10143 25467 10149
rect 25958 10140 25964 10192
rect 26016 10180 26022 10192
rect 26697 10183 26755 10189
rect 26697 10180 26709 10183
rect 26016 10152 26709 10180
rect 26016 10140 26022 10152
rect 26697 10149 26709 10152
rect 26743 10149 26755 10183
rect 26697 10143 26755 10149
rect 28626 10140 28632 10192
rect 28684 10180 28690 10192
rect 28858 10183 28916 10189
rect 28858 10180 28870 10183
rect 28684 10152 28870 10180
rect 28684 10140 28690 10152
rect 28858 10149 28870 10152
rect 28904 10149 28916 10183
rect 28858 10143 28916 10149
rect 30282 10140 30288 10192
rect 30340 10180 30346 10192
rect 30469 10183 30527 10189
rect 30469 10180 30481 10183
rect 30340 10152 30481 10180
rect 30340 10140 30346 10152
rect 30469 10149 30481 10152
rect 30515 10149 30527 10183
rect 30469 10143 30527 10149
rect 30558 10140 30564 10192
rect 30616 10180 30622 10192
rect 30616 10152 30709 10180
rect 30616 10140 30622 10152
rect 32214 10140 32220 10192
rect 32272 10180 32278 10192
rect 33060 10189 33088 10220
rect 33873 10217 33885 10220
rect 33919 10217 33931 10251
rect 36262 10248 36268 10260
rect 36223 10220 36268 10248
rect 33873 10211 33931 10217
rect 36262 10208 36268 10220
rect 36320 10208 36326 10260
rect 33045 10183 33103 10189
rect 33045 10180 33057 10183
rect 32272 10152 33057 10180
rect 32272 10140 32278 10152
rect 33045 10149 33057 10152
rect 33091 10149 33103 10183
rect 33045 10143 33103 10149
rect 33134 10140 33140 10192
rect 33192 10180 33198 10192
rect 33686 10180 33692 10192
rect 33192 10152 33237 10180
rect 33647 10152 33692 10180
rect 33192 10140 33198 10152
rect 33686 10140 33692 10152
rect 33744 10140 33750 10192
rect 34698 10180 34704 10192
rect 34659 10152 34704 10180
rect 34698 10140 34704 10152
rect 34756 10140 34762 10192
rect 34882 10140 34888 10192
rect 34940 10180 34946 10192
rect 36538 10180 36544 10192
rect 34940 10152 36544 10180
rect 34940 10140 34946 10152
rect 36538 10140 36544 10152
rect 36596 10180 36602 10192
rect 36633 10183 36691 10189
rect 36633 10180 36645 10183
rect 36596 10152 36645 10180
rect 36596 10140 36602 10152
rect 36633 10149 36645 10152
rect 36679 10149 36691 10183
rect 36633 10143 36691 10149
rect 26145 10115 26203 10121
rect 26145 10081 26157 10115
rect 26191 10112 26203 10115
rect 26234 10112 26240 10124
rect 26191 10084 26240 10112
rect 26191 10081 26203 10084
rect 26145 10075 26203 10081
rect 26234 10072 26240 10084
rect 26292 10072 26298 10124
rect 36078 10112 36084 10124
rect 36039 10084 36084 10112
rect 36078 10072 36084 10084
rect 36136 10072 36142 10124
rect 21039 10016 22968 10044
rect 21039 10013 21051 10016
rect 20993 10007 21051 10013
rect 23014 10004 23020 10056
rect 23072 10044 23078 10056
rect 23201 10047 23259 10053
rect 23201 10044 23213 10047
rect 23072 10016 23213 10044
rect 23072 10004 23078 10016
rect 23201 10013 23213 10016
rect 23247 10013 23259 10047
rect 23474 10044 23480 10056
rect 23435 10016 23480 10044
rect 23201 10007 23259 10013
rect 23474 10004 23480 10016
rect 23532 10004 23538 10056
rect 26326 10004 26332 10056
rect 26384 10044 26390 10056
rect 26605 10047 26663 10053
rect 26605 10044 26617 10047
rect 26384 10016 26617 10044
rect 26384 10004 26390 10016
rect 26605 10013 26617 10016
rect 26651 10013 26663 10047
rect 26605 10007 26663 10013
rect 26881 10047 26939 10053
rect 26881 10013 26893 10047
rect 26927 10013 26939 10047
rect 28534 10044 28540 10056
rect 28495 10016 28540 10044
rect 26881 10007 26939 10013
rect 15436 9948 16252 9976
rect 23492 9976 23520 10004
rect 25774 9976 25780 9988
rect 23492 9948 25780 9976
rect 15436 9936 15442 9948
rect 25774 9936 25780 9948
rect 25832 9976 25838 9988
rect 26896 9976 26924 10007
rect 28534 10004 28540 10016
rect 28592 10004 28598 10056
rect 31110 10044 31116 10056
rect 31023 10016 31116 10044
rect 31110 10004 31116 10016
rect 31168 10044 31174 10056
rect 34606 10044 34612 10056
rect 31168 10016 34284 10044
rect 34567 10016 34612 10044
rect 31168 10004 31174 10016
rect 32309 9979 32367 9985
rect 32309 9976 32321 9979
rect 25832 9948 26924 9976
rect 28092 9948 32321 9976
rect 25832 9936 25838 9948
rect 28092 9920 28120 9948
rect 32309 9945 32321 9948
rect 32355 9976 32367 9979
rect 32490 9976 32496 9988
rect 32355 9948 32496 9976
rect 32355 9945 32367 9948
rect 32309 9939 32367 9945
rect 32490 9936 32496 9948
rect 32548 9936 32554 9988
rect 34256 9976 34284 10016
rect 34606 10004 34612 10016
rect 34664 10004 34670 10056
rect 34885 10047 34943 10053
rect 34885 10013 34897 10047
rect 34931 10013 34943 10047
rect 34885 10007 34943 10013
rect 34900 9976 34928 10007
rect 35250 9976 35256 9988
rect 34256 9948 35256 9976
rect 35250 9936 35256 9948
rect 35308 9936 35314 9988
rect 1670 9908 1676 9920
rect 1631 9880 1676 9908
rect 1670 9868 1676 9880
rect 1728 9868 1734 9920
rect 8711 9911 8769 9917
rect 8711 9877 8723 9911
rect 8757 9908 8769 9911
rect 8846 9908 8852 9920
rect 8757 9880 8852 9908
rect 8757 9877 8769 9880
rect 8711 9871 8769 9877
rect 8846 9868 8852 9880
rect 8904 9868 8910 9920
rect 9030 9908 9036 9920
rect 8991 9880 9036 9908
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 9953 9911 10011 9917
rect 9953 9877 9965 9911
rect 9999 9908 10011 9911
rect 10042 9908 10048 9920
rect 9999 9880 10048 9908
rect 9999 9877 10011 9880
rect 9953 9871 10011 9877
rect 10042 9868 10048 9880
rect 10100 9908 10106 9920
rect 16114 9908 16120 9920
rect 10100 9880 16120 9908
rect 10100 9868 10106 9880
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 23658 9868 23664 9920
rect 23716 9908 23722 9920
rect 24121 9911 24179 9917
rect 24121 9908 24133 9911
rect 23716 9880 24133 9908
rect 23716 9868 23722 9880
rect 24121 9877 24133 9880
rect 24167 9877 24179 9911
rect 24121 9871 24179 9877
rect 24394 9868 24400 9920
rect 24452 9908 24458 9920
rect 25958 9908 25964 9920
rect 24452 9880 25964 9908
rect 24452 9868 24458 9880
rect 25958 9868 25964 9880
rect 26016 9868 26022 9920
rect 27062 9868 27068 9920
rect 27120 9908 27126 9920
rect 27801 9911 27859 9917
rect 27801 9908 27813 9911
rect 27120 9880 27813 9908
rect 27120 9868 27126 9880
rect 27801 9877 27813 9880
rect 27847 9908 27859 9911
rect 28074 9908 28080 9920
rect 27847 9880 28080 9908
rect 27847 9877 27859 9880
rect 27801 9871 27859 9877
rect 28074 9868 28080 9880
rect 28132 9868 28138 9920
rect 30098 9908 30104 9920
rect 30059 9880 30104 9908
rect 30098 9868 30104 9880
rect 30156 9868 30162 9920
rect 33873 9911 33931 9917
rect 33873 9877 33885 9911
rect 33919 9908 33931 9911
rect 34057 9911 34115 9917
rect 34057 9908 34069 9911
rect 33919 9880 34069 9908
rect 33919 9877 33931 9880
rect 33873 9871 33931 9877
rect 34057 9877 34069 9880
rect 34103 9908 34115 9911
rect 35618 9908 35624 9920
rect 34103 9880 35624 9908
rect 34103 9877 34115 9880
rect 34057 9871 34115 9877
rect 35618 9868 35624 9880
rect 35676 9868 35682 9920
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 2041 9707 2099 9713
rect 2041 9673 2053 9707
rect 2087 9704 2099 9707
rect 2406 9704 2412 9716
rect 2087 9676 2412 9704
rect 2087 9673 2099 9676
rect 2041 9667 2099 9673
rect 2406 9664 2412 9676
rect 2464 9704 2470 9716
rect 3973 9707 4031 9713
rect 3973 9704 3985 9707
rect 2464 9676 3985 9704
rect 2464 9664 2470 9676
rect 3973 9673 3985 9676
rect 4019 9673 4031 9707
rect 5166 9704 5172 9716
rect 5127 9676 5172 9704
rect 3973 9667 4031 9673
rect 3988 9636 4016 9667
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 5902 9664 5908 9716
rect 5960 9704 5966 9716
rect 5997 9707 6055 9713
rect 5997 9704 6009 9707
rect 5960 9676 6009 9704
rect 5960 9664 5966 9676
rect 5997 9673 6009 9676
rect 6043 9673 6055 9707
rect 5997 9667 6055 9673
rect 8846 9664 8852 9716
rect 8904 9704 8910 9716
rect 9585 9707 9643 9713
rect 9585 9704 9597 9707
rect 8904 9676 9597 9704
rect 8904 9664 8910 9676
rect 9585 9673 9597 9676
rect 9631 9704 9643 9707
rect 10502 9704 10508 9716
rect 9631 9676 10508 9704
rect 9631 9673 9643 9676
rect 9585 9667 9643 9673
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 11422 9704 11428 9716
rect 11383 9676 11428 9704
rect 11422 9664 11428 9676
rect 11480 9664 11486 9716
rect 11606 9664 11612 9716
rect 11664 9704 11670 9716
rect 11793 9707 11851 9713
rect 11793 9704 11805 9707
rect 11664 9676 11805 9704
rect 11664 9664 11670 9676
rect 11793 9673 11805 9676
rect 11839 9673 11851 9707
rect 11793 9667 11851 9673
rect 16022 9664 16028 9716
rect 16080 9704 16086 9716
rect 16577 9707 16635 9713
rect 16577 9704 16589 9707
rect 16080 9676 16589 9704
rect 16080 9664 16086 9676
rect 16577 9673 16589 9676
rect 16623 9704 16635 9707
rect 16666 9704 16672 9716
rect 16623 9676 16672 9704
rect 16623 9673 16635 9676
rect 16577 9667 16635 9673
rect 16666 9664 16672 9676
rect 16724 9664 16730 9716
rect 17865 9707 17923 9713
rect 17865 9673 17877 9707
rect 17911 9704 17923 9707
rect 18138 9704 18144 9716
rect 17911 9676 18144 9704
rect 17911 9673 17923 9676
rect 17865 9667 17923 9673
rect 18138 9664 18144 9676
rect 18196 9664 18202 9716
rect 18782 9704 18788 9716
rect 18743 9676 18788 9704
rect 18782 9664 18788 9676
rect 18840 9664 18846 9716
rect 20162 9704 20168 9716
rect 20123 9676 20168 9704
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 21910 9704 21916 9716
rect 21871 9676 21916 9704
rect 21910 9664 21916 9676
rect 21968 9704 21974 9716
rect 22189 9707 22247 9713
rect 22189 9704 22201 9707
rect 21968 9676 22201 9704
rect 21968 9664 21974 9676
rect 22189 9673 22201 9676
rect 22235 9673 22247 9707
rect 22189 9667 22247 9673
rect 22741 9707 22799 9713
rect 22741 9673 22753 9707
rect 22787 9704 22799 9707
rect 23014 9704 23020 9716
rect 22787 9676 23020 9704
rect 22787 9673 22799 9676
rect 22741 9667 22799 9673
rect 23014 9664 23020 9676
rect 23072 9664 23078 9716
rect 23109 9707 23167 9713
rect 23109 9673 23121 9707
rect 23155 9704 23167 9707
rect 23198 9704 23204 9716
rect 23155 9676 23204 9704
rect 23155 9673 23167 9676
rect 23109 9667 23167 9673
rect 23198 9664 23204 9676
rect 23256 9664 23262 9716
rect 24578 9704 24584 9716
rect 24539 9676 24584 9704
rect 24578 9664 24584 9676
rect 24636 9664 24642 9716
rect 24854 9704 24860 9716
rect 24815 9676 24860 9704
rect 24854 9664 24860 9676
rect 24912 9704 24918 9716
rect 25225 9707 25283 9713
rect 25225 9704 25237 9707
rect 24912 9676 25237 9704
rect 24912 9664 24918 9676
rect 25225 9673 25237 9676
rect 25271 9673 25283 9707
rect 25225 9667 25283 9673
rect 25958 9664 25964 9716
rect 26016 9704 26022 9716
rect 26513 9707 26571 9713
rect 26513 9704 26525 9707
rect 26016 9676 26525 9704
rect 26016 9664 26022 9676
rect 26513 9673 26525 9676
rect 26559 9673 26571 9707
rect 26513 9667 26571 9673
rect 30282 9664 30288 9716
rect 30340 9704 30346 9716
rect 30837 9707 30895 9713
rect 30837 9704 30849 9707
rect 30340 9676 30849 9704
rect 30340 9664 30346 9676
rect 30837 9673 30849 9676
rect 30883 9673 30895 9707
rect 30837 9667 30895 9673
rect 31435 9707 31493 9713
rect 31435 9673 31447 9707
rect 31481 9704 31493 9707
rect 32306 9704 32312 9716
rect 31481 9676 32312 9704
rect 31481 9673 31493 9676
rect 31435 9667 31493 9673
rect 32306 9664 32312 9676
rect 32364 9664 32370 9716
rect 33134 9664 33140 9716
rect 33192 9704 33198 9716
rect 33229 9707 33287 9713
rect 33229 9704 33241 9707
rect 33192 9676 33241 9704
rect 33192 9664 33198 9676
rect 33229 9673 33241 9676
rect 33275 9704 33287 9707
rect 33505 9707 33563 9713
rect 33505 9704 33517 9707
rect 33275 9676 33517 9704
rect 33275 9673 33287 9676
rect 33229 9667 33287 9673
rect 33505 9673 33517 9676
rect 33551 9673 33563 9707
rect 33505 9667 33563 9673
rect 33965 9707 34023 9713
rect 33965 9673 33977 9707
rect 34011 9704 34023 9707
rect 34606 9704 34612 9716
rect 34011 9676 34612 9704
rect 34011 9673 34023 9676
rect 33965 9667 34023 9673
rect 34606 9664 34612 9676
rect 34664 9664 34670 9716
rect 6641 9639 6699 9645
rect 3988 9608 4154 9636
rect 2314 9568 2320 9580
rect 2275 9540 2320 9568
rect 2314 9528 2320 9540
rect 2372 9568 2378 9580
rect 3237 9571 3295 9577
rect 3237 9568 3249 9571
rect 2372 9540 3249 9568
rect 2372 9528 2378 9540
rect 3237 9537 3249 9540
rect 3283 9537 3295 9571
rect 4126 9568 4154 9608
rect 6641 9605 6653 9639
rect 6687 9636 6699 9639
rect 7374 9636 7380 9648
rect 6687 9608 7380 9636
rect 6687 9605 6699 9608
rect 6641 9599 6699 9605
rect 7374 9596 7380 9608
rect 7432 9596 7438 9648
rect 9217 9639 9275 9645
rect 9217 9605 9229 9639
rect 9263 9636 9275 9639
rect 12342 9636 12348 9648
rect 9263 9608 12348 9636
rect 9263 9605 9275 9608
rect 9217 9599 9275 9605
rect 12342 9596 12348 9608
rect 12400 9636 12406 9648
rect 13725 9639 13783 9645
rect 12400 9608 12848 9636
rect 12400 9596 12406 9608
rect 8478 9568 8484 9580
rect 4126 9540 8484 9568
rect 3237 9531 3295 9537
rect 4632 9509 4660 9540
rect 8478 9528 8484 9540
rect 8536 9528 8542 9580
rect 8665 9571 8723 9577
rect 8665 9537 8677 9571
rect 8711 9568 8723 9571
rect 9030 9568 9036 9580
rect 8711 9540 9036 9568
rect 8711 9537 8723 9540
rect 8665 9531 8723 9537
rect 9030 9528 9036 9540
rect 9088 9528 9094 9580
rect 10134 9568 10140 9580
rect 10095 9540 10140 9568
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 10962 9528 10968 9580
rect 11020 9568 11026 9580
rect 12250 9568 12256 9580
rect 11020 9540 12256 9568
rect 11020 9528 11026 9540
rect 12250 9528 12256 9540
rect 12308 9568 12314 9580
rect 12820 9577 12848 9608
rect 13725 9605 13737 9639
rect 13771 9636 13783 9639
rect 14182 9636 14188 9648
rect 13771 9608 14188 9636
rect 13771 9605 13783 9608
rect 13725 9599 13783 9605
rect 14182 9596 14188 9608
rect 14240 9596 14246 9648
rect 15930 9596 15936 9648
rect 15988 9636 15994 9648
rect 16209 9639 16267 9645
rect 16209 9636 16221 9639
rect 15988 9608 16221 9636
rect 15988 9596 15994 9608
rect 16209 9605 16221 9608
rect 16255 9605 16267 9639
rect 16209 9599 16267 9605
rect 23290 9596 23296 9648
rect 23348 9636 23354 9648
rect 26326 9636 26332 9648
rect 23348 9608 26332 9636
rect 23348 9596 23354 9608
rect 26326 9596 26332 9608
rect 26384 9596 26390 9648
rect 27062 9636 27068 9648
rect 27023 9608 27068 9636
rect 27062 9596 27068 9608
rect 27120 9596 27126 9648
rect 30193 9639 30251 9645
rect 30193 9605 30205 9639
rect 30239 9636 30251 9639
rect 30558 9636 30564 9648
rect 30239 9608 30564 9636
rect 30239 9605 30251 9608
rect 30193 9599 30251 9605
rect 30558 9596 30564 9608
rect 30616 9596 30622 9648
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 12308 9540 12541 9568
rect 12308 9528 12314 9540
rect 12529 9537 12541 9540
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 12805 9571 12863 9577
rect 12805 9537 12817 9571
rect 12851 9537 12863 9571
rect 12805 9531 12863 9537
rect 13630 9528 13636 9580
rect 13688 9568 13694 9580
rect 15010 9568 15016 9580
rect 13688 9540 15016 9568
rect 13688 9528 13694 9540
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 19150 9528 19156 9580
rect 19208 9568 19214 9580
rect 19245 9571 19303 9577
rect 19245 9568 19257 9571
rect 19208 9540 19257 9568
rect 19208 9528 19214 9540
rect 19245 9537 19257 9540
rect 19291 9537 19303 9571
rect 19245 9531 19303 9537
rect 19886 9528 19892 9580
rect 19944 9568 19950 9580
rect 20993 9571 21051 9577
rect 20993 9568 21005 9571
rect 19944 9540 21005 9568
rect 19944 9528 19950 9540
rect 20993 9537 21005 9540
rect 21039 9568 21051 9571
rect 21818 9568 21824 9580
rect 21039 9540 21824 9568
rect 21039 9537 21051 9540
rect 20993 9531 21051 9537
rect 21818 9528 21824 9540
rect 21876 9528 21882 9580
rect 23658 9568 23664 9580
rect 23446 9540 23664 9568
rect 3697 9503 3755 9509
rect 3697 9469 3709 9503
rect 3743 9500 3755 9503
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 3743 9472 4445 9500
rect 3743 9469 3755 9472
rect 3697 9463 3755 9469
rect 4433 9469 4445 9472
rect 4479 9469 4491 9503
rect 4433 9463 4491 9469
rect 4617 9503 4675 9509
rect 4617 9469 4629 9503
rect 4663 9469 4675 9503
rect 4617 9463 4675 9469
rect 5629 9503 5687 9509
rect 5629 9469 5641 9503
rect 5675 9500 5687 9503
rect 5756 9503 5814 9509
rect 5756 9500 5768 9503
rect 5675 9472 5768 9500
rect 5675 9469 5687 9472
rect 5629 9463 5687 9469
rect 5756 9469 5768 9472
rect 5802 9500 5814 9503
rect 5902 9500 5908 9512
rect 5802 9472 5908 9500
rect 5802 9469 5814 9472
rect 5756 9463 5814 9469
rect 2406 9392 2412 9444
rect 2464 9432 2470 9444
rect 2961 9435 3019 9441
rect 2464 9404 2509 9432
rect 2464 9392 2470 9404
rect 2961 9401 2973 9435
rect 3007 9432 3019 9435
rect 3050 9432 3056 9444
rect 3007 9404 3056 9432
rect 3007 9401 3019 9404
rect 2961 9395 3019 9401
rect 3050 9392 3056 9404
rect 3108 9392 3114 9444
rect 4448 9432 4476 9463
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 5994 9460 6000 9512
rect 6052 9500 6058 9512
rect 6273 9503 6331 9509
rect 6273 9500 6285 9503
rect 6052 9472 6285 9500
rect 6052 9460 6058 9472
rect 6273 9469 6285 9472
rect 6319 9500 6331 9503
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 6319 9472 6837 9500
rect 6319 9469 6331 9472
rect 6273 9463 6331 9469
rect 6825 9469 6837 9472
rect 6871 9469 6883 9503
rect 7374 9500 7380 9512
rect 7335 9472 7380 9500
rect 6825 9463 6883 9469
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 10318 9460 10324 9512
rect 10376 9500 10382 9512
rect 11057 9503 11115 9509
rect 11057 9500 11069 9503
rect 10376 9472 11069 9500
rect 10376 9460 10382 9472
rect 11057 9469 11069 9472
rect 11103 9500 11115 9503
rect 12161 9503 12219 9509
rect 12161 9500 12173 9503
rect 11103 9472 12173 9500
rect 11103 9469 11115 9472
rect 11057 9463 11115 9469
rect 12161 9469 12173 9472
rect 12207 9469 12219 9503
rect 12161 9463 12219 9469
rect 7190 9432 7196 9444
rect 4448 9404 7196 9432
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 7466 9392 7472 9444
rect 7524 9432 7530 9444
rect 8386 9432 8392 9444
rect 7524 9404 8392 9432
rect 7524 9392 7530 9404
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 8754 9432 8760 9444
rect 8715 9404 8760 9432
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 10458 9435 10516 9441
rect 10458 9432 10470 9435
rect 9968 9404 10470 9432
rect 1486 9324 1492 9376
rect 1544 9364 1550 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 1544 9336 1593 9364
rect 1544 9324 1550 9336
rect 1581 9333 1593 9336
rect 1627 9333 1639 9367
rect 1581 9327 1639 9333
rect 4062 9324 4068 9376
rect 4120 9364 4126 9376
rect 4249 9367 4307 9373
rect 4249 9364 4261 9367
rect 4120 9336 4261 9364
rect 4120 9324 4126 9336
rect 4249 9333 4261 9336
rect 4295 9333 4307 9367
rect 4249 9327 4307 9333
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 6917 9367 6975 9373
rect 6917 9364 6929 9367
rect 6788 9336 6929 9364
rect 6788 9324 6794 9336
rect 6917 9333 6929 9336
rect 6963 9333 6975 9367
rect 7834 9364 7840 9376
rect 7795 9336 7840 9364
rect 6917 9327 6975 9333
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 9766 9324 9772 9376
rect 9824 9364 9830 9376
rect 9968 9373 9996 9404
rect 10458 9401 10470 9404
rect 10504 9401 10516 9435
rect 10458 9395 10516 9401
rect 9953 9367 10011 9373
rect 9953 9364 9965 9367
rect 9824 9336 9965 9364
rect 9824 9324 9830 9336
rect 9953 9333 9965 9336
rect 9999 9333 10011 9367
rect 12176 9364 12204 9463
rect 13538 9460 13544 9512
rect 13596 9500 13602 9512
rect 14068 9503 14126 9509
rect 14068 9500 14080 9503
rect 13596 9472 14080 9500
rect 13596 9460 13602 9472
rect 14068 9469 14080 9472
rect 14114 9500 14126 9503
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 14114 9472 14473 9500
rect 14114 9469 14126 9472
rect 14068 9463 14126 9469
rect 14461 9469 14473 9472
rect 14507 9469 14519 9503
rect 14461 9463 14519 9469
rect 15194 9460 15200 9512
rect 15252 9500 15258 9512
rect 15933 9503 15991 9509
rect 15933 9500 15945 9503
rect 15252 9472 15945 9500
rect 15252 9460 15258 9472
rect 15933 9469 15945 9472
rect 15979 9469 15991 9503
rect 15933 9463 15991 9469
rect 17012 9503 17070 9509
rect 17012 9469 17024 9503
rect 17058 9500 17070 9503
rect 17494 9500 17500 9512
rect 17058 9472 17500 9500
rect 17058 9469 17070 9472
rect 17012 9463 17070 9469
rect 17494 9460 17500 9472
rect 17552 9460 17558 9512
rect 18300 9503 18358 9509
rect 18300 9469 18312 9503
rect 18346 9500 18358 9503
rect 18782 9500 18788 9512
rect 18346 9472 18788 9500
rect 18346 9469 18358 9472
rect 18300 9463 18358 9469
rect 18782 9460 18788 9472
rect 18840 9460 18846 9512
rect 23014 9460 23020 9512
rect 23072 9500 23078 9512
rect 23446 9500 23474 9540
rect 23658 9528 23664 9540
rect 23716 9528 23722 9580
rect 24670 9528 24676 9580
rect 24728 9568 24734 9580
rect 25498 9568 25504 9580
rect 24728 9540 25504 9568
rect 24728 9528 24734 9540
rect 25498 9528 25504 9540
rect 25556 9528 25562 9580
rect 25774 9568 25780 9580
rect 25735 9540 25780 9568
rect 25774 9528 25780 9540
rect 25832 9528 25838 9580
rect 28353 9571 28411 9577
rect 28353 9537 28365 9571
rect 28399 9568 28411 9571
rect 28534 9568 28540 9580
rect 28399 9540 28540 9568
rect 28399 9537 28411 9540
rect 28353 9531 28411 9537
rect 28534 9528 28540 9540
rect 28592 9528 28598 9580
rect 29273 9571 29331 9577
rect 29273 9537 29285 9571
rect 29319 9568 29331 9571
rect 29638 9568 29644 9580
rect 29319 9540 29644 9568
rect 29319 9537 29331 9540
rect 29273 9531 29331 9537
rect 29638 9528 29644 9540
rect 29696 9528 29702 9580
rect 32309 9571 32367 9577
rect 32309 9537 32321 9571
rect 32355 9568 32367 9571
rect 32674 9568 32680 9580
rect 32355 9540 32680 9568
rect 32355 9537 32367 9540
rect 32309 9531 32367 9537
rect 32674 9528 32680 9540
rect 32732 9528 32738 9580
rect 34790 9528 34796 9580
rect 34848 9568 34854 9580
rect 34977 9571 35035 9577
rect 34977 9568 34989 9571
rect 34848 9540 34989 9568
rect 34848 9528 34854 9540
rect 34977 9537 34989 9540
rect 35023 9537 35035 9571
rect 35250 9568 35256 9580
rect 35211 9540 35256 9568
rect 34977 9531 35035 9537
rect 35250 9528 35256 9540
rect 35308 9528 35314 9580
rect 35618 9528 35624 9580
rect 35676 9568 35682 9580
rect 36817 9571 36875 9577
rect 36817 9568 36829 9571
rect 35676 9540 36829 9568
rect 35676 9528 35682 9540
rect 36817 9537 36829 9540
rect 36863 9537 36875 9571
rect 36817 9531 36875 9537
rect 23072 9472 23474 9500
rect 27893 9503 27951 9509
rect 23072 9460 23078 9472
rect 27893 9469 27905 9503
rect 27939 9469 27951 9503
rect 28074 9500 28080 9512
rect 28035 9472 28080 9500
rect 27893 9463 27951 9469
rect 12621 9435 12679 9441
rect 12621 9401 12633 9435
rect 12667 9401 12679 9435
rect 12621 9395 12679 9401
rect 14921 9435 14979 9441
rect 14921 9401 14933 9435
rect 14967 9432 14979 9435
rect 15375 9435 15433 9441
rect 15375 9432 15387 9435
rect 14967 9404 15387 9432
rect 14967 9401 14979 9404
rect 14921 9395 14979 9401
rect 15375 9401 15387 9404
rect 15421 9432 15433 9435
rect 15838 9432 15844 9444
rect 15421 9404 15844 9432
rect 15421 9401 15433 9404
rect 15375 9395 15433 9401
rect 12636 9364 12664 9395
rect 15838 9392 15844 9404
rect 15896 9392 15902 9444
rect 21358 9441 21364 9444
rect 19153 9435 19211 9441
rect 19153 9401 19165 9435
rect 19199 9432 19211 9435
rect 19607 9435 19665 9441
rect 19607 9432 19619 9435
rect 19199 9404 19619 9432
rect 19199 9401 19211 9404
rect 19153 9395 19211 9401
rect 19607 9401 19619 9404
rect 19653 9432 19665 9435
rect 20901 9435 20959 9441
rect 20901 9432 20913 9435
rect 19653 9404 20913 9432
rect 19653 9401 19665 9404
rect 19607 9395 19665 9401
rect 20901 9401 20913 9404
rect 20947 9432 20959 9435
rect 21355 9432 21364 9441
rect 20947 9404 21364 9432
rect 20947 9401 20959 9404
rect 20901 9395 20959 9401
rect 21355 9395 21364 9404
rect 21358 9392 21364 9395
rect 21416 9392 21422 9444
rect 23477 9435 23535 9441
rect 23477 9401 23489 9435
rect 23523 9432 23535 9435
rect 23658 9432 23664 9444
rect 23523 9404 23664 9432
rect 23523 9401 23535 9404
rect 23477 9395 23535 9401
rect 23658 9392 23664 9404
rect 23716 9432 23722 9444
rect 23982 9435 24040 9441
rect 23982 9432 23994 9435
rect 23716 9404 23994 9432
rect 23716 9392 23722 9404
rect 23982 9401 23994 9404
rect 24028 9401 24040 9435
rect 23982 9395 24040 9401
rect 25593 9435 25651 9441
rect 25593 9401 25605 9435
rect 25639 9401 25651 9435
rect 25593 9395 25651 9401
rect 27525 9435 27583 9441
rect 27525 9401 27537 9435
rect 27571 9432 27583 9435
rect 27908 9432 27936 9463
rect 28074 9460 28080 9472
rect 28132 9460 28138 9512
rect 31364 9503 31422 9509
rect 31364 9469 31376 9503
rect 31410 9500 31422 9503
rect 31754 9500 31760 9512
rect 31410 9472 31760 9500
rect 31410 9469 31422 9472
rect 31364 9463 31422 9469
rect 28258 9432 28264 9444
rect 27571 9404 28264 9432
rect 27571 9401 27583 9404
rect 27525 9395 27583 9401
rect 12176 9336 12664 9364
rect 9953 9327 10011 9333
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14139 9367 14197 9373
rect 14139 9364 14151 9367
rect 13964 9336 14151 9364
rect 13964 9324 13970 9336
rect 14139 9333 14151 9336
rect 14185 9333 14197 9367
rect 14139 9327 14197 9333
rect 17083 9367 17141 9373
rect 17083 9333 17095 9367
rect 17129 9364 17141 9367
rect 17310 9364 17316 9376
rect 17129 9336 17316 9364
rect 17129 9333 17141 9336
rect 17083 9327 17141 9333
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 17494 9364 17500 9376
rect 17455 9336 17500 9364
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 18371 9367 18429 9373
rect 18371 9333 18383 9367
rect 18417 9364 18429 9367
rect 18598 9364 18604 9376
rect 18417 9336 18604 9364
rect 18417 9333 18429 9336
rect 18371 9327 18429 9333
rect 18598 9324 18604 9336
rect 18656 9324 18662 9376
rect 19518 9324 19524 9376
rect 19576 9364 19582 9376
rect 20533 9367 20591 9373
rect 20533 9364 20545 9367
rect 19576 9336 20545 9364
rect 19576 9324 19582 9336
rect 20533 9333 20545 9336
rect 20579 9364 20591 9367
rect 21726 9364 21732 9376
rect 20579 9336 21732 9364
rect 20579 9333 20591 9336
rect 20533 9327 20591 9333
rect 21726 9324 21732 9336
rect 21784 9324 21790 9376
rect 24854 9324 24860 9376
rect 24912 9364 24918 9376
rect 25608 9364 25636 9395
rect 28258 9392 28264 9404
rect 28316 9392 28322 9444
rect 29594 9435 29652 9441
rect 29594 9432 29606 9435
rect 29012 9404 29606 9432
rect 24912 9336 25636 9364
rect 24912 9324 24918 9336
rect 28626 9324 28632 9376
rect 28684 9364 28690 9376
rect 28721 9367 28779 9373
rect 28721 9364 28733 9367
rect 28684 9336 28733 9364
rect 28684 9324 28690 9336
rect 28721 9333 28733 9336
rect 28767 9364 28779 9367
rect 28810 9364 28816 9376
rect 28767 9336 28816 9364
rect 28767 9333 28779 9336
rect 28721 9327 28779 9333
rect 28810 9324 28816 9336
rect 28868 9364 28874 9376
rect 29012 9373 29040 9404
rect 29594 9401 29606 9404
rect 29640 9401 29652 9435
rect 29594 9395 29652 9401
rect 30742 9392 30748 9444
rect 30800 9432 30806 9444
rect 31379 9432 31407 9463
rect 31754 9460 31760 9472
rect 31812 9460 31818 9512
rect 32630 9435 32688 9441
rect 32630 9432 32642 9435
rect 30800 9404 31407 9432
rect 32140 9404 32642 9432
rect 30800 9392 30806 9404
rect 28997 9367 29055 9373
rect 28997 9364 29009 9367
rect 28868 9336 29009 9364
rect 28868 9324 28874 9336
rect 28997 9333 29009 9336
rect 29043 9333 29055 9367
rect 28997 9327 29055 9333
rect 32030 9324 32036 9376
rect 32088 9364 32094 9376
rect 32140 9373 32168 9404
rect 32630 9401 32642 9404
rect 32676 9401 32688 9435
rect 32630 9395 32688 9401
rect 34701 9435 34759 9441
rect 34701 9401 34713 9435
rect 34747 9432 34759 9435
rect 35066 9432 35072 9444
rect 34747 9404 35072 9432
rect 34747 9401 34759 9404
rect 34701 9395 34759 9401
rect 35066 9392 35072 9404
rect 35124 9432 35130 9444
rect 36354 9432 36360 9444
rect 35124 9404 36360 9432
rect 35124 9392 35130 9404
rect 36354 9392 36360 9404
rect 36412 9392 36418 9444
rect 36538 9432 36544 9444
rect 36499 9404 36544 9432
rect 36538 9392 36544 9404
rect 36596 9392 36602 9444
rect 36630 9392 36636 9444
rect 36688 9432 36694 9444
rect 36688 9404 36733 9432
rect 36688 9392 36694 9404
rect 32125 9367 32183 9373
rect 32125 9364 32137 9367
rect 32088 9336 32137 9364
rect 32088 9324 32094 9336
rect 32125 9333 32137 9336
rect 32171 9333 32183 9367
rect 34330 9364 34336 9376
rect 34291 9336 34336 9364
rect 32125 9327 32183 9333
rect 34330 9324 34336 9336
rect 34388 9324 34394 9376
rect 36078 9364 36084 9376
rect 36039 9336 36084 9364
rect 36078 9324 36084 9336
rect 36136 9324 36142 9376
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 1728 9132 6868 9160
rect 1728 9120 1734 9132
rect 2590 9092 2596 9104
rect 2551 9064 2596 9092
rect 2590 9052 2596 9064
rect 2648 9052 2654 9104
rect 5074 9092 5080 9104
rect 5035 9064 5080 9092
rect 5074 9052 5080 9064
rect 5132 9052 5138 9104
rect 6546 9092 6552 9104
rect 6507 9064 6552 9092
rect 6546 9052 6552 9064
rect 6604 9052 6610 9104
rect 6638 9052 6644 9104
rect 6696 9092 6702 9104
rect 6840 9092 6868 9132
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 7561 9163 7619 9169
rect 7561 9160 7573 9163
rect 6972 9132 7573 9160
rect 6972 9120 6978 9132
rect 7561 9129 7573 9132
rect 7607 9160 7619 9163
rect 8113 9163 8171 9169
rect 8113 9160 8125 9163
rect 7607 9132 8125 9160
rect 7607 9129 7619 9132
rect 7561 9123 7619 9129
rect 8113 9129 8125 9132
rect 8159 9129 8171 9163
rect 10134 9160 10140 9172
rect 10095 9132 10140 9160
rect 8113 9123 8171 9129
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 10778 9120 10784 9172
rect 10836 9160 10842 9172
rect 10873 9163 10931 9169
rect 10873 9160 10885 9163
rect 10836 9132 10885 9160
rect 10836 9120 10842 9132
rect 10873 9129 10885 9132
rect 10919 9129 10931 9163
rect 11422 9160 11428 9172
rect 11383 9132 11428 9160
rect 10873 9123 10931 9129
rect 11422 9120 11428 9132
rect 11480 9120 11486 9172
rect 11606 9120 11612 9172
rect 11664 9160 11670 9172
rect 11977 9163 12035 9169
rect 11977 9160 11989 9163
rect 11664 9132 11989 9160
rect 11664 9120 11670 9132
rect 11977 9129 11989 9132
rect 12023 9129 12035 9163
rect 11977 9123 12035 9129
rect 12250 9120 12256 9172
rect 12308 9160 12314 9172
rect 12437 9163 12495 9169
rect 12437 9160 12449 9163
rect 12308 9132 12449 9160
rect 12308 9120 12314 9132
rect 12437 9129 12449 9132
rect 12483 9129 12495 9163
rect 15010 9160 15016 9172
rect 14971 9132 15016 9160
rect 12437 9123 12495 9129
rect 15010 9120 15016 9132
rect 15068 9120 15074 9172
rect 16666 9160 16672 9172
rect 16627 9132 16672 9160
rect 16666 9120 16672 9132
rect 16724 9120 16730 9172
rect 17678 9160 17684 9172
rect 17639 9132 17684 9160
rect 17678 9120 17684 9132
rect 17736 9120 17742 9172
rect 18598 9120 18604 9172
rect 18656 9160 18662 9172
rect 18693 9163 18751 9169
rect 18693 9160 18705 9163
rect 18656 9132 18705 9160
rect 18656 9120 18662 9132
rect 18693 9129 18705 9132
rect 18739 9160 18751 9163
rect 20714 9160 20720 9172
rect 18739 9132 19012 9160
rect 20675 9132 20720 9160
rect 18739 9129 18751 9132
rect 18693 9123 18751 9129
rect 9815 9095 9873 9101
rect 6696 9064 6741 9092
rect 6840 9064 8610 9092
rect 6696 9052 6702 9064
rect 1464 9027 1522 9033
rect 1464 8993 1476 9027
rect 1510 9024 1522 9027
rect 1670 9024 1676 9036
rect 1510 8996 1676 9024
rect 1510 8993 1522 8996
rect 1464 8987 1522 8993
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 8110 9024 8116 9036
rect 8071 8996 8116 9024
rect 8110 8984 8116 8996
rect 8168 8984 8174 9036
rect 8478 9024 8484 9036
rect 8439 8996 8484 9024
rect 8478 8984 8484 8996
rect 8536 8984 8542 9036
rect 8582 9024 8610 9064
rect 9815 9061 9827 9095
rect 9861 9092 9873 9095
rect 10226 9092 10232 9104
rect 9861 9064 10232 9092
rect 9861 9061 9873 9064
rect 9815 9055 9873 9061
rect 10226 9052 10232 9064
rect 10284 9052 10290 9104
rect 13814 9052 13820 9104
rect 13872 9092 13878 9104
rect 14369 9095 14427 9101
rect 13872 9064 13917 9092
rect 13872 9052 13878 9064
rect 14369 9061 14381 9095
rect 14415 9092 14427 9095
rect 15378 9092 15384 9104
rect 14415 9064 15384 9092
rect 14415 9061 14427 9064
rect 14369 9055 14427 9061
rect 15378 9052 15384 9064
rect 15436 9052 15442 9104
rect 15838 9052 15844 9104
rect 15896 9092 15902 9104
rect 18984 9101 19012 9132
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 21818 9160 21824 9172
rect 21779 9132 21824 9160
rect 21818 9120 21824 9132
rect 21876 9120 21882 9172
rect 24762 9120 24768 9172
rect 24820 9160 24826 9172
rect 25041 9163 25099 9169
rect 25041 9160 25053 9163
rect 24820 9132 25053 9160
rect 24820 9120 24826 9132
rect 25041 9129 25053 9132
rect 25087 9129 25099 9163
rect 25041 9123 25099 9129
rect 25130 9120 25136 9172
rect 25188 9160 25194 9172
rect 26605 9163 26663 9169
rect 26605 9160 26617 9163
rect 25188 9132 26617 9160
rect 25188 9120 25194 9132
rect 26605 9129 26617 9132
rect 26651 9129 26663 9163
rect 28534 9160 28540 9172
rect 28495 9132 28540 9160
rect 26605 9123 26663 9129
rect 28534 9120 28540 9132
rect 28592 9120 28598 9172
rect 29549 9163 29607 9169
rect 29549 9129 29561 9163
rect 29595 9160 29607 9163
rect 30098 9160 30104 9172
rect 29595 9132 30104 9160
rect 29595 9129 29607 9132
rect 29549 9123 29607 9129
rect 30098 9120 30104 9132
rect 30156 9120 30162 9172
rect 34054 9160 34060 9172
rect 34015 9132 34060 9160
rect 34054 9120 34060 9132
rect 34112 9120 34118 9172
rect 34790 9120 34796 9172
rect 34848 9160 34854 9172
rect 35253 9163 35311 9169
rect 35253 9160 35265 9163
rect 34848 9132 35265 9160
rect 34848 9120 34854 9132
rect 35253 9129 35265 9132
rect 35299 9129 35311 9163
rect 35802 9160 35808 9172
rect 35763 9132 35808 9160
rect 35253 9123 35311 9129
rect 35802 9120 35808 9132
rect 35860 9120 35866 9172
rect 36354 9160 36360 9172
rect 36315 9132 36360 9160
rect 36354 9120 36360 9132
rect 36412 9120 36418 9172
rect 36630 9160 36636 9172
rect 36591 9132 36636 9160
rect 36630 9120 36636 9132
rect 36688 9120 36694 9172
rect 16070 9095 16128 9101
rect 16070 9092 16082 9095
rect 15896 9064 16082 9092
rect 15896 9052 15902 9064
rect 16070 9061 16082 9064
rect 16116 9061 16128 9095
rect 16070 9055 16128 9061
rect 18969 9095 19027 9101
rect 18969 9061 18981 9095
rect 19015 9061 19027 9095
rect 18969 9055 19027 9061
rect 19058 9052 19064 9104
rect 19116 9092 19122 9104
rect 19116 9064 19161 9092
rect 19116 9052 19122 9064
rect 19702 9052 19708 9104
rect 19760 9092 19766 9104
rect 19981 9095 20039 9101
rect 19981 9092 19993 9095
rect 19760 9064 19993 9092
rect 19760 9052 19766 9064
rect 19981 9061 19993 9064
rect 20027 9092 20039 9095
rect 23014 9092 23020 9104
rect 20027 9064 22876 9092
rect 22975 9064 23020 9092
rect 20027 9061 20039 9064
rect 19981 9055 20039 9061
rect 9728 9027 9786 9033
rect 9728 9024 9740 9027
rect 8582 8996 9740 9024
rect 9728 8993 9740 8996
rect 9774 9024 9786 9027
rect 9950 9024 9956 9036
rect 9774 8996 9956 9024
rect 9774 8993 9786 8996
rect 9728 8987 9786 8993
rect 9950 8984 9956 8996
rect 10008 9024 10014 9036
rect 11698 9024 11704 9036
rect 10008 8996 11704 9024
rect 10008 8984 10014 8996
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 15746 9024 15752 9036
rect 15707 8996 15752 9024
rect 15746 8984 15752 8996
rect 15804 8984 15810 9036
rect 17773 9027 17831 9033
rect 17773 8993 17785 9027
rect 17819 9024 17831 9027
rect 17954 9024 17960 9036
rect 17819 8996 17960 9024
rect 17819 8993 17831 8996
rect 17773 8987 17831 8993
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 20806 8984 20812 9036
rect 20864 9024 20870 9036
rect 20936 9027 20994 9033
rect 20936 9024 20948 9027
rect 20864 8996 20948 9024
rect 20864 8984 20870 8996
rect 20936 8993 20948 8996
rect 20982 8993 20994 9027
rect 22462 9024 22468 9036
rect 22423 8996 22468 9024
rect 20936 8987 20994 8993
rect 22462 8984 22468 8996
rect 22520 8984 22526 9036
rect 22848 9033 22876 9064
rect 23014 9052 23020 9064
rect 23072 9052 23078 9104
rect 23658 9052 23664 9104
rect 23716 9092 23722 9104
rect 24166 9095 24224 9101
rect 24166 9092 24178 9095
rect 23716 9064 24178 9092
rect 23716 9052 23722 9064
rect 24166 9061 24178 9064
rect 24212 9061 24224 9095
rect 25498 9092 25504 9104
rect 25459 9064 25504 9092
rect 24166 9055 24224 9061
rect 25498 9052 25504 9064
rect 25556 9052 25562 9104
rect 26326 9092 26332 9104
rect 26287 9064 26332 9092
rect 26326 9052 26332 9064
rect 26384 9052 26390 9104
rect 28810 9052 28816 9104
rect 28868 9092 28874 9104
rect 28950 9095 29008 9101
rect 28950 9092 28962 9095
rect 28868 9064 28962 9092
rect 28868 9052 28874 9064
rect 28950 9061 28962 9064
rect 28996 9061 29008 9095
rect 28950 9055 29008 9061
rect 31205 9095 31263 9101
rect 31205 9061 31217 9095
rect 31251 9092 31263 9095
rect 32766 9092 32772 9104
rect 31251 9064 32772 9092
rect 31251 9061 31263 9064
rect 31205 9055 31263 9061
rect 32766 9052 32772 9064
rect 32824 9092 32830 9104
rect 33137 9095 33195 9101
rect 33137 9092 33149 9095
rect 32824 9064 33149 9092
rect 32824 9052 32830 9064
rect 33137 9061 33149 9064
rect 33183 9061 33195 9095
rect 33137 9055 33195 9061
rect 22833 9027 22891 9033
rect 22833 8993 22845 9027
rect 22879 9024 22891 9027
rect 22922 9024 22928 9036
rect 22879 8996 22928 9024
rect 22879 8993 22891 8996
rect 22833 8987 22891 8993
rect 22922 8984 22928 8996
rect 22980 8984 22986 9036
rect 24765 9027 24823 9033
rect 24765 8993 24777 9027
rect 24811 9024 24823 9027
rect 24854 9024 24860 9036
rect 24811 8996 24860 9024
rect 24811 8993 24823 8996
rect 24765 8987 24823 8993
rect 24854 8984 24860 8996
rect 24912 8984 24918 9036
rect 26510 9024 26516 9036
rect 26471 8996 26516 9024
rect 26510 8984 26516 8996
rect 26568 8984 26574 9036
rect 27062 9024 27068 9036
rect 27023 8996 27068 9024
rect 27062 8984 27068 8996
rect 27120 8984 27126 9036
rect 28350 8984 28356 9036
rect 28408 9024 28414 9036
rect 28629 9027 28687 9033
rect 28629 9024 28641 9027
rect 28408 8996 28641 9024
rect 28408 8984 28414 8996
rect 28629 8993 28641 8996
rect 28675 8993 28687 9027
rect 30558 9024 30564 9036
rect 30519 8996 30564 9024
rect 28629 8987 28687 8993
rect 30558 8984 30564 8996
rect 30616 8984 30622 9036
rect 30926 9024 30932 9036
rect 30887 8996 30932 9024
rect 30926 8984 30932 8996
rect 30984 8984 30990 9036
rect 32122 9024 32128 9036
rect 32083 8996 32128 9024
rect 32122 8984 32128 8996
rect 32180 8984 32186 9036
rect 32398 8984 32404 9036
rect 32456 9024 32462 9036
rect 32585 9027 32643 9033
rect 32585 9024 32597 9027
rect 32456 8996 32597 9024
rect 32456 8984 32462 8996
rect 32585 8993 32597 8996
rect 32631 9024 32643 9027
rect 33318 9024 33324 9036
rect 32631 8996 33324 9024
rect 32631 8993 32643 8996
rect 32585 8987 32643 8993
rect 33318 8984 33324 8996
rect 33376 8984 33382 9036
rect 34330 8984 34336 9036
rect 34388 9024 34394 9036
rect 34609 9027 34667 9033
rect 34609 9024 34621 9027
rect 34388 8996 34621 9024
rect 34388 8984 34394 8996
rect 34609 8993 34621 8996
rect 34655 9024 34667 9027
rect 34698 9024 34704 9036
rect 34655 8996 34704 9024
rect 34655 8993 34667 8996
rect 34609 8987 34667 8993
rect 34698 8984 34704 8996
rect 34756 9024 34762 9036
rect 36648 9024 36676 9120
rect 34756 8996 36676 9024
rect 34756 8984 34762 8996
rect 2498 8956 2504 8968
rect 2459 8928 2504 8956
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 2958 8916 2964 8968
rect 3016 8956 3022 8968
rect 3145 8959 3203 8965
rect 3145 8956 3157 8959
rect 3016 8928 3157 8956
rect 3016 8916 3022 8928
rect 3145 8925 3157 8928
rect 3191 8956 3203 8959
rect 4709 8959 4767 8965
rect 4709 8956 4721 8959
rect 3191 8928 4721 8956
rect 3191 8925 3203 8928
rect 3145 8919 3203 8925
rect 4709 8925 4721 8928
rect 4755 8956 4767 8959
rect 4798 8956 4804 8968
rect 4755 8928 4804 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 4798 8916 4804 8928
rect 4856 8956 4862 8968
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 4856 8928 4997 8956
rect 4856 8916 4862 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 5166 8916 5172 8968
rect 5224 8956 5230 8968
rect 5261 8959 5319 8965
rect 5261 8956 5273 8959
rect 5224 8928 5273 8956
rect 5224 8916 5230 8928
rect 5261 8925 5273 8928
rect 5307 8956 5319 8959
rect 6825 8959 6883 8965
rect 6825 8956 6837 8959
rect 5307 8928 6837 8956
rect 5307 8925 5319 8928
rect 5261 8919 5319 8925
rect 6825 8925 6837 8928
rect 6871 8925 6883 8959
rect 11054 8956 11060 8968
rect 11015 8928 11060 8956
rect 6825 8919 6883 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 13170 8916 13176 8968
rect 13228 8956 13234 8968
rect 13725 8959 13783 8965
rect 13725 8956 13737 8959
rect 13228 8928 13737 8956
rect 13228 8916 13234 8928
rect 13725 8925 13737 8928
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8956 23903 8959
rect 25130 8956 25136 8968
rect 23891 8928 25136 8956
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 25130 8916 25136 8928
rect 25188 8916 25194 8968
rect 32861 8959 32919 8965
rect 32861 8925 32873 8959
rect 32907 8956 32919 8959
rect 33505 8959 33563 8965
rect 33505 8956 33517 8959
rect 32907 8928 33517 8956
rect 32907 8925 32919 8928
rect 32861 8919 32919 8925
rect 33505 8925 33517 8928
rect 33551 8956 33563 8959
rect 33689 8959 33747 8965
rect 33689 8956 33701 8959
rect 33551 8928 33701 8956
rect 33551 8925 33563 8928
rect 33505 8919 33563 8925
rect 33689 8925 33701 8928
rect 33735 8925 33747 8959
rect 33689 8919 33747 8925
rect 33778 8916 33784 8968
rect 33836 8956 33842 8968
rect 35437 8959 35495 8965
rect 35437 8956 35449 8959
rect 33836 8928 35449 8956
rect 33836 8916 33842 8928
rect 35437 8925 35449 8928
rect 35483 8956 35495 8959
rect 36262 8956 36268 8968
rect 35483 8928 36268 8956
rect 35483 8925 35495 8928
rect 35437 8919 35495 8925
rect 36262 8916 36268 8928
rect 36320 8916 36326 8968
rect 2038 8848 2044 8900
rect 2096 8888 2102 8900
rect 2096 8860 4154 8888
rect 2096 8848 2102 8860
rect 1535 8823 1593 8829
rect 1535 8789 1547 8823
rect 1581 8820 1593 8823
rect 1854 8820 1860 8832
rect 1581 8792 1860 8820
rect 1581 8789 1593 8792
rect 1535 8783 1593 8789
rect 1854 8780 1860 8792
rect 1912 8780 1918 8832
rect 2314 8820 2320 8832
rect 2275 8792 2320 8820
rect 2314 8780 2320 8792
rect 2372 8780 2378 8832
rect 4126 8820 4154 8860
rect 5534 8848 5540 8900
rect 5592 8888 5598 8900
rect 7834 8888 7840 8900
rect 5592 8860 7840 8888
rect 5592 8848 5598 8860
rect 7834 8848 7840 8860
rect 7892 8848 7898 8900
rect 19518 8888 19524 8900
rect 19479 8860 19524 8888
rect 19518 8848 19524 8860
rect 19576 8848 19582 8900
rect 33410 8848 33416 8900
rect 33468 8888 33474 8900
rect 39574 8888 39580 8900
rect 33468 8860 39580 8888
rect 33468 8848 33474 8860
rect 39574 8848 39580 8860
rect 39632 8848 39638 8900
rect 4706 8820 4712 8832
rect 4126 8792 4712 8820
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 9125 8823 9183 8829
rect 9125 8820 9137 8823
rect 8812 8792 9137 8820
rect 8812 8780 8818 8792
rect 9125 8789 9137 8792
rect 9171 8820 9183 8823
rect 10594 8820 10600 8832
rect 9171 8792 10600 8820
rect 9171 8789 9183 8792
rect 9125 8783 9183 8789
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 12802 8820 12808 8832
rect 12763 8792 12808 8820
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 13446 8820 13452 8832
rect 13407 8792 13452 8820
rect 13446 8780 13452 8792
rect 13504 8820 13510 8832
rect 13722 8820 13728 8832
rect 13504 8792 13728 8820
rect 13504 8780 13510 8792
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 18003 8823 18061 8829
rect 18003 8789 18015 8823
rect 18049 8820 18061 8823
rect 18230 8820 18236 8832
rect 18049 8792 18236 8820
rect 18049 8789 18061 8792
rect 18003 8783 18061 8789
rect 18230 8780 18236 8792
rect 18288 8780 18294 8832
rect 18414 8820 18420 8832
rect 18375 8792 18420 8820
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 20714 8780 20720 8832
rect 20772 8820 20778 8832
rect 21039 8823 21097 8829
rect 21039 8820 21051 8823
rect 20772 8792 21051 8820
rect 20772 8780 20778 8792
rect 21039 8789 21051 8792
rect 21085 8789 21097 8823
rect 21542 8820 21548 8832
rect 21503 8792 21548 8820
rect 21039 8783 21097 8789
rect 21542 8780 21548 8792
rect 21600 8780 21606 8832
rect 23658 8820 23664 8832
rect 23619 8792 23664 8820
rect 23658 8780 23664 8792
rect 23716 8780 23722 8832
rect 27706 8820 27712 8832
rect 27667 8792 27712 8820
rect 27706 8780 27712 8792
rect 27764 8780 27770 8832
rect 30101 8823 30159 8829
rect 30101 8789 30113 8823
rect 30147 8820 30159 8823
rect 30190 8820 30196 8832
rect 30147 8792 30196 8820
rect 30147 8789 30159 8792
rect 30101 8783 30159 8789
rect 30190 8780 30196 8792
rect 30248 8780 30254 8832
rect 34974 8820 34980 8832
rect 34935 8792 34980 8820
rect 34974 8780 34980 8792
rect 35032 8780 35038 8832
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 1670 8616 1676 8628
rect 1631 8588 1676 8616
rect 1670 8576 1676 8588
rect 1728 8576 1734 8628
rect 2590 8576 2596 8628
rect 2648 8616 2654 8628
rect 3142 8616 3148 8628
rect 2648 8588 3148 8616
rect 2648 8576 2654 8588
rect 3142 8576 3148 8588
rect 3200 8616 3206 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 3200 8588 3249 8616
rect 3200 8576 3206 8588
rect 3237 8585 3249 8588
rect 3283 8585 3295 8619
rect 3970 8616 3976 8628
rect 3931 8588 3976 8616
rect 3237 8579 3295 8585
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 6273 8619 6331 8625
rect 6273 8585 6285 8619
rect 6319 8616 6331 8619
rect 6546 8616 6552 8628
rect 6319 8588 6552 8616
rect 6319 8585 6331 8588
rect 6273 8579 6331 8585
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 8110 8616 8116 8628
rect 8071 8588 8116 8616
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 8478 8616 8484 8628
rect 8439 8588 8484 8616
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 9030 8576 9036 8628
rect 9088 8616 9094 8628
rect 9171 8619 9229 8625
rect 9171 8616 9183 8619
rect 9088 8588 9183 8616
rect 9088 8576 9094 8588
rect 9171 8585 9183 8588
rect 9217 8585 9229 8619
rect 9950 8616 9956 8628
rect 9911 8588 9956 8616
rect 9171 8579 9229 8585
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 10652 8588 10977 8616
rect 10652 8576 10658 8588
rect 10965 8585 10977 8588
rect 11011 8585 11023 8619
rect 10965 8579 11023 8585
rect 11054 8576 11060 8628
rect 11112 8616 11118 8628
rect 11701 8619 11759 8625
rect 11701 8616 11713 8619
rect 11112 8588 11713 8616
rect 11112 8576 11118 8588
rect 11701 8585 11713 8588
rect 11747 8616 11759 8619
rect 12526 8616 12532 8628
rect 11747 8588 12532 8616
rect 11747 8585 11759 8588
rect 11701 8579 11759 8585
rect 12526 8576 12532 8588
rect 12584 8576 12590 8628
rect 13725 8619 13783 8625
rect 13725 8585 13737 8619
rect 13771 8616 13783 8619
rect 13814 8616 13820 8628
rect 13771 8588 13820 8616
rect 13771 8585 13783 8588
rect 13725 8579 13783 8585
rect 13814 8576 13820 8588
rect 13872 8616 13878 8628
rect 14001 8619 14059 8625
rect 14001 8616 14013 8619
rect 13872 8588 14013 8616
rect 13872 8576 13878 8588
rect 14001 8585 14013 8588
rect 14047 8585 14059 8619
rect 14001 8579 14059 8585
rect 15746 8576 15752 8628
rect 15804 8616 15810 8628
rect 17313 8619 17371 8625
rect 17313 8616 17325 8619
rect 15804 8588 17325 8616
rect 15804 8576 15810 8588
rect 17313 8585 17325 8588
rect 17359 8585 17371 8619
rect 19242 8616 19248 8628
rect 19203 8588 19248 8616
rect 17313 8579 17371 8585
rect 19242 8576 19248 8588
rect 19300 8576 19306 8628
rect 20622 8616 20628 8628
rect 20583 8588 20628 8616
rect 20622 8576 20628 8588
rect 20680 8576 20686 8628
rect 20806 8576 20812 8628
rect 20864 8616 20870 8628
rect 20901 8619 20959 8625
rect 20901 8616 20913 8619
rect 20864 8588 20913 8616
rect 20864 8576 20870 8588
rect 20901 8585 20913 8588
rect 20947 8585 20959 8619
rect 21266 8616 21272 8628
rect 21227 8588 21272 8616
rect 20901 8579 20959 8585
rect 21266 8576 21272 8588
rect 21324 8576 21330 8628
rect 24394 8576 24400 8628
rect 24452 8616 24458 8628
rect 24581 8619 24639 8625
rect 24581 8616 24593 8619
rect 24452 8588 24593 8616
rect 24452 8576 24458 8588
rect 24581 8585 24593 8588
rect 24627 8585 24639 8619
rect 24581 8579 24639 8585
rect 24949 8619 25007 8625
rect 24949 8585 24961 8619
rect 24995 8616 25007 8619
rect 25130 8616 25136 8628
rect 24995 8588 25136 8616
rect 24995 8585 25007 8588
rect 24949 8579 25007 8585
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 25406 8576 25412 8628
rect 25464 8616 25470 8628
rect 25501 8619 25559 8625
rect 25501 8616 25513 8619
rect 25464 8588 25513 8616
rect 25464 8576 25470 8588
rect 25501 8585 25513 8588
rect 25547 8585 25559 8619
rect 27062 8616 27068 8628
rect 27023 8588 27068 8616
rect 25501 8579 25559 8585
rect 2498 8508 2504 8560
rect 2556 8548 2562 8560
rect 3605 8551 3663 8557
rect 3605 8548 3617 8551
rect 2556 8520 3617 8548
rect 2556 8508 2562 8520
rect 3605 8517 3617 8520
rect 3651 8517 3663 8551
rect 3605 8511 3663 8517
rect 5166 8508 5172 8560
rect 5224 8548 5230 8560
rect 15473 8551 15531 8557
rect 5224 8520 5580 8548
rect 5224 8508 5230 8520
rect 1854 8440 1860 8492
rect 1912 8480 1918 8492
rect 2317 8483 2375 8489
rect 2317 8480 2329 8483
rect 1912 8452 2329 8480
rect 1912 8440 1918 8452
rect 2317 8449 2329 8452
rect 2363 8449 2375 8483
rect 2958 8480 2964 8492
rect 2919 8452 2964 8480
rect 2317 8443 2375 8449
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5442 8480 5448 8492
rect 5307 8452 5448 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 5552 8489 5580 8520
rect 15473 8517 15485 8551
rect 15519 8548 15531 8551
rect 15519 8520 17264 8548
rect 15519 8517 15531 8520
rect 15473 8511 15531 8517
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8449 5595 8483
rect 6914 8480 6920 8492
rect 6875 8452 6920 8480
rect 5537 8443 5595 8449
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 10045 8483 10103 8489
rect 10045 8449 10057 8483
rect 10091 8480 10103 8483
rect 10778 8480 10784 8492
rect 10091 8452 10784 8480
rect 10091 8449 10103 8452
rect 10045 8443 10103 8449
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 16114 8480 16120 8492
rect 16075 8452 16120 8480
rect 16114 8440 16120 8452
rect 16172 8480 16178 8492
rect 17126 8480 17132 8492
rect 16172 8452 17132 8480
rect 16172 8440 16178 8452
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8412 3847 8415
rect 4433 8415 4491 8421
rect 4433 8412 4445 8415
rect 3835 8384 4445 8412
rect 3835 8381 3847 8384
rect 3789 8375 3847 8381
rect 4433 8381 4445 8384
rect 4479 8412 4491 8415
rect 4614 8412 4620 8424
rect 4479 8384 4620 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 4614 8372 4620 8384
rect 4672 8372 4678 8424
rect 9068 8415 9126 8421
rect 9068 8412 9080 8415
rect 6472 8384 9080 8412
rect 2133 8347 2191 8353
rect 2133 8313 2145 8347
rect 2179 8344 2191 8347
rect 2314 8344 2320 8356
rect 2179 8316 2320 8344
rect 2179 8313 2191 8316
rect 2133 8307 2191 8313
rect 2314 8304 2320 8316
rect 2372 8344 2378 8356
rect 2409 8347 2467 8353
rect 2409 8344 2421 8347
rect 2372 8316 2421 8344
rect 2372 8304 2378 8316
rect 2409 8313 2421 8316
rect 2455 8344 2467 8347
rect 2682 8344 2688 8356
rect 2455 8316 2688 8344
rect 2455 8313 2467 8316
rect 2409 8307 2467 8313
rect 2682 8304 2688 8316
rect 2740 8304 2746 8356
rect 5077 8347 5135 8353
rect 5077 8313 5089 8347
rect 5123 8344 5135 8347
rect 5350 8344 5356 8356
rect 5123 8316 5356 8344
rect 5123 8313 5135 8316
rect 5077 8307 5135 8313
rect 5350 8304 5356 8316
rect 5408 8304 5414 8356
rect 6472 8344 6500 8384
rect 9068 8381 9080 8384
rect 9114 8412 9126 8415
rect 9490 8412 9496 8424
rect 9114 8384 9496 8412
rect 9114 8381 9126 8384
rect 9068 8375 9126 8381
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 12802 8412 12808 8424
rect 11296 8384 12808 8412
rect 11296 8372 11302 8384
rect 12802 8372 12808 8384
rect 12860 8372 12866 8424
rect 14553 8415 14611 8421
rect 14553 8381 14565 8415
rect 14599 8412 14611 8415
rect 14642 8412 14648 8424
rect 14599 8384 14648 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 14642 8372 14648 8384
rect 14700 8372 14706 8424
rect 16316 8421 16344 8452
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 16301 8415 16359 8421
rect 16301 8381 16313 8415
rect 16347 8381 16359 8415
rect 16850 8412 16856 8424
rect 16811 8384 16856 8412
rect 16301 8375 16359 8381
rect 16850 8372 16856 8384
rect 16908 8372 16914 8424
rect 5644 8316 6500 8344
rect 6641 8347 6699 8353
rect 4706 8236 4712 8288
rect 4764 8276 4770 8288
rect 5644 8276 5672 8316
rect 6641 8313 6653 8347
rect 6687 8344 6699 8347
rect 7190 8344 7196 8356
rect 6687 8316 7196 8344
rect 6687 8313 6699 8316
rect 6641 8307 6699 8313
rect 7190 8304 7196 8316
rect 7248 8353 7254 8356
rect 7248 8347 7296 8353
rect 7248 8313 7250 8347
rect 7284 8313 7296 8347
rect 7248 8307 7296 8313
rect 7248 8304 7254 8307
rect 9766 8304 9772 8356
rect 9824 8344 9830 8356
rect 10366 8347 10424 8353
rect 10366 8344 10378 8347
rect 9824 8316 10378 8344
rect 9824 8304 9830 8316
rect 10366 8313 10378 8316
rect 10412 8344 10424 8347
rect 11333 8347 11391 8353
rect 11333 8344 11345 8347
rect 10412 8316 11345 8344
rect 10412 8313 10424 8316
rect 10366 8307 10424 8313
rect 11333 8313 11345 8316
rect 11379 8344 11391 8347
rect 11422 8344 11428 8356
rect 11379 8316 11428 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 11422 8304 11428 8316
rect 11480 8344 11486 8356
rect 12621 8347 12679 8353
rect 12621 8344 12633 8347
rect 11480 8316 12633 8344
rect 11480 8304 11486 8316
rect 12621 8313 12633 8316
rect 12667 8344 12679 8347
rect 13126 8347 13184 8353
rect 13126 8344 13138 8347
rect 12667 8316 13138 8344
rect 12667 8313 12679 8316
rect 12621 8307 12679 8313
rect 13126 8313 13138 8316
rect 13172 8344 13184 8347
rect 14915 8347 14973 8353
rect 13172 8316 13814 8344
rect 13172 8313 13184 8316
rect 13126 8307 13184 8313
rect 4764 8248 5672 8276
rect 4764 8236 4770 8248
rect 6822 8236 6828 8288
rect 6880 8276 6886 8288
rect 7837 8279 7895 8285
rect 7837 8276 7849 8279
rect 6880 8248 7849 8276
rect 6880 8236 6886 8248
rect 7837 8245 7849 8248
rect 7883 8245 7895 8279
rect 13786 8276 13814 8316
rect 14915 8313 14927 8347
rect 14961 8313 14973 8347
rect 17034 8344 17040 8356
rect 16995 8316 17040 8344
rect 14915 8307 14973 8313
rect 14461 8279 14519 8285
rect 14461 8276 14473 8279
rect 13786 8248 14473 8276
rect 7837 8239 7895 8245
rect 14461 8245 14473 8248
rect 14507 8276 14519 8279
rect 14930 8276 14958 8307
rect 17034 8304 17040 8316
rect 17092 8304 17098 8356
rect 17236 8344 17264 8520
rect 17310 8440 17316 8492
rect 17368 8480 17374 8492
rect 18233 8483 18291 8489
rect 18233 8480 18245 8483
rect 17368 8452 18245 8480
rect 17368 8440 17374 8452
rect 18233 8449 18245 8452
rect 18279 8480 18291 8483
rect 18506 8480 18512 8492
rect 18279 8452 18512 8480
rect 18279 8449 18291 8452
rect 18233 8443 18291 8449
rect 18506 8440 18512 8452
rect 18564 8440 18570 8492
rect 18598 8440 18604 8492
rect 18656 8480 18662 8492
rect 19260 8480 19288 8576
rect 19705 8483 19763 8489
rect 19705 8480 19717 8483
rect 18656 8452 18701 8480
rect 19260 8452 19717 8480
rect 18656 8440 18662 8452
rect 19705 8449 19717 8452
rect 19751 8449 19763 8483
rect 25516 8480 25544 8579
rect 27062 8576 27068 8588
rect 27120 8576 27126 8628
rect 28350 8576 28356 8628
rect 28408 8616 28414 8628
rect 28997 8619 29055 8625
rect 28997 8616 29009 8619
rect 28408 8588 29009 8616
rect 28408 8576 28414 8588
rect 28997 8585 29009 8588
rect 29043 8585 29055 8619
rect 28997 8579 29055 8585
rect 31202 8576 31208 8628
rect 31260 8616 31266 8628
rect 31711 8619 31769 8625
rect 31711 8616 31723 8619
rect 31260 8588 31723 8616
rect 31260 8576 31266 8588
rect 31711 8585 31723 8588
rect 31757 8585 31769 8619
rect 34054 8616 34060 8628
rect 33967 8588 34060 8616
rect 31711 8579 31769 8585
rect 34054 8576 34060 8588
rect 34112 8616 34118 8628
rect 35802 8616 35808 8628
rect 34112 8588 35808 8616
rect 34112 8576 34118 8588
rect 35802 8576 35808 8588
rect 35860 8616 35866 8628
rect 35897 8619 35955 8625
rect 35897 8616 35909 8619
rect 35860 8588 35909 8616
rect 35860 8576 35866 8588
rect 35897 8585 35909 8588
rect 35943 8585 35955 8619
rect 36262 8616 36268 8628
rect 36223 8588 36268 8616
rect 35897 8579 35955 8585
rect 36262 8576 36268 8588
rect 36320 8576 36326 8628
rect 36630 8616 36636 8628
rect 36591 8588 36636 8616
rect 36630 8576 36636 8588
rect 36688 8576 36694 8628
rect 30282 8548 30288 8560
rect 28092 8520 30288 8548
rect 25777 8483 25835 8489
rect 25777 8480 25789 8483
rect 25516 8452 25789 8480
rect 19705 8443 19763 8449
rect 25777 8449 25789 8452
rect 25823 8449 25835 8483
rect 25777 8443 25835 8449
rect 26421 8483 26479 8489
rect 26421 8449 26433 8483
rect 26467 8480 26479 8483
rect 26970 8480 26976 8492
rect 26467 8452 26976 8480
rect 26467 8449 26479 8452
rect 26421 8443 26479 8449
rect 26970 8440 26976 8452
rect 27028 8440 27034 8492
rect 17865 8415 17923 8421
rect 17865 8381 17877 8415
rect 17911 8412 17923 8415
rect 17954 8412 17960 8424
rect 17911 8384 17960 8412
rect 17911 8381 17923 8384
rect 17865 8375 17923 8381
rect 17954 8372 17960 8384
rect 18012 8372 18018 8424
rect 21266 8372 21272 8424
rect 21324 8412 21330 8424
rect 21453 8415 21511 8421
rect 21453 8412 21465 8415
rect 21324 8384 21465 8412
rect 21324 8372 21330 8384
rect 21453 8381 21465 8384
rect 21499 8381 21511 8415
rect 21453 8375 21511 8381
rect 21542 8372 21548 8424
rect 21600 8412 21606 8424
rect 21913 8415 21971 8421
rect 21913 8412 21925 8415
rect 21600 8384 21925 8412
rect 21600 8372 21606 8384
rect 21913 8381 21925 8384
rect 21959 8381 21971 8415
rect 21913 8375 21971 8381
rect 23661 8415 23719 8421
rect 23661 8381 23673 8415
rect 23707 8412 23719 8415
rect 24210 8412 24216 8424
rect 23707 8384 24216 8412
rect 23707 8381 23719 8384
rect 23661 8375 23719 8381
rect 24210 8372 24216 8384
rect 24268 8372 24274 8424
rect 27522 8412 27528 8424
rect 27435 8384 27528 8412
rect 18325 8347 18383 8353
rect 18325 8344 18337 8347
rect 17236 8316 18337 8344
rect 18325 8313 18337 8316
rect 18371 8344 18383 8347
rect 18414 8344 18420 8356
rect 18371 8316 18420 8344
rect 18371 8313 18383 8316
rect 18325 8307 18383 8313
rect 18414 8304 18420 8316
rect 18472 8344 18478 8356
rect 19242 8344 19248 8356
rect 18472 8316 19248 8344
rect 18472 8304 18478 8316
rect 19242 8304 19248 8316
rect 19300 8304 19306 8356
rect 19613 8347 19671 8353
rect 19613 8313 19625 8347
rect 19659 8344 19671 8347
rect 20067 8347 20125 8353
rect 20067 8344 20079 8347
rect 19659 8316 20079 8344
rect 19659 8313 19671 8316
rect 19613 8307 19671 8313
rect 20067 8313 20079 8316
rect 20113 8344 20125 8347
rect 20113 8316 20346 8344
rect 20113 8313 20125 8316
rect 20067 8307 20125 8313
rect 15746 8276 15752 8288
rect 14507 8248 15752 8276
rect 14507 8245 14519 8248
rect 14461 8239 14519 8245
rect 15746 8236 15752 8248
rect 15804 8236 15810 8288
rect 17862 8236 17868 8288
rect 17920 8276 17926 8288
rect 19058 8276 19064 8288
rect 17920 8248 19064 8276
rect 17920 8236 17926 8248
rect 19058 8236 19064 8248
rect 19116 8236 19122 8288
rect 20318 8276 20346 8316
rect 20530 8304 20536 8356
rect 20588 8344 20594 8356
rect 21560 8344 21588 8372
rect 23750 8344 23756 8356
rect 20588 8316 21588 8344
rect 22480 8316 23756 8344
rect 20588 8304 20594 8316
rect 22480 8288 22508 8316
rect 23750 8304 23756 8316
rect 23808 8304 23814 8356
rect 24023 8347 24081 8353
rect 24023 8313 24035 8347
rect 24069 8313 24081 8347
rect 24023 8307 24081 8313
rect 21358 8276 21364 8288
rect 20318 8248 21364 8276
rect 21358 8236 21364 8248
rect 21416 8236 21422 8288
rect 21542 8276 21548 8288
rect 21503 8248 21548 8276
rect 21542 8236 21548 8248
rect 21600 8236 21606 8288
rect 22462 8276 22468 8288
rect 22423 8248 22468 8276
rect 22462 8236 22468 8248
rect 22520 8236 22526 8288
rect 22922 8276 22928 8288
rect 22883 8248 22928 8276
rect 22922 8236 22928 8248
rect 22980 8236 22986 8288
rect 23477 8279 23535 8285
rect 23477 8245 23489 8279
rect 23523 8276 23535 8279
rect 23658 8276 23664 8288
rect 23523 8248 23664 8276
rect 23523 8245 23535 8248
rect 23477 8239 23535 8245
rect 23658 8236 23664 8248
rect 23716 8276 23722 8288
rect 24038 8276 24066 8307
rect 25866 8304 25872 8356
rect 25924 8344 25930 8356
rect 25924 8316 25969 8344
rect 25924 8304 25930 8316
rect 24670 8276 24676 8288
rect 23716 8248 24676 8276
rect 23716 8236 23722 8248
rect 24670 8236 24676 8248
rect 24728 8236 24734 8288
rect 25130 8236 25136 8288
rect 25188 8276 25194 8288
rect 26510 8276 26516 8288
rect 25188 8248 26516 8276
rect 25188 8236 25194 8248
rect 26510 8236 26516 8248
rect 26568 8276 26574 8288
rect 27448 8285 27476 8384
rect 27522 8372 27528 8384
rect 27580 8412 27586 8424
rect 27617 8415 27675 8421
rect 27617 8412 27629 8415
rect 27580 8384 27629 8412
rect 27580 8372 27586 8384
rect 27617 8381 27629 8384
rect 27663 8381 27675 8415
rect 27617 8375 27675 8381
rect 27706 8372 27712 8424
rect 27764 8412 27770 8424
rect 28092 8421 28120 8520
rect 30282 8508 30288 8520
rect 30340 8548 30346 8560
rect 30926 8548 30932 8560
rect 30340 8520 30932 8548
rect 30340 8508 30346 8520
rect 30926 8508 30932 8520
rect 30984 8548 30990 8560
rect 31021 8551 31079 8557
rect 31021 8548 31033 8551
rect 30984 8520 31033 8548
rect 30984 8508 30990 8520
rect 31021 8517 31033 8520
rect 31067 8517 31079 8551
rect 31021 8511 31079 8517
rect 30745 8483 30803 8489
rect 30745 8449 30757 8483
rect 30791 8480 30803 8483
rect 31481 8483 31539 8489
rect 31481 8480 31493 8483
rect 30791 8452 31493 8480
rect 30791 8449 30803 8452
rect 30745 8443 30803 8449
rect 31481 8449 31493 8452
rect 31527 8480 31539 8483
rect 35253 8483 35311 8489
rect 35253 8480 35265 8483
rect 31527 8452 35265 8480
rect 31527 8449 31539 8452
rect 31481 8443 31539 8449
rect 31680 8421 31708 8452
rect 35253 8449 35265 8452
rect 35299 8480 35311 8483
rect 35618 8480 35624 8492
rect 35299 8452 35624 8480
rect 35299 8449 35311 8452
rect 35253 8443 35311 8449
rect 35618 8440 35624 8452
rect 35676 8440 35682 8492
rect 28077 8415 28135 8421
rect 28077 8412 28089 8415
rect 27764 8384 28089 8412
rect 27764 8372 27770 8384
rect 28077 8381 28089 8384
rect 28123 8381 28135 8415
rect 28077 8375 28135 8381
rect 31640 8415 31708 8421
rect 31640 8381 31652 8415
rect 31686 8384 31708 8415
rect 32766 8412 32772 8424
rect 32727 8384 32772 8412
rect 31686 8381 31698 8384
rect 31640 8375 31698 8381
rect 32766 8372 32772 8384
rect 32824 8372 32830 8424
rect 33689 8415 33747 8421
rect 33689 8381 33701 8415
rect 33735 8412 33747 8415
rect 34609 8415 34667 8421
rect 34609 8412 34621 8415
rect 33735 8384 34621 8412
rect 33735 8381 33747 8384
rect 33689 8375 33747 8381
rect 34609 8381 34621 8384
rect 34655 8381 34667 8415
rect 34609 8375 34667 8381
rect 28353 8347 28411 8353
rect 28353 8313 28365 8347
rect 28399 8344 28411 8347
rect 29638 8344 29644 8356
rect 28399 8316 29644 8344
rect 28399 8313 28411 8316
rect 28353 8307 28411 8313
rect 29638 8304 29644 8316
rect 29696 8304 29702 8356
rect 29917 8347 29975 8353
rect 29917 8313 29929 8347
rect 29963 8344 29975 8347
rect 30098 8344 30104 8356
rect 29963 8316 30104 8344
rect 29963 8313 29975 8316
rect 29917 8307 29975 8313
rect 30098 8304 30104 8316
rect 30156 8304 30162 8356
rect 30190 8304 30196 8356
rect 30248 8344 30254 8356
rect 30248 8316 30293 8344
rect 30248 8304 30254 8316
rect 32030 8304 32036 8356
rect 32088 8344 32094 8356
rect 32585 8347 32643 8353
rect 32585 8344 32597 8347
rect 32088 8316 32597 8344
rect 32088 8304 32094 8316
rect 32585 8313 32597 8316
rect 32631 8344 32643 8347
rect 33131 8347 33189 8353
rect 33131 8344 33143 8347
rect 32631 8316 33143 8344
rect 32631 8313 32643 8316
rect 32585 8307 32643 8313
rect 33131 8313 33143 8316
rect 33177 8344 33189 8347
rect 34054 8344 34060 8356
rect 33177 8316 34060 8344
rect 33177 8313 33189 8316
rect 33131 8307 33189 8313
rect 34054 8304 34060 8316
rect 34112 8304 34118 8356
rect 26697 8279 26755 8285
rect 26697 8276 26709 8279
rect 26568 8248 26709 8276
rect 26568 8236 26574 8248
rect 26697 8245 26709 8248
rect 26743 8276 26755 8279
rect 27433 8279 27491 8285
rect 27433 8276 27445 8279
rect 26743 8248 27445 8276
rect 26743 8245 26755 8248
rect 26697 8239 26755 8245
rect 27433 8245 27445 8248
rect 27479 8245 27491 8279
rect 27433 8239 27491 8245
rect 28721 8279 28779 8285
rect 28721 8245 28733 8279
rect 28767 8276 28779 8279
rect 28810 8276 28816 8288
rect 28767 8248 28816 8276
rect 28767 8245 28779 8248
rect 28721 8239 28779 8245
rect 28810 8236 28816 8248
rect 28868 8236 28874 8288
rect 30466 8236 30472 8288
rect 30524 8276 30530 8288
rect 32122 8276 32128 8288
rect 30524 8248 32128 8276
rect 30524 8236 30530 8248
rect 32122 8236 32128 8248
rect 32180 8236 32186 8288
rect 34624 8276 34652 8375
rect 36262 8372 36268 8424
rect 36320 8412 36326 8424
rect 36449 8415 36507 8421
rect 36449 8412 36461 8415
rect 36320 8384 36461 8412
rect 36320 8372 36326 8384
rect 36449 8381 36461 8384
rect 36495 8412 36507 8415
rect 37001 8415 37059 8421
rect 37001 8412 37013 8415
rect 36495 8384 37013 8412
rect 36495 8381 36507 8384
rect 36449 8375 36507 8381
rect 37001 8381 37013 8384
rect 37047 8381 37059 8415
rect 37001 8375 37059 8381
rect 34974 8344 34980 8356
rect 34935 8316 34980 8344
rect 34974 8304 34980 8316
rect 35032 8304 35038 8356
rect 35069 8347 35127 8353
rect 35069 8313 35081 8347
rect 35115 8313 35127 8347
rect 35069 8307 35127 8313
rect 35084 8276 35112 8307
rect 34624 8248 35112 8276
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 2130 8072 2136 8084
rect 2091 8044 2136 8072
rect 2130 8032 2136 8044
rect 2188 8032 2194 8084
rect 2682 8072 2688 8084
rect 2643 8044 2688 8072
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 4062 8072 4068 8084
rect 3927 8044 4068 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 5810 8072 5816 8084
rect 5771 8044 5816 8072
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 6549 8075 6607 8081
rect 6549 8041 6561 8075
rect 6595 8072 6607 8075
rect 6638 8072 6644 8084
rect 6595 8044 6644 8072
rect 6595 8041 6607 8044
rect 6549 8035 6607 8041
rect 6638 8032 6644 8044
rect 6696 8072 6702 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 6696 8044 7757 8072
rect 6696 8032 6702 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 8711 8075 8769 8081
rect 8711 8041 8723 8075
rect 8757 8072 8769 8075
rect 12158 8072 12164 8084
rect 8757 8044 12164 8072
rect 8757 8041 8769 8044
rect 8711 8035 8769 8041
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 12618 8072 12624 8084
rect 12452 8044 12624 8072
rect 3513 8007 3571 8013
rect 3513 7973 3525 8007
rect 3559 8004 3571 8007
rect 3786 8004 3792 8016
rect 3559 7976 3792 8004
rect 3559 7973 3571 7976
rect 3513 7967 3571 7973
rect 3786 7964 3792 7976
rect 3844 8004 3850 8016
rect 4157 8007 4215 8013
rect 4157 8004 4169 8007
rect 3844 7976 4169 8004
rect 3844 7964 3850 7976
rect 4157 7973 4169 7976
rect 4203 7973 4215 8007
rect 4157 7967 4215 7973
rect 4246 7964 4252 8016
rect 4304 8004 4310 8016
rect 4798 8004 4804 8016
rect 4304 7976 4349 8004
rect 4759 7976 4804 8004
rect 4304 7964 4310 7976
rect 4798 7964 4804 7976
rect 4856 7964 4862 8016
rect 5074 7964 5080 8016
rect 5132 8004 5138 8016
rect 5169 8007 5227 8013
rect 5169 8004 5181 8007
rect 5132 7976 5181 8004
rect 5132 7964 5138 7976
rect 5169 7973 5181 7976
rect 5215 8004 5227 8007
rect 6822 8004 6828 8016
rect 5215 7976 6828 8004
rect 5215 7973 5227 7976
rect 5169 7967 5227 7973
rect 6822 7964 6828 7976
rect 6880 7964 6886 8016
rect 7190 8013 7196 8016
rect 7187 8004 7196 8013
rect 7151 7976 7196 8004
rect 7187 7967 7196 7976
rect 7190 7964 7196 7967
rect 7248 7964 7254 8016
rect 11238 8004 11244 8016
rect 11199 7976 11244 8004
rect 11238 7964 11244 7976
rect 11296 7964 11302 8016
rect 12452 8004 12480 8044
rect 12618 8032 12624 8044
rect 12676 8072 12682 8084
rect 12986 8072 12992 8084
rect 12676 8044 12992 8072
rect 12676 8032 12682 8044
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 13170 8072 13176 8084
rect 13131 8044 13176 8072
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 16945 8075 17003 8081
rect 16945 8041 16957 8075
rect 16991 8072 17003 8075
rect 17034 8072 17040 8084
rect 16991 8044 17040 8072
rect 16991 8041 17003 8044
rect 16945 8035 17003 8041
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 18506 8072 18512 8084
rect 18467 8044 18512 8072
rect 18506 8032 18512 8044
rect 18564 8032 18570 8084
rect 18969 8075 19027 8081
rect 18969 8041 18981 8075
rect 19015 8072 19027 8075
rect 19058 8072 19064 8084
rect 19015 8044 19064 8072
rect 19015 8041 19027 8044
rect 18969 8035 19027 8041
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 20073 8075 20131 8081
rect 20073 8072 20085 8075
rect 19168 8044 20085 8072
rect 14369 8007 14427 8013
rect 11348 7976 12480 8004
rect 12636 7976 13814 8004
rect 1762 7936 1768 7948
rect 1723 7908 1768 7936
rect 1762 7896 1768 7908
rect 1820 7896 1826 7948
rect 5626 7936 5632 7948
rect 5587 7908 5632 7936
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 8640 7939 8698 7945
rect 8640 7905 8652 7939
rect 8686 7936 8698 7939
rect 9030 7936 9036 7948
rect 8686 7908 9036 7936
rect 8686 7905 8698 7908
rect 8640 7899 8698 7905
rect 9030 7896 9036 7908
rect 9088 7896 9094 7948
rect 10778 7936 10784 7948
rect 10739 7908 10784 7936
rect 10778 7896 10784 7908
rect 10836 7896 10842 7948
rect 11057 7939 11115 7945
rect 11057 7905 11069 7939
rect 11103 7936 11115 7939
rect 11348 7936 11376 7976
rect 12066 7936 12072 7948
rect 11103 7908 11376 7936
rect 12027 7908 12072 7936
rect 11103 7905 11115 7908
rect 11057 7899 11115 7905
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 6914 7868 6920 7880
rect 6871 7840 6920 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 6914 7828 6920 7840
rect 6972 7828 6978 7880
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 10042 7868 10048 7880
rect 7432 7840 10048 7868
rect 7432 7828 7438 7840
rect 10042 7828 10048 7840
rect 10100 7868 10106 7880
rect 11072 7868 11100 7899
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 12158 7896 12164 7948
rect 12216 7936 12222 7948
rect 12636 7945 12664 7976
rect 12621 7939 12679 7945
rect 12621 7936 12633 7939
rect 12216 7908 12633 7936
rect 12216 7896 12222 7908
rect 12621 7905 12633 7908
rect 12667 7905 12679 7939
rect 13630 7936 13636 7948
rect 13591 7908 13636 7936
rect 12621 7899 12679 7905
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 13786 7936 13814 7976
rect 14369 7973 14381 8007
rect 14415 8004 14427 8007
rect 14642 8004 14648 8016
rect 14415 7976 14648 8004
rect 14415 7973 14427 7976
rect 14369 7967 14427 7973
rect 14642 7964 14648 7976
rect 14700 7964 14706 8016
rect 15651 8007 15709 8013
rect 15651 7973 15663 8007
rect 15697 8004 15709 8007
rect 15746 8004 15752 8016
rect 15697 7976 15752 8004
rect 15697 7973 15709 7976
rect 15651 7967 15709 7973
rect 15746 7964 15752 7976
rect 15804 7964 15810 8016
rect 17586 8004 17592 8016
rect 17547 7976 17592 8004
rect 17586 7964 17592 7976
rect 17644 7964 17650 8016
rect 17681 8007 17739 8013
rect 17681 7973 17693 8007
rect 17727 8004 17739 8007
rect 17862 8004 17868 8016
rect 17727 7976 17868 8004
rect 17727 7973 17739 7976
rect 17681 7967 17739 7973
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 18230 7964 18236 8016
rect 18288 8004 18294 8016
rect 19168 8013 19196 8044
rect 20073 8041 20085 8044
rect 20119 8041 20131 8075
rect 20073 8035 20131 8041
rect 22922 8032 22928 8084
rect 22980 8072 22986 8084
rect 25409 8075 25467 8081
rect 22980 8044 23474 8072
rect 22980 8032 22986 8044
rect 19153 8007 19211 8013
rect 19153 8004 19165 8007
rect 18288 7976 19165 8004
rect 18288 7964 18294 7976
rect 19153 7973 19165 7976
rect 19199 7973 19211 8007
rect 19153 7967 19211 7973
rect 19242 7964 19248 8016
rect 19300 8004 19306 8016
rect 21634 8004 21640 8016
rect 19300 7976 19345 8004
rect 21595 7976 21640 8004
rect 19300 7964 19306 7976
rect 21634 7964 21640 7976
rect 21692 7964 21698 8016
rect 14090 7936 14096 7948
rect 13786 7908 14096 7936
rect 14090 7896 14096 7908
rect 14148 7936 14154 7948
rect 14185 7939 14243 7945
rect 14185 7936 14197 7939
rect 14148 7908 14197 7936
rect 14148 7896 14154 7908
rect 14185 7905 14197 7908
rect 14231 7936 14243 7939
rect 14231 7908 16160 7936
rect 14231 7905 14243 7908
rect 14185 7899 14243 7905
rect 10100 7840 11100 7868
rect 12805 7871 12863 7877
rect 10100 7828 10106 7840
rect 12805 7837 12817 7871
rect 12851 7868 12863 7871
rect 14550 7868 14556 7880
rect 12851 7840 14556 7868
rect 12851 7837 12863 7840
rect 12805 7831 12863 7837
rect 14550 7828 14556 7840
rect 14608 7868 14614 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 14608 7840 15301 7868
rect 14608 7828 14614 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 3053 7735 3111 7741
rect 3053 7701 3065 7735
rect 3099 7732 3111 7735
rect 3510 7732 3516 7744
rect 3099 7704 3516 7732
rect 3099 7701 3111 7704
rect 3053 7695 3111 7701
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 5442 7732 5448 7744
rect 5403 7704 5448 7732
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 9766 7692 9772 7744
rect 9824 7732 9830 7744
rect 10045 7735 10103 7741
rect 10045 7732 10057 7735
rect 9824 7704 10057 7732
rect 9824 7692 9830 7704
rect 10045 7701 10057 7704
rect 10091 7701 10103 7735
rect 10045 7695 10103 7701
rect 13541 7735 13599 7741
rect 13541 7701 13553 7735
rect 13587 7732 13599 7735
rect 13814 7732 13820 7744
rect 13587 7704 13820 7732
rect 13587 7701 13599 7704
rect 13541 7695 13599 7701
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 16132 7732 16160 7908
rect 22646 7896 22652 7948
rect 22704 7936 22710 7948
rect 23017 7939 23075 7945
rect 23017 7936 23029 7939
rect 22704 7908 23029 7936
rect 22704 7896 22710 7908
rect 23017 7905 23029 7908
rect 23063 7905 23075 7939
rect 23017 7899 23075 7905
rect 23106 7896 23112 7948
rect 23164 7936 23170 7948
rect 23201 7939 23259 7945
rect 23201 7936 23213 7939
rect 23164 7908 23213 7936
rect 23164 7896 23170 7908
rect 23201 7905 23213 7908
rect 23247 7905 23259 7939
rect 23446 7936 23474 8044
rect 25409 8041 25421 8075
rect 25455 8072 25467 8075
rect 25777 8075 25835 8081
rect 25777 8072 25789 8075
rect 25455 8044 25789 8072
rect 25455 8041 25467 8044
rect 25409 8035 25467 8041
rect 25777 8041 25789 8044
rect 25823 8072 25835 8075
rect 25866 8072 25872 8084
rect 25823 8044 25872 8072
rect 25823 8041 25835 8044
rect 25777 8035 25835 8041
rect 25866 8032 25872 8044
rect 25924 8032 25930 8084
rect 30098 8032 30104 8084
rect 30156 8072 30162 8084
rect 30653 8075 30711 8081
rect 30653 8072 30665 8075
rect 30156 8044 30665 8072
rect 30156 8032 30162 8044
rect 30653 8041 30665 8044
rect 30699 8041 30711 8075
rect 32398 8072 32404 8084
rect 32359 8044 32404 8072
rect 30653 8035 30711 8041
rect 32398 8032 32404 8044
rect 32456 8032 32462 8084
rect 34425 8075 34483 8081
rect 34425 8041 34437 8075
rect 34471 8072 34483 8075
rect 34471 8044 35480 8072
rect 34471 8041 34483 8044
rect 34425 8035 34483 8041
rect 35452 8016 35480 8044
rect 24670 7964 24676 8016
rect 24728 8004 24734 8016
rect 24810 8007 24868 8013
rect 24810 8004 24822 8007
rect 24728 7976 24822 8004
rect 24728 7964 24734 7976
rect 24810 7973 24822 7976
rect 24856 7973 24868 8007
rect 24810 7967 24868 7973
rect 26875 8007 26933 8013
rect 26875 7973 26887 8007
rect 26921 8004 26933 8007
rect 27338 8004 27344 8016
rect 26921 7976 27344 8004
rect 26921 7973 26933 7976
rect 26875 7967 26933 7973
rect 27338 7964 27344 7976
rect 27396 8004 27402 8016
rect 28810 8004 28816 8016
rect 27396 7976 28816 8004
rect 27396 7964 27402 7976
rect 28810 7964 28816 7976
rect 28868 8004 28874 8016
rect 29226 8007 29284 8013
rect 29226 8004 29238 8007
rect 28868 7976 29238 8004
rect 28868 7964 28874 7976
rect 29226 7973 29238 7976
rect 29272 7973 29284 8007
rect 29226 7967 29284 7973
rect 33867 8007 33925 8013
rect 33867 7973 33879 8007
rect 33913 8004 33925 8007
rect 34054 8004 34060 8016
rect 33913 7976 34060 8004
rect 33913 7973 33925 7976
rect 33867 7967 33925 7973
rect 34054 7964 34060 7976
rect 34112 7964 34118 8016
rect 35434 8004 35440 8016
rect 35347 7976 35440 8004
rect 35434 7964 35440 7976
rect 35492 7964 35498 8016
rect 23937 7939 23995 7945
rect 23937 7936 23949 7939
rect 23446 7908 23949 7936
rect 23201 7899 23259 7905
rect 23937 7905 23949 7908
rect 23983 7936 23995 7939
rect 24118 7936 24124 7948
rect 23983 7908 24124 7936
rect 23983 7905 23995 7908
rect 23937 7899 23995 7905
rect 24118 7896 24124 7908
rect 24176 7936 24182 7948
rect 27062 7936 27068 7948
rect 24176 7908 27068 7936
rect 24176 7896 24182 7908
rect 27062 7896 27068 7908
rect 27120 7896 27126 7948
rect 29825 7939 29883 7945
rect 29825 7905 29837 7939
rect 29871 7936 29883 7939
rect 30190 7936 30196 7948
rect 29871 7908 30196 7936
rect 29871 7905 29883 7908
rect 29825 7899 29883 7905
rect 30190 7896 30196 7908
rect 30248 7896 30254 7948
rect 32560 7939 32618 7945
rect 32560 7905 32572 7939
rect 32606 7936 32618 7939
rect 32674 7936 32680 7948
rect 32606 7908 32680 7936
rect 32606 7905 32618 7908
rect 32560 7899 32618 7905
rect 32674 7896 32680 7908
rect 32732 7936 32738 7948
rect 35158 7936 35164 7948
rect 32732 7908 35164 7936
rect 32732 7896 32738 7908
rect 35158 7896 35164 7908
rect 35216 7896 35222 7948
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7868 18291 7871
rect 18598 7868 18604 7880
rect 18279 7840 18604 7868
rect 18279 7837 18291 7840
rect 18233 7831 18291 7837
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 19518 7868 19524 7880
rect 19479 7840 19524 7868
rect 19518 7828 19524 7840
rect 19576 7868 19582 7880
rect 21269 7871 21327 7877
rect 21269 7868 21281 7871
rect 19576 7840 21281 7868
rect 19576 7828 19582 7840
rect 21269 7837 21281 7840
rect 21315 7868 21327 7871
rect 21545 7871 21603 7877
rect 21545 7868 21557 7871
rect 21315 7840 21557 7868
rect 21315 7837 21327 7840
rect 21269 7831 21327 7837
rect 21545 7837 21557 7840
rect 21591 7837 21603 7871
rect 21818 7868 21824 7880
rect 21779 7840 21824 7868
rect 21545 7831 21603 7837
rect 21818 7828 21824 7840
rect 21876 7828 21882 7880
rect 23569 7871 23627 7877
rect 23569 7837 23581 7871
rect 23615 7868 23627 7871
rect 24394 7868 24400 7880
rect 23615 7840 24400 7868
rect 23615 7837 23627 7840
rect 23569 7831 23627 7837
rect 24394 7828 24400 7840
rect 24452 7828 24458 7880
rect 24489 7871 24547 7877
rect 24489 7837 24501 7871
rect 24535 7868 24547 7871
rect 25038 7868 25044 7880
rect 24535 7840 25044 7868
rect 24535 7837 24547 7840
rect 24489 7831 24547 7837
rect 25038 7828 25044 7840
rect 25096 7828 25102 7880
rect 26513 7871 26571 7877
rect 26513 7837 26525 7871
rect 26559 7868 26571 7871
rect 26694 7868 26700 7880
rect 26559 7840 26700 7868
rect 26559 7837 26571 7840
rect 26513 7831 26571 7837
rect 26694 7828 26700 7840
rect 26752 7828 26758 7880
rect 28905 7871 28963 7877
rect 28905 7837 28917 7871
rect 28951 7868 28963 7871
rect 29454 7868 29460 7880
rect 28951 7840 29460 7868
rect 28951 7837 28963 7840
rect 28905 7831 28963 7837
rect 29454 7828 29460 7840
rect 29512 7828 29518 7880
rect 29638 7828 29644 7880
rect 29696 7868 29702 7880
rect 30098 7868 30104 7880
rect 29696 7840 30104 7868
rect 29696 7828 29702 7840
rect 30098 7828 30104 7840
rect 30156 7828 30162 7880
rect 33502 7868 33508 7880
rect 33463 7840 33508 7868
rect 33502 7828 33508 7840
rect 33560 7828 33566 7880
rect 35342 7868 35348 7880
rect 35303 7840 35348 7868
rect 35342 7828 35348 7840
rect 35400 7828 35406 7880
rect 35618 7868 35624 7880
rect 35579 7840 35624 7868
rect 35618 7828 35624 7840
rect 35676 7828 35682 7880
rect 16209 7803 16267 7809
rect 16209 7769 16221 7803
rect 16255 7800 16267 7803
rect 17862 7800 17868 7812
rect 16255 7772 17868 7800
rect 16255 7769 16267 7772
rect 16209 7763 16267 7769
rect 17862 7760 17868 7772
rect 17920 7760 17926 7812
rect 25682 7760 25688 7812
rect 25740 7800 25746 7812
rect 30469 7803 30527 7809
rect 30469 7800 30481 7803
rect 25740 7772 30481 7800
rect 25740 7760 25746 7772
rect 30469 7769 30481 7772
rect 30515 7800 30527 7803
rect 30558 7800 30564 7812
rect 30515 7772 30564 7800
rect 30515 7769 30527 7772
rect 30469 7763 30527 7769
rect 30558 7760 30564 7772
rect 30616 7760 30622 7812
rect 33318 7800 33324 7812
rect 33106 7772 33324 7800
rect 16577 7735 16635 7741
rect 16577 7732 16589 7735
rect 16132 7704 16589 7732
rect 16577 7701 16589 7704
rect 16623 7732 16635 7735
rect 16850 7732 16856 7744
rect 16623 7704 16856 7732
rect 16623 7701 16635 7704
rect 16577 7695 16635 7701
rect 16850 7692 16856 7704
rect 16908 7732 16914 7744
rect 20530 7732 20536 7744
rect 16908 7704 20536 7732
rect 16908 7692 16914 7704
rect 20530 7692 20536 7704
rect 20588 7692 20594 7744
rect 24210 7732 24216 7744
rect 24171 7704 24216 7732
rect 24210 7692 24216 7704
rect 24268 7692 24274 7744
rect 27430 7732 27436 7744
rect 27391 7704 27436 7732
rect 27430 7692 27436 7704
rect 27488 7692 27494 7744
rect 27706 7732 27712 7744
rect 27667 7704 27712 7732
rect 27706 7692 27712 7704
rect 27764 7692 27770 7744
rect 32631 7735 32689 7741
rect 32631 7701 32643 7735
rect 32677 7732 32689 7735
rect 33106 7732 33134 7772
rect 33318 7760 33324 7772
rect 33376 7760 33382 7812
rect 32677 7704 33134 7732
rect 33229 7735 33287 7741
rect 32677 7701 32689 7704
rect 32631 7695 32689 7701
rect 33229 7701 33241 7735
rect 33275 7732 33287 7735
rect 33410 7732 33416 7744
rect 33275 7704 33416 7732
rect 33275 7701 33287 7704
rect 33229 7695 33287 7701
rect 33410 7692 33416 7704
rect 33468 7692 33474 7744
rect 34882 7732 34888 7744
rect 34843 7704 34888 7732
rect 34882 7692 34888 7704
rect 34940 7692 34946 7744
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 3142 7528 3148 7540
rect 3103 7500 3148 7528
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 8757 7531 8815 7537
rect 8757 7528 8769 7531
rect 5408 7500 8769 7528
rect 5408 7488 5414 7500
rect 8757 7497 8769 7500
rect 8803 7497 8815 7531
rect 9582 7528 9588 7540
rect 9543 7500 9588 7528
rect 8757 7491 8815 7497
rect 9582 7488 9588 7500
rect 9640 7528 9646 7540
rect 10226 7528 10232 7540
rect 9640 7500 10232 7528
rect 9640 7488 9646 7500
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 11793 7531 11851 7537
rect 11793 7497 11805 7531
rect 11839 7528 11851 7531
rect 12158 7528 12164 7540
rect 11839 7500 12164 7528
rect 11839 7497 11851 7500
rect 11793 7491 11851 7497
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 14182 7528 14188 7540
rect 12268 7500 14188 7528
rect 5902 7420 5908 7472
rect 5960 7460 5966 7472
rect 10134 7460 10140 7472
rect 5960 7432 10140 7460
rect 5960 7420 5966 7432
rect 10134 7420 10140 7432
rect 10192 7420 10198 7472
rect 10778 7420 10784 7472
rect 10836 7460 10842 7472
rect 11241 7463 11299 7469
rect 11241 7460 11253 7463
rect 10836 7432 11253 7460
rect 10836 7420 10842 7432
rect 11241 7429 11253 7432
rect 11287 7460 11299 7463
rect 12268 7460 12296 7500
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 14550 7528 14556 7540
rect 14511 7500 14556 7528
rect 14550 7488 14556 7500
rect 14608 7488 14614 7540
rect 15289 7531 15347 7537
rect 15289 7497 15301 7531
rect 15335 7528 15347 7531
rect 15470 7528 15476 7540
rect 15335 7500 15476 7528
rect 15335 7497 15347 7500
rect 15289 7491 15347 7497
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 17589 7531 17647 7537
rect 17589 7497 17601 7531
rect 17635 7528 17647 7531
rect 17862 7528 17868 7540
rect 17635 7500 17868 7528
rect 17635 7497 17647 7500
rect 17589 7491 17647 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 19242 7488 19248 7540
rect 19300 7528 19306 7540
rect 19613 7531 19671 7537
rect 19613 7528 19625 7531
rect 19300 7500 19625 7528
rect 19300 7488 19306 7500
rect 19613 7497 19625 7500
rect 19659 7497 19671 7531
rect 19613 7491 19671 7497
rect 20073 7531 20131 7537
rect 20073 7497 20085 7531
rect 20119 7528 20131 7531
rect 20714 7528 20720 7540
rect 20119 7500 20720 7528
rect 20119 7497 20131 7500
rect 20073 7491 20131 7497
rect 16114 7460 16120 7472
rect 11287 7432 12296 7460
rect 13141 7432 16120 7460
rect 11287 7429 11299 7432
rect 11241 7423 11299 7429
rect 4062 7352 4068 7404
rect 4120 7392 4126 7404
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 4120 7364 4169 7392
rect 4120 7352 4126 7364
rect 4157 7361 4169 7364
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 5626 7352 5632 7404
rect 5684 7392 5690 7404
rect 5721 7395 5779 7401
rect 5721 7392 5733 7395
rect 5684 7364 5733 7392
rect 5684 7352 5690 7364
rect 5721 7361 5733 7364
rect 5767 7392 5779 7395
rect 8294 7392 8300 7404
rect 5767 7364 8300 7392
rect 5767 7361 5779 7364
rect 5721 7355 5779 7361
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 9858 7392 9864 7404
rect 9088 7364 9864 7392
rect 9088 7352 9094 7364
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 10226 7352 10232 7404
rect 10284 7392 10290 7404
rect 10284 7364 10329 7392
rect 10284 7352 10290 7364
rect 10410 7352 10416 7404
rect 10468 7392 10474 7404
rect 13141 7392 13169 7432
rect 10468 7364 13169 7392
rect 13633 7395 13691 7401
rect 10468 7352 10474 7364
rect 13633 7361 13645 7395
rect 13679 7392 13691 7395
rect 13814 7392 13820 7404
rect 13679 7364 13820 7392
rect 13679 7361 13691 7364
rect 13633 7355 13691 7361
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 13924 7401 13952 7432
rect 16114 7420 16120 7432
rect 16172 7420 16178 7472
rect 20088 7460 20116 7491
rect 20714 7488 20720 7500
rect 20772 7488 20778 7540
rect 21634 7488 21640 7540
rect 21692 7528 21698 7540
rect 22373 7531 22431 7537
rect 22373 7528 22385 7531
rect 21692 7500 22385 7528
rect 21692 7488 21698 7500
rect 22373 7497 22385 7500
rect 22419 7497 22431 7531
rect 22373 7491 22431 7497
rect 23474 7488 23480 7540
rect 23532 7528 23538 7540
rect 28902 7528 28908 7540
rect 23532 7500 28908 7528
rect 23532 7488 23538 7500
rect 18708 7432 20116 7460
rect 13909 7395 13967 7401
rect 13909 7361 13921 7395
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 16209 7395 16267 7401
rect 16209 7361 16221 7395
rect 16255 7392 16267 7395
rect 17034 7392 17040 7404
rect 16255 7364 17040 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 17034 7352 17040 7364
rect 17092 7352 17098 7404
rect 18708 7401 18736 7432
rect 18693 7395 18751 7401
rect 18693 7361 18705 7395
rect 18739 7361 18751 7395
rect 18693 7355 18751 7361
rect 19337 7395 19395 7401
rect 19337 7361 19349 7395
rect 19383 7392 19395 7395
rect 19518 7392 19524 7404
rect 19383 7364 19524 7392
rect 19383 7361 19395 7364
rect 19337 7355 19395 7361
rect 19518 7352 19524 7364
rect 19576 7352 19582 7404
rect 21453 7395 21511 7401
rect 21453 7361 21465 7395
rect 21499 7392 21511 7395
rect 21542 7392 21548 7404
rect 21499 7364 21548 7392
rect 21499 7361 21511 7364
rect 21453 7355 21511 7361
rect 21542 7352 21548 7364
rect 21600 7352 21606 7404
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7324 2283 7327
rect 3510 7324 3516 7336
rect 2271 7296 3516 7324
rect 2271 7293 2283 7296
rect 2225 7287 2283 7293
rect 3510 7284 3516 7296
rect 3568 7284 3574 7336
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7324 6699 7327
rect 6822 7324 6828 7336
rect 6687 7296 6828 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 7837 7327 7895 7333
rect 7837 7293 7849 7327
rect 7883 7324 7895 7327
rect 8018 7324 8024 7336
rect 7883 7296 8024 7324
rect 7883 7293 7895 7296
rect 7837 7287 7895 7293
rect 8018 7284 8024 7296
rect 8076 7284 8082 7336
rect 10042 7324 10048 7336
rect 10003 7296 10048 7324
rect 10042 7284 10048 7296
rect 10100 7284 10106 7336
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 10919 7296 10977 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 10965 7287 11023 7293
rect 12342 7284 12348 7336
rect 12400 7324 12406 7336
rect 12564 7327 12622 7333
rect 12564 7324 12576 7327
rect 12400 7296 12576 7324
rect 12400 7284 12406 7296
rect 12564 7293 12576 7296
rect 12610 7324 12622 7327
rect 12989 7327 13047 7333
rect 12989 7324 13001 7327
rect 12610 7296 13001 7324
rect 12610 7293 12622 7296
rect 12564 7287 12622 7293
rect 12989 7293 13001 7296
rect 13035 7293 13047 7327
rect 12989 7287 13047 7293
rect 15105 7327 15163 7333
rect 15105 7293 15117 7327
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 1857 7259 1915 7265
rect 1857 7225 1869 7259
rect 1903 7256 1915 7259
rect 2130 7256 2136 7268
rect 1903 7228 2136 7256
rect 1903 7225 1915 7228
rect 1857 7219 1915 7225
rect 2130 7216 2136 7228
rect 2188 7256 2194 7268
rect 2587 7259 2645 7265
rect 2587 7256 2599 7259
rect 2188 7228 2599 7256
rect 2188 7216 2194 7228
rect 2587 7225 2599 7228
rect 2633 7256 2645 7259
rect 3694 7256 3700 7268
rect 2633 7228 3700 7256
rect 2633 7225 2645 7228
rect 2587 7219 2645 7225
rect 3528 7197 3556 7228
rect 3694 7216 3700 7228
rect 3752 7256 3758 7268
rect 4065 7259 4123 7265
rect 4065 7256 4077 7259
rect 3752 7228 4077 7256
rect 3752 7216 3758 7228
rect 4065 7225 4077 7228
rect 4111 7256 4123 7259
rect 4519 7259 4577 7265
rect 4519 7256 4531 7259
rect 4111 7228 4531 7256
rect 4111 7225 4123 7228
rect 4065 7219 4123 7225
rect 4519 7225 4531 7228
rect 4565 7256 4577 7259
rect 7190 7256 7196 7268
rect 4565 7228 7196 7256
rect 4565 7225 4577 7228
rect 4519 7219 4577 7225
rect 7190 7216 7196 7228
rect 7248 7256 7254 7268
rect 7377 7259 7435 7265
rect 7377 7256 7389 7259
rect 7248 7228 7389 7256
rect 7248 7216 7254 7228
rect 7377 7225 7389 7228
rect 7423 7256 7435 7259
rect 7745 7259 7803 7265
rect 7745 7256 7757 7259
rect 7423 7228 7757 7256
rect 7423 7225 7435 7228
rect 7377 7219 7435 7225
rect 7745 7225 7757 7228
rect 7791 7256 7803 7259
rect 8110 7256 8116 7268
rect 7791 7228 8116 7256
rect 7791 7225 7803 7228
rect 7745 7219 7803 7225
rect 8110 7216 8116 7228
rect 8168 7265 8174 7268
rect 8168 7259 8216 7265
rect 8168 7225 8170 7259
rect 8204 7225 8216 7259
rect 8168 7219 8216 7225
rect 9309 7259 9367 7265
rect 9309 7225 9321 7259
rect 9355 7256 9367 7259
rect 10321 7259 10379 7265
rect 9355 7228 9674 7256
rect 9355 7225 9367 7228
rect 9309 7219 9367 7225
rect 8168 7216 8174 7219
rect 3513 7191 3571 7197
rect 3513 7157 3525 7191
rect 3559 7157 3571 7191
rect 5074 7188 5080 7200
rect 5035 7160 5080 7188
rect 3513 7151 3571 7157
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 6273 7191 6331 7197
rect 6273 7157 6285 7191
rect 6319 7188 6331 7191
rect 6914 7188 6920 7200
rect 6319 7160 6920 7188
rect 6319 7157 6331 7160
rect 6273 7151 6331 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7009 7191 7067 7197
rect 7009 7157 7021 7191
rect 7055 7188 7067 7191
rect 7098 7188 7104 7200
rect 7055 7160 7104 7188
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 9646 7188 9674 7228
rect 10321 7225 10333 7259
rect 10367 7225 10379 7259
rect 10321 7219 10379 7225
rect 10042 7188 10048 7200
rect 9646 7160 10048 7188
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10336 7188 10364 7219
rect 10410 7216 10416 7268
rect 10468 7256 10474 7268
rect 12434 7256 12440 7268
rect 10468 7228 12440 7256
rect 10468 7216 10474 7228
rect 12434 7216 12440 7228
rect 12492 7256 12498 7268
rect 13357 7259 13415 7265
rect 13357 7256 13369 7259
rect 12492 7228 13369 7256
rect 12492 7216 12498 7228
rect 13357 7225 13369 7228
rect 13403 7256 13415 7259
rect 13630 7256 13636 7268
rect 13403 7228 13636 7256
rect 13403 7225 13415 7228
rect 13357 7219 13415 7225
rect 13630 7216 13636 7228
rect 13688 7216 13694 7268
rect 13725 7259 13783 7265
rect 13725 7225 13737 7259
rect 13771 7256 13783 7259
rect 13998 7256 14004 7268
rect 13771 7228 14004 7256
rect 13771 7225 13783 7228
rect 13725 7219 13783 7225
rect 13998 7216 14004 7228
rect 14056 7216 14062 7268
rect 15013 7259 15071 7265
rect 15013 7225 15025 7259
rect 15059 7256 15071 7259
rect 15120 7256 15148 7287
rect 15286 7284 15292 7336
rect 15344 7324 15350 7336
rect 15657 7327 15715 7333
rect 15657 7324 15669 7327
rect 15344 7296 15669 7324
rect 15344 7284 15350 7296
rect 15657 7293 15669 7296
rect 15703 7324 15715 7327
rect 15746 7324 15752 7336
rect 15703 7296 15752 7324
rect 15703 7293 15715 7296
rect 15657 7287 15715 7293
rect 15746 7284 15752 7296
rect 15804 7324 15810 7336
rect 16117 7327 16175 7333
rect 16117 7324 16129 7327
rect 15804 7296 16129 7324
rect 15804 7284 15810 7296
rect 16117 7293 16129 7296
rect 16163 7324 16175 7327
rect 17129 7327 17187 7333
rect 16163 7296 16614 7324
rect 16163 7293 16175 7296
rect 16117 7287 16175 7293
rect 16206 7256 16212 7268
rect 15059 7228 16212 7256
rect 15059 7225 15071 7228
rect 15013 7219 15071 7225
rect 16206 7216 16212 7228
rect 16264 7216 16270 7268
rect 16586 7265 16614 7296
rect 17129 7293 17141 7327
rect 17175 7324 17187 7327
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 17175 7296 18429 7324
rect 17175 7293 17187 7296
rect 17129 7287 17187 7293
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 18417 7287 18475 7293
rect 20216 7327 20274 7333
rect 20216 7293 20228 7327
rect 20262 7324 20274 7327
rect 20622 7324 20628 7336
rect 20262 7296 20628 7324
rect 20262 7293 20274 7296
rect 20216 7287 20274 7293
rect 16571 7259 16629 7265
rect 16571 7225 16583 7259
rect 16617 7256 16629 7259
rect 16666 7256 16672 7268
rect 16617 7228 16672 7256
rect 16617 7225 16629 7228
rect 16571 7219 16629 7225
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 10962 7188 10968 7200
rect 10192 7160 10364 7188
rect 10923 7160 10968 7188
rect 10192 7148 10198 7160
rect 10962 7148 10968 7160
rect 11020 7148 11026 7200
rect 12158 7188 12164 7200
rect 12119 7160 12164 7188
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 12667 7191 12725 7197
rect 12667 7157 12679 7191
rect 12713 7188 12725 7191
rect 12894 7188 12900 7200
rect 12713 7160 12900 7188
rect 12713 7157 12725 7160
rect 12667 7151 12725 7157
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 18432 7188 18460 7287
rect 20622 7284 20628 7296
rect 20680 7324 20686 7336
rect 22830 7324 22836 7336
rect 20680 7296 22836 7324
rect 20680 7284 20686 7296
rect 22830 7284 22836 7296
rect 22888 7284 22894 7336
rect 23952 7333 23980 7500
rect 28902 7488 28908 7500
rect 28960 7488 28966 7540
rect 32674 7528 32680 7540
rect 32635 7500 32680 7528
rect 32674 7488 32680 7500
rect 32732 7488 32738 7540
rect 34054 7488 34060 7540
rect 34112 7528 34118 7540
rect 34241 7531 34299 7537
rect 34241 7528 34253 7531
rect 34112 7500 34253 7528
rect 34112 7488 34118 7500
rect 34241 7497 34253 7500
rect 34287 7497 34299 7531
rect 34241 7491 34299 7497
rect 35434 7488 35440 7540
rect 35492 7528 35498 7540
rect 35897 7531 35955 7537
rect 35897 7528 35909 7531
rect 35492 7500 35909 7528
rect 35492 7488 35498 7500
rect 35897 7497 35909 7500
rect 35943 7497 35955 7531
rect 36630 7528 36636 7540
rect 36591 7500 36636 7528
rect 35897 7491 35955 7497
rect 36630 7488 36636 7500
rect 36688 7488 36694 7540
rect 26970 7420 26976 7472
rect 27028 7460 27034 7472
rect 27522 7460 27528 7472
rect 27028 7432 27528 7460
rect 27028 7420 27034 7432
rect 27522 7420 27528 7432
rect 27580 7460 27586 7472
rect 28261 7463 28319 7469
rect 28261 7460 28273 7463
rect 27580 7432 28273 7460
rect 27580 7420 27586 7432
rect 28261 7429 28273 7432
rect 28307 7429 28319 7463
rect 28261 7423 28319 7429
rect 32355 7463 32413 7469
rect 32355 7429 32367 7463
rect 32401 7460 32413 7463
rect 34882 7460 34888 7472
rect 32401 7432 34888 7460
rect 32401 7429 32413 7432
rect 32355 7423 32413 7429
rect 34882 7420 34888 7432
rect 34940 7460 34946 7472
rect 34940 7432 35020 7460
rect 34940 7420 34946 7432
rect 24210 7392 24216 7404
rect 24171 7364 24216 7392
rect 24210 7352 24216 7364
rect 24268 7352 24274 7404
rect 25869 7395 25927 7401
rect 25869 7361 25881 7395
rect 25915 7392 25927 7395
rect 26142 7392 26148 7404
rect 25915 7364 26148 7392
rect 25915 7361 25927 7364
rect 25869 7355 25927 7361
rect 26142 7352 26148 7364
rect 26200 7352 26206 7404
rect 27706 7392 27712 7404
rect 27667 7364 27712 7392
rect 27706 7352 27712 7364
rect 27764 7392 27770 7404
rect 27982 7392 27988 7404
rect 27764 7364 27988 7392
rect 27764 7352 27770 7364
rect 27982 7352 27988 7364
rect 28040 7352 28046 7404
rect 28810 7352 28816 7404
rect 28868 7392 28874 7404
rect 28905 7395 28963 7401
rect 28905 7392 28917 7395
rect 28868 7364 28917 7392
rect 28868 7352 28874 7364
rect 28905 7361 28917 7364
rect 28951 7392 28963 7395
rect 29917 7395 29975 7401
rect 29917 7392 29929 7395
rect 28951 7364 29929 7392
rect 28951 7361 28963 7364
rect 28905 7355 28963 7361
rect 29917 7361 29929 7364
rect 29963 7361 29975 7395
rect 30098 7392 30104 7404
rect 30059 7364 30104 7392
rect 29917 7355 29975 7361
rect 23937 7327 23995 7333
rect 23937 7293 23949 7327
rect 23983 7293 23995 7327
rect 24118 7324 24124 7336
rect 24079 7296 24124 7324
rect 23937 7287 23995 7293
rect 24118 7284 24124 7296
rect 24176 7284 24182 7336
rect 26789 7327 26847 7333
rect 26789 7293 26801 7327
rect 26835 7324 26847 7327
rect 27433 7327 27491 7333
rect 27433 7324 27445 7327
rect 26835 7296 27445 7324
rect 26835 7293 26847 7296
rect 26789 7287 26847 7293
rect 27433 7293 27445 7296
rect 27479 7293 27491 7327
rect 27433 7287 27491 7293
rect 18785 7259 18843 7265
rect 18785 7225 18797 7259
rect 18831 7225 18843 7259
rect 18785 7219 18843 7225
rect 18598 7188 18604 7200
rect 18432 7160 18604 7188
rect 18598 7148 18604 7160
rect 18656 7188 18662 7200
rect 18800 7188 18828 7219
rect 19426 7216 19432 7268
rect 19484 7256 19490 7268
rect 20303 7259 20361 7265
rect 20303 7256 20315 7259
rect 19484 7228 20315 7256
rect 19484 7216 19490 7228
rect 20303 7225 20315 7228
rect 20349 7225 20361 7259
rect 21358 7256 21364 7268
rect 21271 7228 21364 7256
rect 20303 7219 20361 7225
rect 21358 7216 21364 7228
rect 21416 7256 21422 7268
rect 21815 7259 21873 7265
rect 21815 7256 21827 7259
rect 21416 7228 21827 7256
rect 21416 7216 21422 7228
rect 21815 7225 21827 7228
rect 21861 7256 21873 7259
rect 25685 7259 25743 7265
rect 25685 7256 25697 7259
rect 21861 7228 25697 7256
rect 21861 7225 21873 7228
rect 21815 7219 21873 7225
rect 24688 7200 24716 7228
rect 25685 7225 25697 7228
rect 25731 7256 25743 7259
rect 26190 7259 26248 7265
rect 26190 7256 26202 7259
rect 25731 7228 26202 7256
rect 25731 7225 25743 7228
rect 25685 7219 25743 7225
rect 26190 7225 26202 7228
rect 26236 7256 26248 7259
rect 27065 7259 27123 7265
rect 27065 7256 27077 7259
rect 26236 7228 27077 7256
rect 26236 7225 26248 7228
rect 26190 7219 26248 7225
rect 27065 7225 27077 7228
rect 27111 7256 27123 7259
rect 27338 7256 27344 7268
rect 27111 7228 27344 7256
rect 27111 7225 27123 7228
rect 27065 7219 27123 7225
rect 27338 7216 27344 7228
rect 27396 7216 27402 7268
rect 18656 7160 18828 7188
rect 18656 7148 18662 7160
rect 22002 7148 22008 7200
rect 22060 7188 22066 7200
rect 22646 7188 22652 7200
rect 22060 7160 22652 7188
rect 22060 7148 22066 7160
rect 22646 7148 22652 7160
rect 22704 7148 22710 7200
rect 23014 7188 23020 7200
rect 22975 7160 23020 7188
rect 23014 7148 23020 7160
rect 23072 7148 23078 7200
rect 24670 7188 24676 7200
rect 24631 7160 24676 7188
rect 24670 7148 24676 7160
rect 24728 7148 24734 7200
rect 25038 7188 25044 7200
rect 24999 7160 25044 7188
rect 25038 7148 25044 7160
rect 25096 7148 25102 7200
rect 27448 7188 27476 7287
rect 27801 7259 27859 7265
rect 27801 7225 27813 7259
rect 27847 7225 27859 7259
rect 29932 7256 29960 7355
rect 30098 7352 30104 7364
rect 30156 7352 30162 7404
rect 33410 7392 33416 7404
rect 33106 7364 33416 7392
rect 31754 7284 31760 7336
rect 31812 7324 31818 7336
rect 32252 7327 32310 7333
rect 32252 7324 32264 7327
rect 31812 7296 32264 7324
rect 31812 7284 31818 7296
rect 32252 7293 32264 7296
rect 32298 7324 32310 7327
rect 32493 7327 32551 7333
rect 32493 7324 32505 7327
rect 32298 7296 32505 7324
rect 32298 7293 32310 7296
rect 32252 7287 32310 7293
rect 32493 7293 32505 7296
rect 32539 7293 32551 7327
rect 32493 7287 32551 7293
rect 30422 7259 30480 7265
rect 30422 7256 30434 7259
rect 29932 7228 30434 7256
rect 27801 7219 27859 7225
rect 30422 7225 30434 7228
rect 30468 7256 30480 7259
rect 32030 7256 32036 7268
rect 30468 7228 32036 7256
rect 30468 7225 30480 7228
rect 30422 7219 30480 7225
rect 27816 7188 27844 7219
rect 32030 7216 32036 7228
rect 32088 7216 32094 7268
rect 33106 7256 33134 7364
rect 33410 7352 33416 7364
rect 33468 7392 33474 7404
rect 34992 7401 35020 7432
rect 34609 7395 34667 7401
rect 34609 7392 34621 7395
rect 33468 7364 34621 7392
rect 33468 7352 33474 7364
rect 34609 7361 34621 7364
rect 34655 7361 34667 7395
rect 34609 7355 34667 7361
rect 34977 7395 35035 7401
rect 34977 7361 34989 7395
rect 35023 7361 35035 7395
rect 35342 7392 35348 7404
rect 35303 7364 35348 7392
rect 34977 7355 35035 7361
rect 33318 7256 33324 7268
rect 32278 7228 33134 7256
rect 33279 7228 33324 7256
rect 29454 7188 29460 7200
rect 27448 7160 27844 7188
rect 29415 7160 29460 7188
rect 29454 7148 29460 7160
rect 29512 7148 29518 7200
rect 31021 7191 31079 7197
rect 31021 7157 31033 7191
rect 31067 7188 31079 7191
rect 32278 7188 32306 7228
rect 33318 7216 33324 7228
rect 33376 7216 33382 7268
rect 33410 7216 33416 7268
rect 33468 7256 33474 7268
rect 33965 7259 34023 7265
rect 33468 7228 33513 7256
rect 33468 7216 33474 7228
rect 33965 7225 33977 7259
rect 34011 7256 34023 7259
rect 34624 7256 34652 7355
rect 35342 7352 35348 7364
rect 35400 7352 35406 7404
rect 36449 7327 36507 7333
rect 36449 7293 36461 7327
rect 36495 7293 36507 7327
rect 36449 7287 36507 7293
rect 35069 7259 35127 7265
rect 35069 7256 35081 7259
rect 34011 7228 34376 7256
rect 34624 7228 35081 7256
rect 34011 7225 34023 7228
rect 33965 7219 34023 7225
rect 31067 7160 32306 7188
rect 32493 7191 32551 7197
rect 31067 7157 31079 7160
rect 31021 7151 31079 7157
rect 32493 7157 32505 7191
rect 32539 7188 32551 7191
rect 33137 7191 33195 7197
rect 33137 7188 33149 7191
rect 32539 7160 33149 7188
rect 32539 7157 32551 7160
rect 32493 7151 32551 7157
rect 33137 7157 33149 7160
rect 33183 7188 33195 7191
rect 34054 7188 34060 7200
rect 33183 7160 34060 7188
rect 33183 7157 33195 7160
rect 33137 7151 33195 7157
rect 34054 7148 34060 7160
rect 34112 7148 34118 7200
rect 34348 7188 34376 7228
rect 35069 7225 35081 7228
rect 35115 7225 35127 7259
rect 35069 7219 35127 7225
rect 35158 7216 35164 7268
rect 35216 7256 35222 7268
rect 36464 7256 36492 7287
rect 37001 7259 37059 7265
rect 37001 7256 37013 7259
rect 35216 7228 37013 7256
rect 35216 7216 35222 7228
rect 37001 7225 37013 7228
rect 37047 7225 37059 7259
rect 37001 7219 37059 7225
rect 34974 7188 34980 7200
rect 34348 7160 34980 7188
rect 34974 7148 34980 7160
rect 35032 7188 35038 7200
rect 36354 7188 36360 7200
rect 35032 7160 36360 7188
rect 35032 7148 35038 7160
rect 36354 7148 36360 7160
rect 36412 7148 36418 7200
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 1762 6984 1768 6996
rect 1723 6956 1768 6984
rect 1762 6944 1768 6956
rect 1820 6944 1826 6996
rect 2866 6944 2872 6996
rect 2924 6984 2930 6996
rect 3421 6987 3479 6993
rect 3421 6984 3433 6987
rect 2924 6956 3433 6984
rect 2924 6944 2930 6956
rect 3421 6953 3433 6956
rect 3467 6953 3479 6987
rect 3421 6947 3479 6953
rect 8757 6987 8815 6993
rect 8757 6953 8769 6987
rect 8803 6984 8815 6987
rect 10410 6984 10416 6996
rect 8803 6956 10416 6984
rect 8803 6953 8815 6956
rect 8757 6947 8815 6953
rect 10410 6944 10416 6956
rect 10468 6944 10474 6996
rect 13998 6984 14004 6996
rect 13959 6956 14004 6984
rect 13998 6944 14004 6956
rect 14056 6944 14062 6996
rect 14182 6944 14188 6996
rect 14240 6984 14246 6996
rect 14369 6987 14427 6993
rect 14369 6984 14381 6987
rect 14240 6956 14381 6984
rect 14240 6944 14246 6956
rect 14369 6953 14381 6956
rect 14415 6953 14427 6987
rect 14369 6947 14427 6953
rect 17497 6987 17555 6993
rect 17497 6953 17509 6987
rect 17543 6984 17555 6987
rect 17586 6984 17592 6996
rect 17543 6956 17592 6984
rect 17543 6953 17555 6956
rect 17497 6947 17555 6953
rect 17586 6944 17592 6956
rect 17644 6944 17650 6996
rect 18506 6984 18512 6996
rect 18419 6956 18512 6984
rect 18506 6944 18512 6956
rect 18564 6984 18570 6996
rect 19426 6984 19432 6996
rect 18564 6956 19432 6984
rect 18564 6944 18570 6956
rect 19426 6944 19432 6956
rect 19484 6944 19490 6996
rect 19889 6987 19947 6993
rect 19889 6953 19901 6987
rect 19935 6984 19947 6987
rect 19935 6956 21128 6984
rect 19935 6953 19947 6956
rect 19889 6947 19947 6953
rect 2130 6876 2136 6928
rect 2188 6916 2194 6928
rect 2546 6919 2604 6925
rect 2546 6916 2558 6919
rect 2188 6888 2558 6916
rect 2188 6876 2194 6888
rect 2546 6885 2558 6888
rect 2592 6885 2604 6919
rect 2546 6879 2604 6885
rect 3881 6919 3939 6925
rect 3881 6885 3893 6919
rect 3927 6916 3939 6919
rect 4154 6916 4160 6928
rect 3927 6888 4160 6916
rect 3927 6885 3939 6888
rect 3881 6879 3939 6885
rect 4154 6876 4160 6888
rect 4212 6916 4218 6928
rect 4525 6919 4583 6925
rect 4525 6916 4537 6919
rect 4212 6888 4537 6916
rect 4212 6876 4218 6888
rect 4525 6885 4537 6888
rect 4571 6916 4583 6919
rect 5074 6916 5080 6928
rect 4571 6888 5080 6916
rect 4571 6885 4583 6888
rect 4525 6879 4583 6885
rect 5074 6876 5080 6888
rect 5132 6876 5138 6928
rect 6911 6919 6969 6925
rect 6911 6885 6923 6919
rect 6957 6916 6969 6919
rect 7190 6916 7196 6928
rect 6957 6888 7196 6916
rect 6957 6885 6969 6888
rect 6911 6879 6969 6885
rect 7190 6876 7196 6888
rect 7248 6876 7254 6928
rect 9766 6876 9772 6928
rect 9824 6916 9830 6928
rect 9998 6919 10056 6925
rect 9998 6916 10010 6919
rect 9824 6888 10010 6916
rect 9824 6876 9830 6888
rect 9998 6885 10010 6888
rect 10044 6885 10056 6919
rect 9998 6879 10056 6885
rect 12158 6876 12164 6928
rect 12216 6916 12222 6928
rect 12298 6919 12356 6925
rect 12298 6916 12310 6919
rect 12216 6888 12310 6916
rect 12216 6876 12222 6888
rect 12298 6885 12310 6888
rect 12344 6885 12356 6919
rect 12298 6879 12356 6885
rect 13725 6919 13783 6925
rect 13725 6885 13737 6919
rect 13771 6916 13783 6919
rect 14090 6916 14096 6928
rect 13771 6888 14096 6916
rect 13771 6885 13783 6888
rect 13725 6879 13783 6885
rect 14090 6876 14096 6888
rect 14148 6876 14154 6928
rect 15841 6919 15899 6925
rect 15841 6885 15853 6919
rect 15887 6916 15899 6919
rect 16117 6919 16175 6925
rect 16117 6916 16129 6919
rect 15887 6888 16129 6916
rect 15887 6885 15899 6888
rect 15841 6879 15899 6885
rect 16117 6885 16129 6888
rect 16163 6916 16175 6919
rect 16298 6916 16304 6928
rect 16163 6888 16304 6916
rect 16163 6885 16175 6888
rect 16117 6879 16175 6885
rect 16298 6876 16304 6888
rect 16356 6876 16362 6928
rect 16666 6876 16672 6928
rect 16724 6916 16730 6928
rect 19222 6919 19280 6925
rect 19222 6916 19234 6919
rect 16724 6888 19234 6916
rect 16724 6876 16730 6888
rect 19222 6885 19234 6888
rect 19268 6916 19280 6919
rect 19334 6916 19340 6928
rect 19268 6888 19340 6916
rect 19268 6885 19280 6888
rect 19222 6879 19280 6885
rect 19334 6876 19340 6888
rect 19392 6876 19398 6928
rect 21100 6925 21128 6956
rect 21542 6944 21548 6996
rect 21600 6944 21606 6996
rect 21634 6944 21640 6996
rect 21692 6984 21698 6996
rect 21913 6987 21971 6993
rect 21913 6984 21925 6987
rect 21692 6956 21925 6984
rect 21692 6944 21698 6956
rect 21913 6953 21925 6956
rect 21959 6953 21971 6987
rect 25961 6987 26019 6993
rect 21913 6947 21971 6953
rect 24044 6956 25176 6984
rect 20993 6919 21051 6925
rect 20993 6916 21005 6919
rect 20640 6888 21005 6916
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 6730 6848 6736 6860
rect 6595 6820 6736 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 6730 6808 6736 6820
rect 6788 6808 6794 6860
rect 8570 6848 8576 6860
rect 8531 6820 8576 6848
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 10134 6808 10140 6860
rect 10192 6848 10198 6860
rect 10597 6851 10655 6857
rect 10597 6848 10609 6851
rect 10192 6820 10609 6848
rect 10192 6808 10198 6820
rect 10597 6817 10609 6820
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 14185 6851 14243 6857
rect 14185 6817 14197 6851
rect 14231 6848 14243 6851
rect 14734 6848 14740 6860
rect 14231 6820 14740 6848
rect 14231 6817 14243 6820
rect 14185 6811 14243 6817
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 17586 6848 17592 6860
rect 17547 6820 17592 6848
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 17770 6848 17776 6860
rect 17731 6820 17776 6848
rect 17770 6808 17776 6820
rect 17828 6808 17834 6860
rect 18690 6808 18696 6860
rect 18748 6848 18754 6860
rect 20640 6857 20668 6888
rect 20993 6885 21005 6888
rect 21039 6885 21051 6919
rect 20993 6879 21051 6885
rect 21085 6919 21143 6925
rect 21085 6885 21097 6919
rect 21131 6916 21143 6919
rect 21266 6916 21272 6928
rect 21131 6888 21272 6916
rect 21131 6885 21143 6888
rect 21085 6879 21143 6885
rect 21266 6876 21272 6888
rect 21324 6876 21330 6928
rect 21560 6916 21588 6944
rect 22281 6919 22339 6925
rect 22281 6916 22293 6919
rect 21560 6888 22293 6916
rect 22281 6885 22293 6888
rect 22327 6885 22339 6919
rect 22281 6879 22339 6885
rect 20625 6851 20683 6857
rect 20625 6848 20637 6851
rect 18748 6820 20637 6848
rect 18748 6808 18754 6820
rect 20625 6817 20637 6820
rect 20671 6817 20683 6851
rect 20625 6811 20683 6817
rect 21637 6851 21695 6857
rect 21637 6817 21649 6851
rect 21683 6848 21695 6851
rect 21818 6848 21824 6860
rect 21683 6820 21824 6848
rect 21683 6817 21695 6820
rect 21637 6811 21695 6817
rect 21818 6808 21824 6820
rect 21876 6848 21882 6860
rect 22462 6848 22468 6860
rect 22520 6857 22526 6860
rect 22520 6851 22558 6857
rect 21876 6820 22468 6848
rect 21876 6808 21882 6820
rect 22462 6808 22468 6820
rect 22546 6817 22558 6851
rect 22520 6811 22558 6817
rect 22520 6808 22526 6811
rect 23106 6808 23112 6860
rect 23164 6848 23170 6860
rect 24044 6857 24072 6956
rect 24489 6919 24547 6925
rect 24489 6885 24501 6919
rect 24535 6916 24547 6919
rect 25038 6916 25044 6928
rect 24535 6888 25044 6916
rect 24535 6885 24547 6888
rect 24489 6879 24547 6885
rect 25038 6876 25044 6888
rect 25096 6876 25102 6928
rect 25148 6916 25176 6956
rect 25961 6953 25973 6987
rect 26007 6984 26019 6987
rect 26142 6984 26148 6996
rect 26007 6956 26148 6984
rect 26007 6953 26019 6956
rect 25961 6947 26019 6953
rect 26142 6944 26148 6956
rect 26200 6944 26206 6996
rect 28258 6984 28264 6996
rect 26528 6956 28264 6984
rect 26528 6916 26556 6956
rect 28258 6944 28264 6956
rect 28316 6944 28322 6996
rect 30282 6984 30288 6996
rect 30243 6956 30288 6984
rect 30282 6944 30288 6956
rect 30340 6944 30346 6996
rect 33318 6944 33324 6996
rect 33376 6984 33382 6996
rect 33873 6987 33931 6993
rect 33873 6984 33885 6987
rect 33376 6956 33885 6984
rect 33376 6944 33382 6956
rect 33873 6953 33885 6956
rect 33919 6953 33931 6987
rect 35342 6984 35348 6996
rect 33873 6947 33931 6953
rect 35176 6956 35348 6984
rect 25148 6888 26556 6916
rect 27249 6919 27307 6925
rect 27249 6885 27261 6919
rect 27295 6916 27307 6919
rect 27430 6916 27436 6928
rect 27295 6888 27436 6916
rect 27295 6885 27307 6888
rect 27249 6879 27307 6885
rect 27430 6876 27436 6888
rect 27488 6876 27494 6928
rect 28810 6916 28816 6928
rect 28771 6888 28816 6916
rect 28810 6876 28816 6888
rect 28868 6876 28874 6928
rect 30300 6916 30328 6944
rect 30300 6888 30972 6916
rect 24029 6851 24087 6857
rect 24029 6848 24041 6851
rect 23164 6820 24041 6848
rect 23164 6808 23170 6820
rect 24029 6817 24041 6820
rect 24075 6817 24087 6851
rect 24029 6811 24087 6817
rect 24305 6851 24363 6857
rect 24305 6817 24317 6851
rect 24351 6817 24363 6851
rect 24305 6811 24363 6817
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 3234 6780 3240 6792
rect 2271 6752 3240 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 4430 6780 4436 6792
rect 3936 6752 4436 6780
rect 3936 6740 3942 6752
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 5442 6780 5448 6792
rect 4755 6752 5448 6780
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 3050 6672 3056 6724
rect 3108 6712 3114 6724
rect 4724 6712 4752 6743
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 9674 6780 9680 6792
rect 9635 6752 9680 6780
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 11974 6780 11980 6792
rect 11935 6752 11980 6780
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 14826 6740 14832 6792
rect 14884 6780 14890 6792
rect 16022 6780 16028 6792
rect 14884 6752 16028 6780
rect 14884 6740 14890 6752
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 16114 6740 16120 6792
rect 16172 6780 16178 6792
rect 16301 6783 16359 6789
rect 16301 6780 16313 6783
rect 16172 6752 16313 6780
rect 16172 6740 16178 6752
rect 16301 6749 16313 6752
rect 16347 6749 16359 6783
rect 16301 6743 16359 6749
rect 18141 6783 18199 6789
rect 18141 6749 18153 6783
rect 18187 6780 18199 6783
rect 18874 6780 18880 6792
rect 18187 6752 18880 6780
rect 18187 6749 18199 6752
rect 18141 6743 18199 6749
rect 18874 6740 18880 6752
rect 18932 6740 18938 6792
rect 18969 6783 19027 6789
rect 18969 6749 18981 6783
rect 19015 6749 19027 6783
rect 24320 6780 24348 6811
rect 24394 6808 24400 6860
rect 24452 6848 24458 6860
rect 25314 6848 25320 6860
rect 24452 6820 25320 6848
rect 24452 6808 24458 6820
rect 25314 6808 25320 6820
rect 25372 6808 25378 6860
rect 30466 6848 30472 6860
rect 30427 6820 30472 6848
rect 30466 6808 30472 6820
rect 30524 6808 30530 6860
rect 30944 6857 30972 6888
rect 32030 6876 32036 6928
rect 32088 6916 32094 6928
rect 32446 6919 32504 6925
rect 32446 6916 32458 6919
rect 32088 6888 32458 6916
rect 32088 6876 32094 6888
rect 32446 6885 32458 6888
rect 32492 6885 32504 6919
rect 34606 6916 34612 6928
rect 34567 6888 34612 6916
rect 32446 6879 32504 6885
rect 34606 6876 34612 6888
rect 34664 6876 34670 6928
rect 35176 6925 35204 6956
rect 35342 6944 35348 6956
rect 35400 6984 35406 6996
rect 35437 6987 35495 6993
rect 35437 6984 35449 6987
rect 35400 6956 35449 6984
rect 35400 6944 35406 6956
rect 35437 6953 35449 6956
rect 35483 6953 35495 6987
rect 35437 6947 35495 6953
rect 35161 6919 35219 6925
rect 35161 6885 35173 6919
rect 35207 6885 35219 6919
rect 36170 6916 36176 6928
rect 36131 6888 36176 6916
rect 35161 6879 35219 6885
rect 36170 6876 36176 6888
rect 36228 6876 36234 6928
rect 30929 6851 30987 6857
rect 30929 6817 30941 6851
rect 30975 6848 30987 6851
rect 31110 6848 31116 6860
rect 30975 6820 31116 6848
rect 30975 6817 30987 6820
rect 30929 6811 30987 6817
rect 31110 6808 31116 6820
rect 31168 6808 31174 6860
rect 24320 6752 24992 6780
rect 18969 6743 19027 6749
rect 3108 6684 4752 6712
rect 3108 6672 3114 6684
rect 18984 6656 19012 6743
rect 24964 6724 24992 6752
rect 26326 6740 26332 6792
rect 26384 6780 26390 6792
rect 27157 6783 27215 6789
rect 27157 6780 27169 6783
rect 26384 6752 27169 6780
rect 26384 6740 26390 6752
rect 27157 6749 27169 6752
rect 27203 6749 27215 6783
rect 27522 6780 27528 6792
rect 27483 6752 27528 6780
rect 27157 6743 27215 6749
rect 27522 6740 27528 6752
rect 27580 6740 27586 6792
rect 28537 6783 28595 6789
rect 28537 6749 28549 6783
rect 28583 6780 28595 6783
rect 28718 6780 28724 6792
rect 28583 6752 28724 6780
rect 28583 6749 28595 6752
rect 28537 6743 28595 6749
rect 28718 6740 28724 6752
rect 28776 6740 28782 6792
rect 29365 6783 29423 6789
rect 29365 6749 29377 6783
rect 29411 6780 29423 6783
rect 29638 6780 29644 6792
rect 29411 6752 29644 6780
rect 29411 6749 29423 6752
rect 29365 6743 29423 6749
rect 29638 6740 29644 6752
rect 29696 6740 29702 6792
rect 31205 6783 31263 6789
rect 31205 6749 31217 6783
rect 31251 6780 31263 6783
rect 32125 6783 32183 6789
rect 32125 6780 32137 6783
rect 31251 6752 32137 6780
rect 31251 6749 31263 6752
rect 31205 6743 31263 6749
rect 32125 6749 32137 6752
rect 32171 6780 32183 6783
rect 33870 6780 33876 6792
rect 32171 6752 33876 6780
rect 32171 6749 32183 6752
rect 32125 6743 32183 6749
rect 33870 6740 33876 6752
rect 33928 6740 33934 6792
rect 34146 6740 34152 6792
rect 34204 6780 34210 6792
rect 34517 6783 34575 6789
rect 34517 6780 34529 6783
rect 34204 6752 34529 6780
rect 34204 6740 34210 6752
rect 34517 6749 34529 6752
rect 34563 6749 34575 6783
rect 36078 6780 36084 6792
rect 36039 6752 36084 6780
rect 34517 6743 34575 6749
rect 36078 6740 36084 6752
rect 36136 6740 36142 6792
rect 36354 6780 36360 6792
rect 36315 6752 36360 6780
rect 36354 6740 36360 6752
rect 36412 6740 36418 6792
rect 24946 6672 24952 6724
rect 25004 6712 25010 6724
rect 25501 6715 25559 6721
rect 25501 6712 25513 6715
rect 25004 6684 25513 6712
rect 25004 6672 25010 6684
rect 25501 6681 25513 6684
rect 25547 6712 25559 6715
rect 26234 6712 26240 6724
rect 25547 6684 26240 6712
rect 25547 6681 25559 6684
rect 25501 6675 25559 6681
rect 26234 6672 26240 6684
rect 26292 6672 26298 6724
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 3145 6647 3203 6653
rect 3145 6644 3157 6647
rect 3016 6616 3157 6644
rect 3016 6604 3022 6616
rect 3145 6613 3157 6616
rect 3191 6613 3203 6647
rect 3145 6607 3203 6613
rect 7006 6604 7012 6656
rect 7064 6644 7070 6656
rect 7469 6647 7527 6653
rect 7469 6644 7481 6647
rect 7064 6616 7481 6644
rect 7064 6604 7070 6616
rect 7469 6613 7481 6616
rect 7515 6613 7527 6647
rect 7469 6607 7527 6613
rect 7929 6647 7987 6653
rect 7929 6613 7941 6647
rect 7975 6644 7987 6647
rect 8018 6644 8024 6656
rect 7975 6616 8024 6644
rect 7975 6613 7987 6616
rect 7929 6607 7987 6613
rect 8018 6604 8024 6616
rect 8076 6644 8082 6656
rect 8478 6644 8484 6656
rect 8076 6616 8484 6644
rect 8076 6604 8082 6616
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 9030 6644 9036 6656
rect 8991 6616 9036 6644
rect 9030 6604 9036 6616
rect 9088 6604 9094 6656
rect 10870 6604 10876 6656
rect 10928 6644 10934 6656
rect 12897 6647 12955 6653
rect 12897 6644 12909 6647
rect 10928 6616 12909 6644
rect 10928 6604 10934 6616
rect 12897 6613 12909 6616
rect 12943 6613 12955 6647
rect 16942 6644 16948 6656
rect 16903 6616 16948 6644
rect 12897 6607 12955 6613
rect 16942 6604 16948 6616
rect 17000 6604 17006 6656
rect 18877 6647 18935 6653
rect 18877 6613 18889 6647
rect 18923 6644 18935 6647
rect 18966 6644 18972 6656
rect 18923 6616 18972 6644
rect 18923 6613 18935 6616
rect 18877 6607 18935 6613
rect 18966 6604 18972 6616
rect 19024 6604 19030 6656
rect 22603 6647 22661 6653
rect 22603 6613 22615 6647
rect 22649 6644 22661 6647
rect 25406 6644 25412 6656
rect 22649 6616 25412 6644
rect 22649 6613 22661 6616
rect 22603 6607 22661 6613
rect 25406 6604 25412 6616
rect 25464 6604 25470 6656
rect 26694 6644 26700 6656
rect 26655 6616 26700 6644
rect 26694 6604 26700 6616
rect 26752 6604 26758 6656
rect 33042 6644 33048 6656
rect 33003 6616 33048 6644
rect 33042 6604 33048 6616
rect 33100 6604 33106 6656
rect 33318 6604 33324 6656
rect 33376 6644 33382 6656
rect 33502 6644 33508 6656
rect 33376 6616 33508 6644
rect 33376 6604 33382 6616
rect 33502 6604 33508 6616
rect 33560 6604 33566 6656
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 2130 6400 2136 6452
rect 2188 6440 2194 6452
rect 2317 6443 2375 6449
rect 2317 6440 2329 6443
rect 2188 6412 2329 6440
rect 2188 6400 2194 6412
rect 2317 6409 2329 6412
rect 2363 6409 2375 6443
rect 2317 6403 2375 6409
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4212 6412 4257 6440
rect 4212 6400 4218 6412
rect 4430 6400 4436 6452
rect 4488 6440 4494 6452
rect 5261 6443 5319 6449
rect 5261 6440 5273 6443
rect 4488 6412 5273 6440
rect 4488 6400 4494 6412
rect 5261 6409 5273 6412
rect 5307 6409 5319 6443
rect 5261 6403 5319 6409
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6440 6699 6443
rect 7190 6440 7196 6452
rect 6687 6412 7196 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 7190 6400 7196 6412
rect 7248 6400 7254 6452
rect 8297 6443 8355 6449
rect 8297 6409 8309 6443
rect 8343 6440 8355 6443
rect 8386 6440 8392 6452
rect 8343 6412 8392 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 9950 6440 9956 6452
rect 9732 6412 9956 6440
rect 9732 6400 9738 6412
rect 9950 6400 9956 6412
rect 10008 6440 10014 6452
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 10008 6412 10057 6440
rect 10008 6400 10014 6412
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 10045 6403 10103 6409
rect 13357 6443 13415 6449
rect 13357 6409 13369 6443
rect 13403 6440 13415 6443
rect 13998 6440 14004 6452
rect 13403 6412 14004 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 15286 6440 15292 6452
rect 15247 6412 15292 6440
rect 15286 6400 15292 6412
rect 15344 6400 15350 6452
rect 16298 6440 16304 6452
rect 16259 6412 16304 6440
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 17681 6443 17739 6449
rect 17681 6409 17693 6443
rect 17727 6440 17739 6443
rect 17770 6440 17776 6452
rect 17727 6412 17776 6440
rect 17727 6409 17739 6412
rect 17681 6403 17739 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 21266 6440 21272 6452
rect 21227 6412 21272 6440
rect 21266 6400 21272 6412
rect 21324 6400 21330 6452
rect 23106 6440 23112 6452
rect 23067 6412 23112 6440
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 24946 6440 24952 6452
rect 24907 6412 24952 6440
rect 24946 6400 24952 6412
rect 25004 6400 25010 6452
rect 25314 6440 25320 6452
rect 25275 6412 25320 6440
rect 25314 6400 25320 6412
rect 25372 6400 25378 6452
rect 27157 6443 27215 6449
rect 27157 6409 27169 6443
rect 27203 6440 27215 6443
rect 27430 6440 27436 6452
rect 27203 6412 27436 6440
rect 27203 6409 27215 6412
rect 27157 6403 27215 6409
rect 27430 6400 27436 6412
rect 27488 6400 27494 6452
rect 28721 6443 28779 6449
rect 27632 6412 28212 6440
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 11977 6375 12035 6381
rect 11977 6372 11989 6375
rect 9824 6344 11989 6372
rect 9824 6332 9830 6344
rect 11977 6341 11989 6344
rect 12023 6372 12035 6375
rect 12158 6372 12164 6384
rect 12023 6344 12164 6372
rect 12023 6341 12035 6344
rect 11977 6335 12035 6341
rect 12158 6332 12164 6344
rect 12216 6332 12222 6384
rect 12250 6332 12256 6384
rect 12308 6372 12314 6384
rect 13446 6372 13452 6384
rect 12308 6344 13452 6372
rect 12308 6332 12314 6344
rect 13446 6332 13452 6344
rect 13504 6372 13510 6384
rect 14369 6375 14427 6381
rect 14369 6372 14381 6375
rect 13504 6344 14381 6372
rect 13504 6332 13510 6344
rect 14369 6341 14381 6344
rect 14415 6341 14427 6375
rect 14369 6335 14427 6341
rect 16022 6332 16028 6384
rect 16080 6372 16086 6384
rect 16945 6375 17003 6381
rect 16945 6372 16957 6375
rect 16080 6344 16957 6372
rect 16080 6332 16086 6344
rect 16945 6341 16957 6344
rect 16991 6341 17003 6375
rect 16945 6335 17003 6341
rect 17586 6332 17592 6384
rect 17644 6372 17650 6384
rect 18230 6372 18236 6384
rect 17644 6344 18236 6372
rect 17644 6332 17650 6344
rect 18230 6332 18236 6344
rect 18288 6332 18294 6384
rect 21821 6375 21879 6381
rect 21821 6372 21833 6375
rect 18340 6344 21833 6372
rect 2038 6304 2044 6316
rect 1412 6276 2044 6304
rect 1412 6245 1440 6276
rect 2038 6264 2044 6276
rect 2096 6264 2102 6316
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6304 2835 6307
rect 2866 6304 2872 6316
rect 2823 6276 2872 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 2866 6264 2872 6276
rect 2924 6264 2930 6316
rect 3050 6304 3056 6316
rect 3011 6276 3056 6304
rect 3050 6264 3056 6276
rect 3108 6264 3114 6316
rect 4430 6304 4436 6316
rect 3712 6276 4436 6304
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6205 1455 6239
rect 1397 6199 1455 6205
rect 2869 6171 2927 6177
rect 2869 6137 2881 6171
rect 2915 6168 2927 6171
rect 3142 6168 3148 6180
rect 2915 6140 3148 6168
rect 2915 6137 2927 6140
rect 2869 6131 2927 6137
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 2958 6060 2964 6112
rect 3016 6100 3022 6112
rect 3712 6109 3740 6276
rect 4430 6264 4436 6276
rect 4488 6264 4494 6316
rect 6273 6307 6331 6313
rect 6273 6273 6285 6307
rect 6319 6304 6331 6307
rect 7006 6304 7012 6316
rect 6319 6276 7012 6304
rect 6319 6273 6331 6276
rect 6273 6267 6331 6273
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 9030 6304 9036 6316
rect 7607 6276 9036 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 9030 6264 9036 6276
rect 9088 6304 9094 6316
rect 11057 6307 11115 6313
rect 11057 6304 11069 6307
rect 9088 6276 11069 6304
rect 9088 6264 9094 6276
rect 11057 6273 11069 6276
rect 11103 6273 11115 6307
rect 14734 6304 14740 6316
rect 14647 6276 14740 6304
rect 11057 6267 11115 6273
rect 14734 6264 14740 6276
rect 14792 6304 14798 6316
rect 16850 6304 16856 6316
rect 14792 6276 16856 6304
rect 14792 6264 14798 6276
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 17126 6264 17132 6316
rect 17184 6304 17190 6316
rect 18340 6304 18368 6344
rect 21821 6341 21833 6344
rect 21867 6341 21879 6375
rect 21821 6335 21879 6341
rect 18506 6304 18512 6316
rect 17184 6276 18368 6304
rect 18467 6276 18512 6304
rect 17184 6264 17190 6276
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 18690 6264 18696 6316
rect 18748 6304 18754 6316
rect 18785 6307 18843 6313
rect 18785 6304 18797 6307
rect 18748 6276 18797 6304
rect 18748 6264 18754 6276
rect 18785 6273 18797 6276
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 21836 6304 21864 6335
rect 23750 6332 23756 6384
rect 23808 6372 23814 6384
rect 27632 6372 27660 6412
rect 28074 6372 28080 6384
rect 23808 6344 27660 6372
rect 27724 6344 28080 6372
rect 23808 6332 23814 6344
rect 23474 6304 23480 6316
rect 21836 6276 23480 6304
rect 8662 6236 8668 6248
rect 8623 6208 8668 6236
rect 8662 6196 8668 6208
rect 8720 6196 8726 6248
rect 8849 6239 8907 6245
rect 8849 6205 8861 6239
rect 8895 6205 8907 6239
rect 8849 6199 8907 6205
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 12986 6236 12992 6248
rect 12483 6208 12992 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 4338 6168 4344 6180
rect 4299 6140 4344 6168
rect 4338 6128 4344 6140
rect 4396 6128 4402 6180
rect 4430 6128 4436 6180
rect 4488 6168 4494 6180
rect 4488 6140 4533 6168
rect 4488 6128 4494 6140
rect 4798 6128 4804 6180
rect 4856 6168 4862 6180
rect 4985 6171 5043 6177
rect 4985 6168 4997 6171
rect 4856 6140 4997 6168
rect 4856 6128 4862 6140
rect 4985 6137 4997 6140
rect 5031 6168 5043 6171
rect 6917 6171 6975 6177
rect 6917 6168 6929 6171
rect 5031 6140 6929 6168
rect 5031 6137 5043 6140
rect 4985 6131 5043 6137
rect 6917 6137 6929 6140
rect 6963 6137 6975 6171
rect 6917 6131 6975 6137
rect 3697 6103 3755 6109
rect 3697 6100 3709 6103
rect 3016 6072 3709 6100
rect 3016 6060 3022 6072
rect 3697 6069 3709 6072
rect 3743 6069 3755 6103
rect 6932 6100 6960 6131
rect 7006 6128 7012 6180
rect 7064 6168 7070 6180
rect 7064 6140 7109 6168
rect 7064 6128 7070 6140
rect 8386 6128 8392 6180
rect 8444 6168 8450 6180
rect 8864 6168 8892 6199
rect 12986 6196 12992 6208
rect 13044 6236 13050 6248
rect 13633 6239 13691 6245
rect 13633 6236 13645 6239
rect 13044 6208 13645 6236
rect 13044 6196 13050 6208
rect 13633 6205 13645 6208
rect 13679 6205 13691 6239
rect 14090 6236 14096 6248
rect 14003 6208 14096 6236
rect 13633 6199 13691 6205
rect 14090 6196 14096 6208
rect 14148 6236 14154 6248
rect 14185 6239 14243 6245
rect 14185 6236 14197 6239
rect 14148 6208 14197 6236
rect 14148 6196 14154 6208
rect 14185 6205 14197 6208
rect 14231 6205 14243 6239
rect 15378 6236 15384 6248
rect 15339 6208 15384 6236
rect 14185 6199 14243 6205
rect 10778 6168 10784 6180
rect 8444 6140 8892 6168
rect 10739 6140 10784 6168
rect 8444 6128 8450 6140
rect 10778 6128 10784 6140
rect 10836 6128 10842 6180
rect 10870 6128 10876 6180
rect 10928 6168 10934 6180
rect 12758 6171 12816 6177
rect 10928 6140 10973 6168
rect 10928 6128 10934 6140
rect 12758 6137 12770 6171
rect 12804 6168 12816 6171
rect 13078 6168 13084 6180
rect 12804 6140 13084 6168
rect 12804 6137 12816 6140
rect 12758 6131 12816 6137
rect 13078 6128 13084 6140
rect 13136 6168 13142 6180
rect 14200 6168 14228 6199
rect 15378 6196 15384 6208
rect 15436 6196 15442 6248
rect 17678 6236 17684 6248
rect 15488 6208 17684 6236
rect 15488 6168 15516 6208
rect 17678 6196 17684 6208
rect 17736 6196 17742 6248
rect 19981 6239 20039 6245
rect 19981 6205 19993 6239
rect 20027 6236 20039 6239
rect 20162 6236 20168 6248
rect 20027 6208 20168 6236
rect 20027 6205 20039 6208
rect 19981 6199 20039 6205
rect 20162 6196 20168 6208
rect 20220 6196 20226 6248
rect 21836 6236 21864 6276
rect 23474 6264 23480 6276
rect 23532 6264 23538 6316
rect 27724 6313 27752 6344
rect 28074 6332 28080 6344
rect 28132 6332 28138 6384
rect 28184 6372 28212 6412
rect 28721 6409 28733 6443
rect 28767 6440 28779 6443
rect 28810 6440 28816 6452
rect 28767 6412 28816 6440
rect 28767 6409 28779 6412
rect 28721 6403 28779 6409
rect 28810 6400 28816 6412
rect 28868 6400 28874 6452
rect 28902 6400 28908 6452
rect 28960 6440 28966 6452
rect 31021 6443 31079 6449
rect 31021 6440 31033 6443
rect 28960 6412 31033 6440
rect 28960 6400 28966 6412
rect 31021 6409 31033 6412
rect 31067 6440 31079 6443
rect 32950 6440 32956 6452
rect 31067 6412 32956 6440
rect 31067 6409 31079 6412
rect 31021 6403 31079 6409
rect 30466 6372 30472 6384
rect 28184 6344 30472 6372
rect 30466 6332 30472 6344
rect 30524 6332 30530 6384
rect 27709 6307 27767 6313
rect 27709 6273 27721 6307
rect 27755 6273 27767 6307
rect 27982 6304 27988 6316
rect 27943 6276 27988 6304
rect 27709 6267 27767 6273
rect 27982 6264 27988 6276
rect 28040 6264 28046 6316
rect 29178 6264 29184 6316
rect 29236 6304 29242 6316
rect 29638 6304 29644 6316
rect 29236 6276 29644 6304
rect 29236 6264 29242 6276
rect 29638 6264 29644 6276
rect 29696 6264 29702 6316
rect 22005 6239 22063 6245
rect 22005 6236 22017 6239
rect 21836 6208 22017 6236
rect 22005 6205 22017 6208
rect 22051 6205 22063 6239
rect 22005 6199 22063 6205
rect 22094 6196 22100 6248
rect 22152 6236 22158 6248
rect 22465 6239 22523 6245
rect 22465 6236 22477 6239
rect 22152 6208 22477 6236
rect 22152 6196 22158 6208
rect 22465 6205 22477 6208
rect 22511 6205 22523 6239
rect 23658 6236 23664 6248
rect 23619 6208 23664 6236
rect 22465 6199 22523 6205
rect 23658 6196 23664 6208
rect 23716 6196 23722 6248
rect 25866 6236 25872 6248
rect 25827 6208 25872 6236
rect 25866 6196 25872 6208
rect 25924 6196 25930 6248
rect 31128 6245 31156 6412
rect 32950 6400 32956 6412
rect 33008 6400 33014 6452
rect 33870 6440 33876 6452
rect 33831 6412 33876 6440
rect 33870 6400 33876 6412
rect 33928 6400 33934 6452
rect 36078 6400 36084 6452
rect 36136 6440 36142 6452
rect 36446 6440 36452 6452
rect 36136 6412 36452 6440
rect 36136 6400 36142 6412
rect 36446 6400 36452 6412
rect 36504 6440 36510 6452
rect 36587 6443 36645 6449
rect 36587 6440 36599 6443
rect 36504 6412 36599 6440
rect 36504 6400 36510 6412
rect 36587 6409 36599 6412
rect 36633 6409 36645 6443
rect 36587 6403 36645 6409
rect 32030 6332 32036 6384
rect 32088 6372 32094 6384
rect 32217 6375 32275 6381
rect 32217 6372 32229 6375
rect 32088 6344 32229 6372
rect 32088 6332 32094 6344
rect 32217 6341 32229 6344
rect 32263 6372 32275 6375
rect 32401 6375 32459 6381
rect 32401 6372 32413 6375
rect 32263 6344 32413 6372
rect 32263 6341 32275 6344
rect 32217 6335 32275 6341
rect 32401 6341 32413 6344
rect 32447 6372 32459 6375
rect 32493 6375 32551 6381
rect 32493 6372 32505 6375
rect 32447 6344 32505 6372
rect 32447 6341 32459 6344
rect 32401 6335 32459 6341
rect 32493 6341 32505 6344
rect 32539 6341 32551 6375
rect 32493 6335 32551 6341
rect 33042 6332 33048 6384
rect 33100 6372 33106 6384
rect 34241 6375 34299 6381
rect 34241 6372 34253 6375
rect 33100 6344 34253 6372
rect 33100 6332 33106 6344
rect 34241 6341 34253 6344
rect 34287 6372 34299 6375
rect 34606 6372 34612 6384
rect 34287 6344 34612 6372
rect 34287 6341 34299 6344
rect 34241 6335 34299 6341
rect 34606 6332 34612 6344
rect 34664 6372 34670 6384
rect 35989 6375 36047 6381
rect 35989 6372 36001 6375
rect 34664 6344 36001 6372
rect 34664 6332 34670 6344
rect 35989 6341 36001 6344
rect 36035 6372 36047 6375
rect 36170 6372 36176 6384
rect 36035 6344 36176 6372
rect 36035 6341 36047 6344
rect 35989 6335 36047 6341
rect 36170 6332 36176 6344
rect 36228 6332 36234 6384
rect 32122 6264 32128 6316
rect 32180 6304 32186 6316
rect 35158 6304 35164 6316
rect 32180 6276 35164 6304
rect 32180 6264 32186 6276
rect 35158 6264 35164 6276
rect 35216 6264 35222 6316
rect 35342 6304 35348 6316
rect 35303 6276 35348 6304
rect 35342 6264 35348 6276
rect 35400 6264 35406 6316
rect 31113 6239 31171 6245
rect 31113 6205 31125 6239
rect 31159 6205 31171 6239
rect 31113 6199 31171 6205
rect 31202 6196 31208 6248
rect 31260 6236 31266 6248
rect 31573 6239 31631 6245
rect 31573 6236 31585 6239
rect 31260 6208 31585 6236
rect 31260 6196 31266 6208
rect 31573 6205 31585 6208
rect 31619 6205 31631 6239
rect 31573 6199 31631 6205
rect 31849 6239 31907 6245
rect 31849 6205 31861 6239
rect 31895 6236 31907 6239
rect 32674 6236 32680 6248
rect 31895 6208 32680 6236
rect 31895 6205 31907 6208
rect 31849 6199 31907 6205
rect 32674 6196 32680 6208
rect 32732 6196 32738 6248
rect 33597 6239 33655 6245
rect 33597 6205 33609 6239
rect 33643 6236 33655 6239
rect 34606 6236 34612 6248
rect 33643 6208 34612 6236
rect 33643 6205 33655 6208
rect 33597 6199 33655 6205
rect 34606 6196 34612 6208
rect 34664 6196 34670 6248
rect 36516 6239 36574 6245
rect 36516 6205 36528 6239
rect 36562 6236 36574 6239
rect 36562 6208 36952 6236
rect 36562 6205 36574 6208
rect 36516 6199 36574 6205
rect 13136 6140 13814 6168
rect 14200 6140 15516 6168
rect 15702 6171 15760 6177
rect 13136 6128 13142 6140
rect 7837 6103 7895 6109
rect 7837 6100 7849 6103
rect 6932 6072 7849 6100
rect 3697 6063 3755 6069
rect 7837 6069 7849 6072
rect 7883 6069 7895 6103
rect 8478 6100 8484 6112
rect 8439 6072 8484 6100
rect 7837 6063 7895 6069
rect 8478 6060 8484 6072
rect 8536 6060 8542 6112
rect 9766 6100 9772 6112
rect 9727 6072 9772 6100
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10597 6103 10655 6109
rect 10597 6069 10609 6103
rect 10643 6100 10655 6103
rect 10888 6100 10916 6128
rect 10643 6072 10916 6100
rect 13786 6100 13814 6140
rect 15702 6137 15714 6171
rect 15748 6137 15760 6171
rect 18598 6168 18604 6180
rect 18559 6140 18604 6168
rect 15702 6131 15760 6137
rect 15286 6100 15292 6112
rect 13786 6072 15292 6100
rect 10643 6069 10655 6072
rect 10597 6063 10655 6069
rect 15286 6060 15292 6072
rect 15344 6100 15350 6112
rect 15717 6100 15745 6131
rect 18598 6128 18604 6140
rect 18656 6128 18662 6180
rect 19334 6128 19340 6180
rect 19392 6168 19398 6180
rect 19521 6171 19579 6177
rect 19521 6168 19533 6171
rect 19392 6140 19533 6168
rect 19392 6128 19398 6140
rect 19521 6137 19533 6140
rect 19567 6168 19579 6171
rect 19889 6171 19947 6177
rect 19889 6168 19901 6171
rect 19567 6140 19901 6168
rect 19567 6137 19579 6140
rect 19521 6131 19579 6137
rect 19889 6137 19901 6140
rect 19935 6168 19947 6171
rect 20343 6171 20401 6177
rect 20343 6168 20355 6171
rect 19935 6140 20355 6168
rect 19935 6137 19947 6140
rect 19889 6131 19947 6137
rect 20343 6137 20355 6140
rect 20389 6168 20401 6171
rect 21358 6168 21364 6180
rect 20389 6140 21364 6168
rect 20389 6137 20401 6140
rect 20343 6131 20401 6137
rect 21358 6128 21364 6140
rect 21416 6128 21422 6180
rect 24023 6171 24081 6177
rect 24023 6168 24035 6171
rect 23584 6140 24035 6168
rect 23584 6112 23612 6140
rect 24023 6137 24035 6140
rect 24069 6168 24081 6171
rect 24670 6168 24676 6180
rect 24069 6140 24676 6168
rect 24069 6137 24081 6140
rect 24023 6131 24081 6137
rect 24670 6128 24676 6140
rect 24728 6168 24734 6180
rect 25685 6171 25743 6177
rect 25685 6168 25697 6171
rect 24728 6140 25697 6168
rect 24728 6128 24734 6140
rect 25685 6137 25697 6140
rect 25731 6168 25743 6171
rect 26190 6171 26248 6177
rect 26190 6168 26202 6171
rect 25731 6140 26202 6168
rect 25731 6137 25743 6140
rect 25685 6131 25743 6137
rect 26190 6137 26202 6140
rect 26236 6137 26248 6171
rect 26190 6131 26248 6137
rect 27801 6171 27859 6177
rect 27801 6137 27813 6171
rect 27847 6168 27859 6171
rect 28810 6168 28816 6180
rect 27847 6140 28816 6168
rect 27847 6137 27859 6140
rect 27801 6131 27859 6137
rect 15344 6072 15745 6100
rect 15344 6060 15350 6072
rect 16206 6060 16212 6112
rect 16264 6100 16270 6112
rect 16577 6103 16635 6109
rect 16577 6100 16589 6103
rect 16264 6072 16589 6100
rect 16264 6060 16270 6072
rect 16577 6069 16589 6072
rect 16623 6069 16635 6103
rect 16577 6063 16635 6069
rect 20622 6060 20628 6112
rect 20680 6100 20686 6112
rect 20901 6103 20959 6109
rect 20901 6100 20913 6103
rect 20680 6072 20913 6100
rect 20680 6060 20686 6072
rect 20901 6069 20913 6072
rect 20947 6069 20959 6103
rect 22278 6100 22284 6112
rect 22239 6072 22284 6100
rect 20901 6063 20959 6069
rect 22278 6060 22284 6072
rect 22336 6060 22342 6112
rect 23477 6103 23535 6109
rect 23477 6069 23489 6103
rect 23523 6100 23535 6103
rect 23566 6100 23572 6112
rect 23523 6072 23572 6100
rect 23523 6069 23535 6072
rect 23477 6063 23535 6069
rect 23566 6060 23572 6072
rect 23624 6060 23630 6112
rect 24578 6100 24584 6112
rect 24539 6072 24584 6100
rect 24578 6060 24584 6072
rect 24636 6060 24642 6112
rect 26789 6103 26847 6109
rect 26789 6069 26801 6103
rect 26835 6100 26847 6103
rect 27525 6103 27583 6109
rect 27525 6100 27537 6103
rect 26835 6072 27537 6100
rect 26835 6069 26847 6072
rect 26789 6063 26847 6069
rect 27525 6069 27537 6072
rect 27571 6100 27583 6103
rect 27816 6100 27844 6131
rect 28810 6128 28816 6140
rect 28868 6128 28874 6180
rect 29362 6168 29368 6180
rect 29323 6140 29368 6168
rect 29362 6128 29368 6140
rect 29420 6128 29426 6180
rect 29457 6171 29515 6177
rect 29457 6137 29469 6171
rect 29503 6137 29515 6171
rect 29457 6131 29515 6137
rect 32401 6171 32459 6177
rect 32401 6137 32413 6171
rect 32447 6168 32459 6171
rect 32998 6171 33056 6177
rect 32998 6168 33010 6171
rect 32447 6140 33010 6168
rect 32447 6137 32459 6140
rect 32401 6131 32459 6137
rect 32998 6137 33010 6140
rect 33044 6137 33056 6171
rect 34974 6168 34980 6180
rect 34935 6140 34980 6168
rect 32998 6131 33056 6137
rect 28994 6100 29000 6112
rect 27571 6072 27844 6100
rect 28955 6072 29000 6100
rect 27571 6069 27583 6072
rect 27525 6063 27583 6069
rect 28994 6060 29000 6072
rect 29052 6100 29058 6112
rect 29472 6100 29500 6131
rect 34974 6128 34980 6140
rect 35032 6128 35038 6180
rect 35069 6171 35127 6177
rect 35069 6137 35081 6171
rect 35115 6137 35127 6171
rect 35069 6131 35127 6137
rect 29052 6072 29500 6100
rect 29052 6060 29058 6072
rect 34606 6060 34612 6112
rect 34664 6100 34670 6112
rect 35084 6100 35112 6131
rect 36924 6112 36952 6208
rect 36906 6100 36912 6112
rect 34664 6072 35112 6100
rect 36867 6072 36912 6100
rect 34664 6060 34670 6072
rect 36906 6060 36912 6072
rect 36964 6060 36970 6112
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 1673 5899 1731 5905
rect 1673 5865 1685 5899
rect 1719 5896 1731 5899
rect 2130 5896 2136 5908
rect 1719 5868 2136 5896
rect 1719 5865 1731 5868
rect 1673 5859 1731 5865
rect 2130 5856 2136 5868
rect 2188 5856 2194 5908
rect 2961 5899 3019 5905
rect 2961 5865 2973 5899
rect 3007 5896 3019 5899
rect 3142 5896 3148 5908
rect 3007 5868 3148 5896
rect 3007 5865 3019 5868
rect 2961 5859 3019 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3234 5856 3240 5908
rect 3292 5896 3298 5908
rect 3292 5868 3337 5896
rect 3292 5856 3298 5868
rect 3418 5856 3424 5908
rect 3476 5896 3482 5908
rect 4338 5896 4344 5908
rect 3476 5868 4344 5896
rect 3476 5856 3482 5868
rect 4338 5856 4344 5868
rect 4396 5896 4402 5908
rect 5077 5899 5135 5905
rect 5077 5896 5089 5899
rect 4396 5868 5089 5896
rect 4396 5856 4402 5868
rect 5077 5865 5089 5868
rect 5123 5865 5135 5899
rect 6730 5896 6736 5908
rect 6691 5868 6736 5896
rect 5077 5859 5135 5865
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7285 5899 7343 5905
rect 7285 5896 7297 5899
rect 6972 5868 7297 5896
rect 6972 5856 6978 5868
rect 7285 5865 7297 5868
rect 7331 5865 7343 5899
rect 7285 5859 7343 5865
rect 8481 5899 8539 5905
rect 8481 5865 8493 5899
rect 8527 5896 8539 5899
rect 8662 5896 8668 5908
rect 8527 5868 8668 5896
rect 8527 5865 8539 5868
rect 8481 5859 8539 5865
rect 8662 5856 8668 5868
rect 8720 5856 8726 5908
rect 10597 5899 10655 5905
rect 10597 5865 10609 5899
rect 10643 5896 10655 5899
rect 12066 5896 12072 5908
rect 10643 5868 12072 5896
rect 10643 5865 10655 5868
rect 10597 5859 10655 5865
rect 12066 5856 12072 5868
rect 12124 5896 12130 5908
rect 13078 5896 13084 5908
rect 12124 5868 12296 5896
rect 13039 5868 13084 5896
rect 12124 5856 12130 5868
rect 2038 5828 2044 5840
rect 1999 5800 2044 5828
rect 2038 5788 2044 5800
rect 2096 5788 2102 5840
rect 2682 5788 2688 5840
rect 2740 5828 2746 5840
rect 3252 5828 3280 5856
rect 2740 5800 3280 5828
rect 4249 5831 4307 5837
rect 2740 5788 2746 5800
rect 4249 5797 4261 5831
rect 4295 5828 4307 5831
rect 5810 5828 5816 5840
rect 4295 5800 5816 5828
rect 4295 5797 4307 5800
rect 4249 5791 4307 5797
rect 5810 5788 5816 5800
rect 5868 5788 5874 5840
rect 7484 5800 8610 5828
rect 3605 5763 3663 5769
rect 3605 5760 3617 5763
rect 2602 5732 3617 5760
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5692 2007 5695
rect 2602 5692 2630 5732
rect 3605 5729 3617 5732
rect 3651 5760 3663 5763
rect 3786 5760 3792 5772
rect 3651 5732 3792 5760
rect 3651 5729 3663 5732
rect 3605 5723 3663 5729
rect 3786 5720 3792 5732
rect 3844 5720 3850 5772
rect 4798 5720 4804 5772
rect 4856 5760 4862 5772
rect 7098 5760 7104 5772
rect 4856 5732 4901 5760
rect 7011 5732 7104 5760
rect 4856 5720 4862 5732
rect 7098 5720 7104 5732
rect 7156 5760 7162 5772
rect 7484 5769 7512 5800
rect 7469 5763 7527 5769
rect 7469 5760 7481 5763
rect 7156 5732 7481 5760
rect 7156 5720 7162 5732
rect 7469 5729 7481 5732
rect 7515 5729 7527 5763
rect 7469 5723 7527 5729
rect 7745 5763 7803 5769
rect 7745 5729 7757 5763
rect 7791 5760 7803 5763
rect 8386 5760 8392 5772
rect 7791 5732 8392 5760
rect 7791 5729 7803 5732
rect 7745 5723 7803 5729
rect 1995 5664 2630 5692
rect 1995 5661 2007 5664
rect 1949 5655 2007 5661
rect 3234 5652 3240 5704
rect 3292 5692 3298 5704
rect 4157 5695 4215 5701
rect 4157 5692 4169 5695
rect 3292 5664 4169 5692
rect 3292 5652 3298 5664
rect 4157 5661 4169 5664
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 2501 5627 2559 5633
rect 2501 5593 2513 5627
rect 2547 5624 2559 5627
rect 4816 5624 4844 5720
rect 5718 5692 5724 5704
rect 5679 5664 5724 5692
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 5997 5695 6055 5701
rect 5997 5661 6009 5695
rect 6043 5661 6055 5695
rect 5997 5655 6055 5661
rect 2547 5596 4844 5624
rect 2547 5593 2559 5596
rect 2501 5587 2559 5593
rect 5350 5584 5356 5636
rect 5408 5624 5414 5636
rect 6012 5624 6040 5655
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 7760 5692 7788 5723
rect 8386 5720 8392 5732
rect 8444 5720 8450 5772
rect 8582 5760 8610 5800
rect 9766 5788 9772 5840
rect 9824 5828 9830 5840
rect 12268 5837 12296 5868
rect 13078 5856 13084 5868
rect 13136 5856 13142 5908
rect 13541 5899 13599 5905
rect 13541 5865 13553 5899
rect 13587 5896 13599 5899
rect 13906 5896 13912 5908
rect 13587 5868 13912 5896
rect 13587 5865 13599 5868
rect 13541 5859 13599 5865
rect 13906 5856 13912 5868
rect 13964 5896 13970 5908
rect 14921 5899 14979 5905
rect 14921 5896 14933 5899
rect 13964 5868 14933 5896
rect 13964 5856 13970 5868
rect 14921 5865 14933 5868
rect 14967 5865 14979 5899
rect 14921 5859 14979 5865
rect 18509 5899 18567 5905
rect 18509 5865 18521 5899
rect 18555 5896 18567 5899
rect 18598 5896 18604 5908
rect 18555 5868 18604 5896
rect 18555 5865 18567 5868
rect 18509 5859 18567 5865
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 18690 5856 18696 5908
rect 18748 5896 18754 5908
rect 21450 5896 21456 5908
rect 18748 5868 21456 5896
rect 18748 5856 18754 5868
rect 21450 5856 21456 5868
rect 21508 5856 21514 5908
rect 22462 5896 22468 5908
rect 21652 5868 22468 5896
rect 9998 5831 10056 5837
rect 9998 5828 10010 5831
rect 9824 5800 10010 5828
rect 9824 5788 9830 5800
rect 9998 5797 10010 5800
rect 10044 5797 10056 5831
rect 9998 5791 10056 5797
rect 12253 5831 12311 5837
rect 12253 5797 12265 5831
rect 12299 5797 12311 5831
rect 12253 5791 12311 5797
rect 12894 5788 12900 5840
rect 12952 5828 12958 5840
rect 13446 5828 13452 5840
rect 12952 5800 13452 5828
rect 12952 5788 12958 5800
rect 13446 5788 13452 5800
rect 13504 5828 13510 5840
rect 13725 5831 13783 5837
rect 13725 5828 13737 5831
rect 13504 5800 13737 5828
rect 13504 5788 13510 5800
rect 13725 5797 13737 5800
rect 13771 5797 13783 5831
rect 13725 5791 13783 5797
rect 13817 5831 13875 5837
rect 13817 5797 13829 5831
rect 13863 5828 13875 5831
rect 14550 5828 14556 5840
rect 13863 5800 14556 5828
rect 13863 5797 13875 5800
rect 13817 5791 13875 5797
rect 14550 5788 14556 5800
rect 14608 5828 14614 5840
rect 15473 5831 15531 5837
rect 15473 5828 15485 5831
rect 14608 5800 15485 5828
rect 14608 5788 14614 5800
rect 15473 5797 15485 5800
rect 15519 5797 15531 5831
rect 16942 5828 16948 5840
rect 16903 5800 16948 5828
rect 15473 5791 15531 5797
rect 16942 5788 16948 5800
rect 17000 5788 17006 5840
rect 17037 5831 17095 5837
rect 17037 5797 17049 5831
rect 17083 5828 17095 5831
rect 18963 5831 19021 5837
rect 17083 5800 18000 5828
rect 17083 5797 17095 5800
rect 17037 5791 17095 5797
rect 10410 5760 10416 5772
rect 8582 5732 10416 5760
rect 10410 5720 10416 5732
rect 10468 5720 10474 5772
rect 9674 5692 9680 5704
rect 6696 5664 7788 5692
rect 9635 5664 9680 5692
rect 6696 5652 6702 5664
rect 9674 5652 9680 5664
rect 9732 5652 9738 5704
rect 12158 5692 12164 5704
rect 12119 5664 12164 5692
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5692 14427 5695
rect 14826 5692 14832 5704
rect 14415 5664 14832 5692
rect 14415 5661 14427 5664
rect 14369 5655 14427 5661
rect 14826 5652 14832 5664
rect 14884 5652 14890 5704
rect 14921 5695 14979 5701
rect 14921 5661 14933 5695
rect 14967 5692 14979 5695
rect 15381 5695 15439 5701
rect 15381 5692 15393 5695
rect 14967 5664 15393 5692
rect 14967 5661 14979 5664
rect 14921 5655 14979 5661
rect 15381 5661 15393 5664
rect 15427 5661 15439 5695
rect 15657 5695 15715 5701
rect 15657 5692 15669 5695
rect 15381 5655 15439 5661
rect 15488 5664 15669 5692
rect 10778 5624 10784 5636
rect 5408 5596 10784 5624
rect 5408 5584 5414 5596
rect 10778 5584 10784 5596
rect 10836 5624 10842 5636
rect 10873 5627 10931 5633
rect 10873 5624 10885 5627
rect 10836 5596 10885 5624
rect 10836 5584 10842 5596
rect 10873 5593 10885 5596
rect 10919 5593 10931 5627
rect 10873 5587 10931 5593
rect 12713 5627 12771 5633
rect 12713 5593 12725 5627
rect 12759 5624 12771 5627
rect 13814 5624 13820 5636
rect 12759 5596 13820 5624
rect 12759 5593 12771 5596
rect 12713 5587 12771 5593
rect 13814 5584 13820 5596
rect 13872 5624 13878 5636
rect 15488 5624 15516 5664
rect 15657 5661 15669 5664
rect 15703 5661 15715 5695
rect 15657 5655 15715 5661
rect 16114 5652 16120 5704
rect 16172 5692 16178 5704
rect 17221 5695 17279 5701
rect 17221 5692 17233 5695
rect 16172 5664 17233 5692
rect 16172 5652 16178 5664
rect 17221 5661 17233 5664
rect 17267 5661 17279 5695
rect 17221 5655 17279 5661
rect 17972 5633 18000 5800
rect 18963 5797 18975 5831
rect 19009 5828 19021 5831
rect 19334 5828 19340 5840
rect 19009 5800 19340 5828
rect 19009 5797 19021 5800
rect 18963 5791 19021 5797
rect 19334 5788 19340 5800
rect 19392 5788 19398 5840
rect 20622 5788 20628 5840
rect 20680 5828 20686 5840
rect 21652 5837 21680 5868
rect 22462 5856 22468 5868
rect 22520 5856 22526 5908
rect 23566 5896 23572 5908
rect 23527 5868 23572 5896
rect 23566 5856 23572 5868
rect 23624 5856 23630 5908
rect 23658 5856 23664 5908
rect 23716 5896 23722 5908
rect 24397 5899 24455 5905
rect 24397 5896 24409 5899
rect 23716 5868 24409 5896
rect 23716 5856 23722 5868
rect 24397 5865 24409 5868
rect 24443 5865 24455 5899
rect 26326 5896 26332 5908
rect 26287 5868 26332 5896
rect 24397 5859 24455 5865
rect 26326 5856 26332 5868
rect 26384 5896 26390 5908
rect 29178 5896 29184 5908
rect 26384 5868 29184 5896
rect 26384 5856 26390 5868
rect 29178 5856 29184 5868
rect 29236 5856 29242 5908
rect 31110 5896 31116 5908
rect 30668 5868 31116 5896
rect 21085 5831 21143 5837
rect 21085 5828 21097 5831
rect 20680 5800 21097 5828
rect 20680 5788 20686 5800
rect 21085 5797 21097 5800
rect 21131 5797 21143 5831
rect 21085 5791 21143 5797
rect 21637 5831 21695 5837
rect 21637 5797 21649 5831
rect 21683 5797 21695 5831
rect 21637 5791 21695 5797
rect 24578 5788 24584 5840
rect 24636 5828 24642 5840
rect 27157 5831 27215 5837
rect 27157 5828 27169 5831
rect 24636 5800 27169 5828
rect 24636 5788 24642 5800
rect 27157 5797 27169 5800
rect 27203 5828 27215 5831
rect 27522 5828 27528 5840
rect 27203 5800 27528 5828
rect 27203 5797 27215 5800
rect 27157 5791 27215 5797
rect 27522 5788 27528 5800
rect 27580 5788 27586 5840
rect 27709 5831 27767 5837
rect 27709 5797 27721 5831
rect 27755 5828 27767 5831
rect 27982 5828 27988 5840
rect 27755 5800 27988 5828
rect 27755 5797 27767 5800
rect 27709 5791 27767 5797
rect 27982 5788 27988 5800
rect 28040 5788 28046 5840
rect 28442 5788 28448 5840
rect 28500 5828 28506 5840
rect 28721 5831 28779 5837
rect 28721 5828 28733 5831
rect 28500 5800 28733 5828
rect 28500 5788 28506 5800
rect 28721 5797 28733 5800
rect 28767 5797 28779 5831
rect 28721 5791 28779 5797
rect 18322 5720 18328 5772
rect 18380 5760 18386 5772
rect 18601 5763 18659 5769
rect 18601 5760 18613 5763
rect 18380 5732 18613 5760
rect 18380 5720 18386 5732
rect 18601 5729 18613 5732
rect 18647 5729 18659 5763
rect 18601 5723 18659 5729
rect 24670 5720 24676 5772
rect 24728 5760 24734 5772
rect 24949 5763 25007 5769
rect 24949 5760 24961 5763
rect 24728 5732 24961 5760
rect 24728 5720 24734 5732
rect 24949 5729 24961 5732
rect 24995 5729 25007 5763
rect 25130 5760 25136 5772
rect 25091 5732 25136 5760
rect 24949 5723 25007 5729
rect 25130 5720 25136 5732
rect 25188 5720 25194 5772
rect 30098 5760 30104 5772
rect 30059 5732 30104 5760
rect 30098 5720 30104 5732
rect 30156 5720 30162 5772
rect 30190 5720 30196 5772
rect 30248 5760 30254 5772
rect 30668 5769 30696 5868
rect 31110 5856 31116 5868
rect 31168 5856 31174 5908
rect 32674 5896 32680 5908
rect 32635 5868 32680 5896
rect 32674 5856 32680 5868
rect 32732 5856 32738 5908
rect 33551 5899 33609 5905
rect 33551 5865 33563 5899
rect 33597 5896 33609 5899
rect 34146 5896 34152 5908
rect 33597 5868 34152 5896
rect 33597 5865 33609 5868
rect 33551 5859 33609 5865
rect 34146 5856 34152 5868
rect 34204 5896 34210 5908
rect 34241 5899 34299 5905
rect 34241 5896 34253 5899
rect 34204 5868 34253 5896
rect 34204 5856 34210 5868
rect 34241 5865 34253 5868
rect 34287 5865 34299 5899
rect 34241 5859 34299 5865
rect 34974 5856 34980 5908
rect 35032 5896 35038 5908
rect 35437 5899 35495 5905
rect 35437 5896 35449 5899
rect 35032 5868 35449 5896
rect 35032 5856 35038 5868
rect 35437 5865 35449 5868
rect 35483 5865 35495 5899
rect 36446 5896 36452 5908
rect 36407 5868 36452 5896
rect 35437 5859 35495 5865
rect 36446 5856 36452 5868
rect 36504 5856 36510 5908
rect 30837 5831 30895 5837
rect 30837 5797 30849 5831
rect 30883 5828 30895 5831
rect 33318 5828 33324 5840
rect 30883 5800 33324 5828
rect 30883 5797 30895 5800
rect 30837 5791 30895 5797
rect 33318 5788 33324 5800
rect 33376 5788 33382 5840
rect 34606 5828 34612 5840
rect 34567 5800 34612 5828
rect 34606 5788 34612 5800
rect 34664 5788 34670 5840
rect 35161 5831 35219 5837
rect 35161 5797 35173 5831
rect 35207 5828 35219 5831
rect 36354 5828 36360 5840
rect 35207 5800 36360 5828
rect 35207 5797 35219 5800
rect 35161 5791 35219 5797
rect 36354 5788 36360 5800
rect 36412 5788 36418 5840
rect 30653 5763 30711 5769
rect 30653 5760 30665 5763
rect 30248 5732 30665 5760
rect 30248 5720 30254 5732
rect 30653 5729 30665 5732
rect 30699 5729 30711 5763
rect 30653 5723 30711 5729
rect 32033 5763 32091 5769
rect 32033 5729 32045 5763
rect 32079 5760 32091 5763
rect 32122 5760 32128 5772
rect 32079 5732 32128 5760
rect 32079 5729 32091 5732
rect 32033 5723 32091 5729
rect 32122 5720 32128 5732
rect 32180 5720 32186 5772
rect 33480 5763 33538 5769
rect 33480 5729 33492 5763
rect 33526 5760 33538 5763
rect 33594 5760 33600 5772
rect 33526 5732 33600 5760
rect 33526 5729 33538 5732
rect 33480 5723 33538 5729
rect 33594 5720 33600 5732
rect 33652 5720 33658 5772
rect 36040 5763 36098 5769
rect 36040 5729 36052 5763
rect 36086 5760 36098 5763
rect 36262 5760 36268 5772
rect 36086 5732 36268 5760
rect 36086 5729 36098 5732
rect 36040 5723 36098 5729
rect 36262 5720 36268 5732
rect 36320 5720 36326 5772
rect 20806 5652 20812 5704
rect 20864 5692 20870 5704
rect 20993 5695 21051 5701
rect 20993 5692 21005 5695
rect 20864 5664 21005 5692
rect 20864 5652 20870 5664
rect 20993 5661 21005 5664
rect 21039 5661 21051 5695
rect 20993 5655 21051 5661
rect 22278 5652 22284 5704
rect 22336 5692 22342 5704
rect 23201 5695 23259 5701
rect 23201 5692 23213 5695
rect 22336 5664 23213 5692
rect 22336 5652 22342 5664
rect 23201 5661 23213 5664
rect 23247 5661 23259 5695
rect 25498 5692 25504 5704
rect 25459 5664 25504 5692
rect 23201 5655 23259 5661
rect 25498 5652 25504 5664
rect 25556 5652 25562 5704
rect 26881 5695 26939 5701
rect 26881 5661 26893 5695
rect 26927 5692 26939 5695
rect 27062 5692 27068 5704
rect 26927 5664 27068 5692
rect 26927 5661 26939 5664
rect 26881 5655 26939 5661
rect 27062 5652 27068 5664
rect 27120 5652 27126 5704
rect 28626 5692 28632 5704
rect 28587 5664 28632 5692
rect 28626 5652 28632 5664
rect 28684 5652 28690 5704
rect 29362 5652 29368 5704
rect 29420 5692 29426 5704
rect 29641 5695 29699 5701
rect 29641 5692 29653 5695
rect 29420 5664 29653 5692
rect 29420 5652 29426 5664
rect 29641 5661 29653 5664
rect 29687 5692 29699 5695
rect 32263 5695 32321 5701
rect 32263 5692 32275 5695
rect 29687 5664 32275 5692
rect 29687 5661 29699 5664
rect 29641 5655 29699 5661
rect 32263 5661 32275 5664
rect 32309 5661 32321 5695
rect 32263 5655 32321 5661
rect 34146 5652 34152 5704
rect 34204 5692 34210 5704
rect 34517 5695 34575 5701
rect 34517 5692 34529 5695
rect 34204 5664 34529 5692
rect 34204 5652 34210 5664
rect 34517 5661 34529 5664
rect 34563 5692 34575 5695
rect 36127 5695 36185 5701
rect 36127 5692 36139 5695
rect 34563 5664 36139 5692
rect 34563 5661 34575 5664
rect 34517 5655 34575 5661
rect 36127 5661 36139 5664
rect 36173 5661 36185 5695
rect 36127 5655 36185 5661
rect 13872 5596 15516 5624
rect 17957 5627 18015 5633
rect 13872 5584 13878 5596
rect 17957 5593 17969 5627
rect 18003 5624 18015 5627
rect 19521 5627 19579 5633
rect 19521 5624 19533 5627
rect 18003 5596 19533 5624
rect 18003 5593 18015 5596
rect 17957 5587 18015 5593
rect 19521 5593 19533 5596
rect 19567 5593 19579 5627
rect 19521 5587 19579 5593
rect 19610 5584 19616 5636
rect 19668 5624 19674 5636
rect 19889 5627 19947 5633
rect 19889 5624 19901 5627
rect 19668 5596 19901 5624
rect 19668 5584 19674 5596
rect 19889 5593 19901 5596
rect 19935 5624 19947 5627
rect 23106 5624 23112 5636
rect 19935 5596 23112 5624
rect 19935 5593 19947 5596
rect 19889 5587 19947 5593
rect 23106 5584 23112 5596
rect 23164 5584 23170 5636
rect 29178 5624 29184 5636
rect 29139 5596 29184 5624
rect 29178 5584 29184 5596
rect 29236 5584 29242 5636
rect 8570 5516 8576 5568
rect 8628 5556 8634 5568
rect 8849 5559 8907 5565
rect 8849 5556 8861 5559
rect 8628 5528 8861 5556
rect 8628 5516 8634 5528
rect 8849 5525 8861 5528
rect 8895 5556 8907 5559
rect 9030 5556 9036 5568
rect 8895 5528 9036 5556
rect 8895 5525 8907 5528
rect 8849 5519 8907 5525
rect 9030 5516 9036 5528
rect 9088 5516 9094 5568
rect 11974 5556 11980 5568
rect 11887 5528 11980 5556
rect 11974 5516 11980 5528
rect 12032 5556 12038 5568
rect 12342 5556 12348 5568
rect 12032 5528 12348 5556
rect 12032 5516 12038 5528
rect 12342 5516 12348 5528
rect 12400 5516 12406 5568
rect 14734 5556 14740 5568
rect 14695 5528 14740 5556
rect 14734 5516 14740 5528
rect 14792 5516 14798 5568
rect 15105 5559 15163 5565
rect 15105 5525 15117 5559
rect 15151 5556 15163 5559
rect 15378 5556 15384 5568
rect 15151 5528 15384 5556
rect 15151 5525 15163 5528
rect 15105 5519 15163 5525
rect 15378 5516 15384 5528
rect 15436 5556 15442 5568
rect 16298 5556 16304 5568
rect 15436 5528 16304 5556
rect 15436 5516 15442 5528
rect 16298 5516 16304 5528
rect 16356 5516 16362 5568
rect 16485 5559 16543 5565
rect 16485 5525 16497 5559
rect 16531 5556 16543 5559
rect 16666 5556 16672 5568
rect 16531 5528 16672 5556
rect 16531 5525 16543 5528
rect 16485 5519 16543 5525
rect 16666 5516 16672 5528
rect 16724 5556 16730 5568
rect 17770 5556 17776 5568
rect 16724 5528 17776 5556
rect 16724 5516 16730 5528
rect 17770 5516 17776 5528
rect 17828 5516 17834 5568
rect 20162 5556 20168 5568
rect 20123 5528 20168 5556
rect 20162 5516 20168 5528
rect 20220 5516 20226 5568
rect 20714 5556 20720 5568
rect 20675 5528 20720 5556
rect 20714 5516 20720 5528
rect 20772 5516 20778 5568
rect 22094 5556 22100 5568
rect 22055 5528 22100 5556
rect 22094 5516 22100 5528
rect 22152 5516 22158 5568
rect 24118 5556 24124 5568
rect 24079 5528 24124 5556
rect 24118 5516 24124 5528
rect 24176 5516 24182 5568
rect 25866 5556 25872 5568
rect 25827 5528 25872 5556
rect 25866 5516 25872 5528
rect 25924 5516 25930 5568
rect 28074 5556 28080 5568
rect 28035 5528 28080 5556
rect 28074 5516 28080 5528
rect 28132 5516 28138 5568
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 2038 5312 2044 5364
rect 2096 5352 2102 5364
rect 2501 5355 2559 5361
rect 2501 5352 2513 5355
rect 2096 5324 2513 5352
rect 2096 5312 2102 5324
rect 2501 5321 2513 5324
rect 2547 5321 2559 5355
rect 2501 5315 2559 5321
rect 3605 5355 3663 5361
rect 3605 5321 3617 5355
rect 3651 5352 3663 5355
rect 3694 5352 3700 5364
rect 3651 5324 3700 5352
rect 3651 5321 3663 5324
rect 3605 5315 3663 5321
rect 3694 5312 3700 5324
rect 3752 5312 3758 5364
rect 4617 5355 4675 5361
rect 4617 5321 4629 5355
rect 4663 5352 4675 5355
rect 4985 5355 5043 5361
rect 4985 5352 4997 5355
rect 4663 5324 4997 5352
rect 4663 5321 4675 5324
rect 4617 5315 4675 5321
rect 4985 5321 4997 5324
rect 5031 5352 5043 5355
rect 5629 5355 5687 5361
rect 5629 5352 5641 5355
rect 5031 5324 5641 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 5629 5321 5641 5324
rect 5675 5352 5687 5355
rect 5810 5352 5816 5364
rect 5675 5324 5816 5352
rect 5675 5321 5687 5324
rect 5629 5315 5687 5321
rect 5810 5312 5816 5324
rect 5868 5312 5874 5364
rect 5905 5355 5963 5361
rect 5905 5321 5917 5355
rect 5951 5352 5963 5355
rect 8662 5352 8668 5364
rect 5951 5324 8668 5352
rect 5951 5321 5963 5324
rect 5905 5315 5963 5321
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 10321 5355 10379 5361
rect 10321 5352 10333 5355
rect 9824 5324 10333 5352
rect 9824 5312 9830 5324
rect 10321 5321 10333 5324
rect 10367 5352 10379 5355
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 10367 5324 10425 5352
rect 10367 5321 10379 5324
rect 10321 5315 10379 5321
rect 10413 5321 10425 5324
rect 10459 5321 10471 5355
rect 12066 5352 12072 5364
rect 12027 5324 12072 5352
rect 10413 5315 10471 5321
rect 12066 5312 12072 5324
rect 12124 5352 12130 5364
rect 14185 5355 14243 5361
rect 12124 5324 13814 5352
rect 12124 5312 12130 5324
rect 3712 5216 3740 5312
rect 6638 5284 6644 5296
rect 6599 5256 6644 5284
rect 6638 5244 6644 5256
rect 6696 5244 6702 5296
rect 7285 5287 7343 5293
rect 7285 5253 7297 5287
rect 7331 5284 7343 5287
rect 7374 5284 7380 5296
rect 7331 5256 7380 5284
rect 7331 5253 7343 5256
rect 7285 5247 7343 5253
rect 7374 5244 7380 5256
rect 7432 5244 7438 5296
rect 9125 5287 9183 5293
rect 9125 5253 9137 5287
rect 9171 5284 9183 5287
rect 11422 5284 11428 5296
rect 9171 5256 11428 5284
rect 9171 5253 9183 5256
rect 9125 5247 9183 5253
rect 11422 5244 11428 5256
rect 11480 5244 11486 5296
rect 13786 5216 13814 5324
rect 14185 5321 14197 5355
rect 14231 5352 14243 5355
rect 14550 5352 14556 5364
rect 14231 5324 14556 5352
rect 14231 5321 14243 5324
rect 14185 5315 14243 5321
rect 14550 5312 14556 5324
rect 14608 5312 14614 5364
rect 17313 5355 17371 5361
rect 17313 5321 17325 5355
rect 17359 5352 17371 5355
rect 17770 5352 17776 5364
rect 17359 5324 17776 5352
rect 17359 5321 17371 5324
rect 17313 5315 17371 5321
rect 17770 5312 17776 5324
rect 17828 5352 17834 5364
rect 18325 5355 18383 5361
rect 18325 5352 18337 5355
rect 17828 5324 18337 5352
rect 17828 5312 17834 5324
rect 18325 5321 18337 5324
rect 18371 5321 18383 5355
rect 18325 5315 18383 5321
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 20530 5352 20536 5364
rect 19392 5324 19437 5352
rect 20491 5324 20536 5352
rect 19392 5312 19398 5324
rect 20530 5312 20536 5324
rect 20588 5312 20594 5364
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 20901 5355 20959 5361
rect 20901 5352 20913 5355
rect 20864 5324 20913 5352
rect 20864 5312 20870 5324
rect 20901 5321 20913 5324
rect 20947 5321 20959 5355
rect 20901 5315 20959 5321
rect 22278 5312 22284 5364
rect 22336 5352 22342 5364
rect 22465 5355 22523 5361
rect 22465 5352 22477 5355
rect 22336 5324 22477 5352
rect 22336 5312 22342 5324
rect 22465 5321 22477 5324
rect 22511 5321 22523 5355
rect 22465 5315 22523 5321
rect 24118 5312 24124 5364
rect 24176 5352 24182 5364
rect 26881 5355 26939 5361
rect 26881 5352 26893 5355
rect 24176 5324 26893 5352
rect 24176 5312 24182 5324
rect 26881 5321 26893 5324
rect 26927 5352 26939 5355
rect 27246 5352 27252 5364
rect 26927 5324 27252 5352
rect 26927 5321 26939 5324
rect 26881 5315 26939 5321
rect 27246 5312 27252 5324
rect 27304 5312 27310 5364
rect 27522 5312 27528 5364
rect 27580 5352 27586 5364
rect 28442 5352 28448 5364
rect 27580 5324 28448 5352
rect 27580 5312 27586 5324
rect 28442 5312 28448 5324
rect 28500 5352 28506 5364
rect 28537 5355 28595 5361
rect 28537 5352 28549 5355
rect 28500 5324 28549 5352
rect 28500 5312 28506 5324
rect 28537 5321 28549 5324
rect 28583 5321 28595 5355
rect 28537 5315 28595 5321
rect 28718 5312 28724 5364
rect 28776 5352 28782 5364
rect 29411 5355 29469 5361
rect 29411 5352 29423 5355
rect 28776 5324 29423 5352
rect 28776 5312 28782 5324
rect 29411 5321 29423 5324
rect 29457 5321 29469 5355
rect 29822 5352 29828 5364
rect 29783 5324 29828 5352
rect 29411 5315 29469 5321
rect 29822 5312 29828 5324
rect 29880 5312 29886 5364
rect 30098 5352 30104 5364
rect 30059 5324 30104 5352
rect 30098 5312 30104 5324
rect 30156 5312 30162 5364
rect 30742 5352 30748 5364
rect 30703 5324 30748 5352
rect 30742 5312 30748 5324
rect 30800 5312 30806 5364
rect 33505 5355 33563 5361
rect 33505 5321 33517 5355
rect 33551 5352 33563 5355
rect 33594 5352 33600 5364
rect 33551 5324 33600 5352
rect 33551 5321 33563 5324
rect 33505 5315 33563 5321
rect 33594 5312 33600 5324
rect 33652 5312 33658 5364
rect 34146 5352 34152 5364
rect 34107 5324 34152 5352
rect 34146 5312 34152 5324
rect 34204 5312 34210 5364
rect 34517 5355 34575 5361
rect 34517 5321 34529 5355
rect 34563 5352 34575 5355
rect 34606 5352 34612 5364
rect 34563 5324 34612 5352
rect 34563 5321 34575 5324
rect 34517 5315 34575 5321
rect 34606 5312 34612 5324
rect 34664 5312 34670 5364
rect 34974 5312 34980 5364
rect 35032 5352 35038 5364
rect 35161 5355 35219 5361
rect 35161 5352 35173 5355
rect 35032 5324 35173 5352
rect 35032 5312 35038 5324
rect 35161 5321 35173 5324
rect 35207 5321 35219 5355
rect 35161 5315 35219 5321
rect 35986 5312 35992 5364
rect 36044 5352 36050 5364
rect 36081 5355 36139 5361
rect 36081 5352 36093 5355
rect 36044 5324 36093 5352
rect 36044 5312 36050 5324
rect 36081 5321 36093 5324
rect 36127 5352 36139 5355
rect 36262 5352 36268 5364
rect 36127 5324 36268 5352
rect 36127 5321 36139 5324
rect 36081 5315 36139 5321
rect 36262 5312 36268 5324
rect 36320 5312 36326 5364
rect 25038 5284 25044 5296
rect 24999 5256 25044 5284
rect 25038 5244 25044 5256
rect 25096 5244 25102 5296
rect 26234 5284 26240 5296
rect 26195 5256 26240 5284
rect 26234 5244 26240 5256
rect 26292 5244 26298 5296
rect 27062 5244 27068 5296
rect 27120 5284 27126 5296
rect 30423 5287 30481 5293
rect 30423 5284 30435 5287
rect 27120 5256 30435 5284
rect 27120 5244 27126 5256
rect 30423 5253 30435 5256
rect 30469 5253 30481 5287
rect 30423 5247 30481 5253
rect 14734 5216 14740 5228
rect 3528 5188 4108 5216
rect 13786 5188 14504 5216
rect 14695 5188 14740 5216
rect 1581 5151 1639 5157
rect 1581 5117 1593 5151
rect 1627 5148 1639 5151
rect 1762 5148 1768 5160
rect 1627 5120 1768 5148
rect 1627 5117 1639 5120
rect 1581 5111 1639 5117
rect 1762 5108 1768 5120
rect 1820 5148 1826 5160
rect 2777 5151 2835 5157
rect 2777 5148 2789 5151
rect 1820 5120 2789 5148
rect 1820 5108 1826 5120
rect 2777 5117 2789 5120
rect 2823 5117 2835 5151
rect 2777 5111 2835 5117
rect 1943 5083 2001 5089
rect 1943 5049 1955 5083
rect 1989 5080 2001 5083
rect 3528 5080 3556 5188
rect 3694 5148 3700 5160
rect 3655 5120 3700 5148
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 4080 5089 4108 5188
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 5767 5120 6316 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 1989 5052 3556 5080
rect 4059 5083 4117 5089
rect 1989 5049 2001 5052
rect 1943 5043 2001 5049
rect 4059 5049 4071 5083
rect 4105 5049 4117 5083
rect 4059 5043 4117 5049
rect 3234 5012 3240 5024
rect 3195 4984 3240 5012
rect 3234 4972 3240 4984
rect 3292 4972 3298 5024
rect 6288 5021 6316 5120
rect 6362 5108 6368 5160
rect 6420 5148 6426 5160
rect 7101 5151 7159 5157
rect 7101 5148 7113 5151
rect 6420 5120 7113 5148
rect 6420 5108 6426 5120
rect 7101 5117 7113 5120
rect 7147 5148 7159 5151
rect 7561 5151 7619 5157
rect 7561 5148 7573 5151
rect 7147 5120 7573 5148
rect 7147 5117 7159 5120
rect 7101 5111 7159 5117
rect 7561 5117 7573 5120
rect 7607 5117 7619 5151
rect 7561 5111 7619 5117
rect 8205 5151 8263 5157
rect 8205 5117 8217 5151
rect 8251 5148 8263 5151
rect 8846 5148 8852 5160
rect 8251 5120 8852 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 8846 5108 8852 5120
rect 8904 5108 8910 5160
rect 10597 5151 10655 5157
rect 10597 5148 10609 5151
rect 10060 5120 10609 5148
rect 8110 5080 8116 5092
rect 8023 5052 8116 5080
rect 8110 5040 8116 5052
rect 8168 5080 8174 5092
rect 8567 5083 8625 5089
rect 8567 5080 8579 5083
rect 8168 5052 8579 5080
rect 8168 5040 8174 5052
rect 8567 5049 8579 5052
rect 8613 5080 8625 5083
rect 9677 5083 9735 5089
rect 9677 5080 9689 5083
rect 8613 5052 9689 5080
rect 8613 5049 8625 5052
rect 8567 5043 8625 5049
rect 9677 5049 9689 5052
rect 9723 5080 9735 5083
rect 9766 5080 9772 5092
rect 9723 5052 9772 5080
rect 9723 5049 9735 5052
rect 9677 5043 9735 5049
rect 9766 5040 9772 5052
rect 9824 5040 9830 5092
rect 10060 5024 10088 5120
rect 10597 5117 10609 5120
rect 10643 5117 10655 5151
rect 10597 5111 10655 5117
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 13872 5120 13917 5148
rect 13872 5108 13878 5120
rect 10321 5083 10379 5089
rect 10321 5049 10333 5083
rect 10367 5080 10379 5083
rect 10918 5083 10976 5089
rect 10918 5080 10930 5083
rect 10367 5052 10930 5080
rect 10367 5049 10379 5052
rect 10321 5043 10379 5049
rect 10918 5049 10930 5052
rect 10964 5049 10976 5083
rect 13170 5080 13176 5092
rect 13131 5052 13176 5080
rect 10918 5043 10976 5049
rect 13170 5040 13176 5052
rect 13228 5040 13234 5092
rect 13262 5040 13268 5092
rect 13320 5080 13326 5092
rect 14476 5080 14504 5188
rect 14734 5176 14740 5188
rect 14792 5176 14798 5228
rect 14826 5176 14832 5228
rect 14884 5216 14890 5228
rect 15381 5219 15439 5225
rect 15381 5216 15393 5219
rect 14884 5188 15393 5216
rect 14884 5176 14890 5188
rect 15381 5185 15393 5188
rect 15427 5216 15439 5219
rect 16942 5216 16948 5228
rect 15427 5188 16948 5216
rect 15427 5185 15439 5188
rect 15381 5179 15439 5185
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 18782 5176 18788 5228
rect 18840 5216 18846 5228
rect 20162 5216 20168 5228
rect 18840 5188 20024 5216
rect 20123 5188 20168 5216
rect 18840 5176 18846 5188
rect 16206 5148 16212 5160
rect 16167 5120 16212 5148
rect 16206 5108 16212 5120
rect 16264 5108 16270 5160
rect 16761 5151 16819 5157
rect 16761 5117 16773 5151
rect 16807 5148 16819 5151
rect 18138 5148 18144 5160
rect 16807 5120 18144 5148
rect 16807 5117 16819 5120
rect 16761 5111 16819 5117
rect 14826 5080 14832 5092
rect 13320 5052 13365 5080
rect 14476 5052 14832 5080
rect 13320 5040 13326 5052
rect 14826 5040 14832 5052
rect 14884 5040 14890 5092
rect 16117 5083 16175 5089
rect 16117 5080 16129 5083
rect 14936 5052 16129 5080
rect 6273 5015 6331 5021
rect 6273 4981 6285 5015
rect 6319 5012 6331 5015
rect 6454 5012 6460 5024
rect 6319 4984 6460 5012
rect 6319 4981 6331 4984
rect 6273 4975 6331 4981
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 10042 5012 10048 5024
rect 10003 4984 10048 5012
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 11517 5015 11575 5021
rect 11517 4981 11529 5015
rect 11563 5012 11575 5015
rect 12894 5012 12900 5024
rect 11563 4984 12900 5012
rect 11563 4981 11575 4984
rect 11517 4975 11575 4981
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 13814 4972 13820 5024
rect 13872 5012 13878 5024
rect 14936 5012 14964 5052
rect 16117 5049 16129 5052
rect 16163 5080 16175 5083
rect 16776 5080 16804 5111
rect 18138 5108 18144 5120
rect 18196 5108 18202 5160
rect 18233 5151 18291 5157
rect 18233 5117 18245 5151
rect 18279 5148 18291 5151
rect 18969 5151 19027 5157
rect 18969 5148 18981 5151
rect 18279 5120 18981 5148
rect 18279 5117 18291 5120
rect 18233 5111 18291 5117
rect 18969 5117 18981 5120
rect 19015 5148 19027 5151
rect 19242 5148 19248 5160
rect 19015 5120 19248 5148
rect 19015 5117 19027 5120
rect 18969 5111 19027 5117
rect 19242 5108 19248 5120
rect 19300 5108 19306 5160
rect 19610 5148 19616 5160
rect 19571 5120 19616 5148
rect 19610 5108 19616 5120
rect 19668 5108 19674 5160
rect 19996 5157 20024 5188
rect 20162 5176 20168 5188
rect 20220 5176 20226 5228
rect 19981 5151 20039 5157
rect 19981 5117 19993 5151
rect 20027 5148 20039 5151
rect 20530 5148 20536 5160
rect 20027 5120 20536 5148
rect 20027 5117 20039 5120
rect 19981 5111 20039 5117
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 20714 5108 20720 5160
rect 20772 5148 20778 5160
rect 21361 5151 21419 5157
rect 21361 5148 21373 5151
rect 20772 5120 21373 5148
rect 20772 5108 20778 5120
rect 21361 5117 21373 5120
rect 21407 5148 21419 5151
rect 21450 5148 21456 5160
rect 21407 5120 21456 5148
rect 21407 5117 21419 5120
rect 21361 5111 21419 5117
rect 21450 5108 21456 5120
rect 21508 5108 21514 5160
rect 23750 5148 23756 5160
rect 23711 5120 23756 5148
rect 23750 5108 23756 5120
rect 23808 5108 23814 5160
rect 24213 5151 24271 5157
rect 24213 5117 24225 5151
rect 24259 5117 24271 5151
rect 25056 5148 25084 5244
rect 25866 5216 25872 5228
rect 25827 5188 25872 5216
rect 25866 5176 25872 5188
rect 25924 5176 25930 5228
rect 25225 5151 25283 5157
rect 25225 5148 25237 5151
rect 25056 5120 25237 5148
rect 24213 5111 24271 5117
rect 25225 5117 25237 5120
rect 25271 5117 25283 5151
rect 25225 5111 25283 5117
rect 25777 5151 25835 5157
rect 25777 5117 25789 5151
rect 25823 5148 25835 5151
rect 26252 5148 26280 5244
rect 27801 5219 27859 5225
rect 27801 5185 27813 5219
rect 27847 5216 27859 5219
rect 27982 5216 27988 5228
rect 27847 5188 27988 5216
rect 27847 5185 27859 5188
rect 27801 5179 27859 5185
rect 27982 5176 27988 5188
rect 28040 5176 28046 5228
rect 28626 5176 28632 5228
rect 28684 5216 28690 5228
rect 28997 5219 29055 5225
rect 28997 5216 29009 5219
rect 28684 5188 29009 5216
rect 28684 5176 28690 5188
rect 28997 5185 29009 5188
rect 29043 5216 29055 5219
rect 31435 5219 31493 5225
rect 31435 5216 31447 5219
rect 29043 5188 31447 5216
rect 29043 5185 29055 5188
rect 28997 5179 29055 5185
rect 31435 5185 31447 5188
rect 31481 5185 31493 5219
rect 31754 5216 31760 5228
rect 31715 5188 31760 5216
rect 31435 5179 31493 5185
rect 31754 5176 31760 5188
rect 31812 5176 31818 5228
rect 25823 5120 26280 5148
rect 29340 5151 29398 5157
rect 25823 5117 25835 5120
rect 25777 5111 25835 5117
rect 29340 5117 29352 5151
rect 29386 5148 29398 5151
rect 29822 5148 29828 5160
rect 29386 5120 29828 5148
rect 29386 5117 29398 5120
rect 29340 5111 29398 5117
rect 16163 5052 16804 5080
rect 17865 5083 17923 5089
rect 16163 5049 16175 5052
rect 16117 5043 16175 5049
rect 17865 5049 17877 5083
rect 17911 5080 17923 5083
rect 18049 5083 18107 5089
rect 18049 5080 18061 5083
rect 17911 5052 18061 5080
rect 17911 5049 17923 5052
rect 17865 5043 17923 5049
rect 18049 5049 18061 5052
rect 18095 5080 18107 5083
rect 18506 5080 18512 5092
rect 18095 5052 18512 5080
rect 18095 5049 18107 5052
rect 18049 5043 18107 5049
rect 18506 5040 18512 5052
rect 18564 5040 18570 5092
rect 19702 5040 19708 5092
rect 19760 5080 19766 5092
rect 21269 5083 21327 5089
rect 21269 5080 21281 5083
rect 19760 5052 21281 5080
rect 19760 5040 19766 5052
rect 21269 5049 21281 5052
rect 21315 5049 21327 5083
rect 21269 5043 21327 5049
rect 22094 5040 22100 5092
rect 22152 5080 22158 5092
rect 22925 5083 22983 5089
rect 22925 5080 22937 5083
rect 22152 5052 22937 5080
rect 22152 5040 22158 5052
rect 22925 5049 22937 5052
rect 22971 5080 22983 5083
rect 24026 5080 24032 5092
rect 22971 5052 24032 5080
rect 22971 5049 22983 5052
rect 22925 5043 22983 5049
rect 24026 5040 24032 5052
rect 24084 5080 24090 5092
rect 24228 5080 24256 5111
rect 25314 5080 25320 5092
rect 24084 5052 25320 5080
rect 24084 5040 24090 5052
rect 25314 5040 25320 5052
rect 25372 5080 25378 5092
rect 25792 5080 25820 5111
rect 29822 5108 29828 5120
rect 29880 5108 29886 5160
rect 30352 5151 30410 5157
rect 30352 5117 30364 5151
rect 30398 5148 30410 5151
rect 30742 5148 30748 5160
rect 30398 5120 30748 5148
rect 30398 5117 30410 5120
rect 30352 5111 30410 5117
rect 30742 5108 30748 5120
rect 30800 5108 30806 5160
rect 31348 5151 31406 5157
rect 31348 5117 31360 5151
rect 31394 5148 31406 5151
rect 31772 5148 31800 5176
rect 31394 5120 31800 5148
rect 34952 5151 35010 5157
rect 31394 5117 31406 5120
rect 31348 5111 31406 5117
rect 34952 5117 34964 5151
rect 34998 5148 35010 5151
rect 34998 5120 35480 5148
rect 34998 5117 35010 5120
rect 34952 5111 35010 5117
rect 25372 5052 25820 5080
rect 27157 5083 27215 5089
rect 25372 5040 25378 5052
rect 27157 5049 27169 5083
rect 27203 5049 27215 5083
rect 27157 5043 27215 5049
rect 15746 5012 15752 5024
rect 13872 4984 14964 5012
rect 15707 4984 15752 5012
rect 13872 4972 13878 4984
rect 15746 4972 15752 4984
rect 15804 4972 15810 5024
rect 16298 5012 16304 5024
rect 16259 4984 16304 5012
rect 16298 4972 16304 4984
rect 16356 4972 16362 5024
rect 23293 5015 23351 5021
rect 23293 4981 23305 5015
rect 23339 5012 23351 5015
rect 23566 5012 23572 5024
rect 23339 4984 23572 5012
rect 23339 4981 23351 4984
rect 23293 4975 23351 4981
rect 23566 4972 23572 4984
rect 23624 4972 23630 5024
rect 23658 4972 23664 5024
rect 23716 5012 23722 5024
rect 23753 5015 23811 5021
rect 23753 5012 23765 5015
rect 23716 4984 23765 5012
rect 23716 4972 23722 4984
rect 23753 4981 23765 4984
rect 23799 4981 23811 5015
rect 24670 5012 24676 5024
rect 24631 4984 24676 5012
rect 23753 4975 23811 4981
rect 24670 4972 24676 4984
rect 24728 4972 24734 5024
rect 27172 5012 27200 5043
rect 27246 5040 27252 5092
rect 27304 5080 27310 5092
rect 28994 5080 29000 5092
rect 27304 5052 29000 5080
rect 27304 5040 27310 5052
rect 28994 5040 29000 5052
rect 29052 5040 29058 5092
rect 35452 5024 35480 5120
rect 28166 5012 28172 5024
rect 27172 4984 28172 5012
rect 28166 4972 28172 4984
rect 28224 4972 28230 5024
rect 32122 5012 32128 5024
rect 32083 4984 32128 5012
rect 32122 4972 32128 4984
rect 32180 4972 32186 5024
rect 35434 5012 35440 5024
rect 35395 4984 35440 5012
rect 35434 4972 35440 4984
rect 35492 4972 35498 5024
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 1949 4811 2007 4817
rect 1949 4777 1961 4811
rect 1995 4808 2007 4811
rect 2038 4808 2044 4820
rect 1995 4780 2044 4808
rect 1995 4777 2007 4780
rect 1949 4771 2007 4777
rect 2038 4768 2044 4780
rect 2096 4808 2102 4820
rect 2225 4811 2283 4817
rect 2225 4808 2237 4811
rect 2096 4780 2237 4808
rect 2096 4768 2102 4780
rect 2225 4777 2237 4780
rect 2271 4777 2283 4811
rect 3694 4808 3700 4820
rect 3655 4780 3700 4808
rect 2225 4771 2283 4777
rect 3694 4768 3700 4780
rect 3752 4808 3758 4820
rect 4157 4811 4215 4817
rect 4157 4808 4169 4811
rect 3752 4780 4169 4808
rect 3752 4768 3758 4780
rect 4157 4777 4169 4780
rect 4203 4777 4215 4811
rect 4157 4771 4215 4777
rect 5442 4768 5448 4820
rect 5500 4808 5506 4820
rect 5537 4811 5595 4817
rect 5537 4808 5549 4811
rect 5500 4780 5549 4808
rect 5500 4768 5506 4780
rect 5537 4777 5549 4780
rect 5583 4808 5595 4811
rect 5718 4808 5724 4820
rect 5583 4780 5724 4808
rect 5583 4777 5595 4780
rect 5537 4771 5595 4777
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 7653 4811 7711 4817
rect 7653 4808 7665 4811
rect 6880 4780 7665 4808
rect 6880 4768 6886 4780
rect 7653 4777 7665 4780
rect 7699 4777 7711 4811
rect 7653 4771 7711 4777
rect 9493 4811 9551 4817
rect 9493 4777 9505 4811
rect 9539 4808 9551 4811
rect 9674 4808 9680 4820
rect 9539 4780 9680 4808
rect 9539 4777 9551 4780
rect 9493 4771 9551 4777
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 11882 4768 11888 4820
rect 11940 4808 11946 4820
rect 11977 4811 12035 4817
rect 11977 4808 11989 4811
rect 11940 4780 11989 4808
rect 11940 4768 11946 4780
rect 11977 4777 11989 4780
rect 12023 4808 12035 4811
rect 12158 4808 12164 4820
rect 12023 4780 12164 4808
rect 12023 4777 12035 4780
rect 11977 4771 12035 4777
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 12342 4808 12348 4820
rect 12303 4780 12348 4808
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 13170 4808 13176 4820
rect 13131 4780 13176 4808
rect 13170 4768 13176 4780
rect 13228 4768 13234 4820
rect 13446 4808 13452 4820
rect 13407 4780 13452 4808
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 14737 4811 14795 4817
rect 14737 4777 14749 4811
rect 14783 4808 14795 4811
rect 14826 4808 14832 4820
rect 14783 4780 14832 4808
rect 14783 4777 14795 4780
rect 14737 4771 14795 4777
rect 14826 4768 14832 4780
rect 14884 4768 14890 4820
rect 16577 4811 16635 4817
rect 16577 4777 16589 4811
rect 16623 4808 16635 4811
rect 18138 4808 18144 4820
rect 16623 4780 18144 4808
rect 16623 4777 16635 4780
rect 16577 4771 16635 4777
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 18322 4768 18328 4820
rect 18380 4808 18386 4820
rect 19245 4811 19303 4817
rect 19245 4808 19257 4811
rect 18380 4780 19257 4808
rect 18380 4768 18386 4780
rect 19245 4777 19257 4780
rect 19291 4777 19303 4811
rect 20622 4808 20628 4820
rect 20583 4780 20628 4808
rect 19245 4771 19303 4777
rect 20622 4768 20628 4780
rect 20680 4768 20686 4820
rect 20806 4768 20812 4820
rect 20864 4808 20870 4820
rect 20901 4811 20959 4817
rect 20901 4808 20913 4811
rect 20864 4780 20913 4808
rect 20864 4768 20870 4780
rect 20901 4777 20913 4780
rect 20947 4777 20959 4811
rect 23750 4808 23756 4820
rect 23711 4780 23756 4808
rect 20901 4771 20959 4777
rect 23750 4768 23756 4780
rect 23808 4768 23814 4820
rect 27522 4808 27528 4820
rect 27483 4780 27528 4808
rect 27522 4768 27528 4780
rect 27580 4768 27586 4820
rect 28074 4768 28080 4820
rect 28132 4808 28138 4820
rect 29779 4811 29837 4817
rect 29779 4808 29791 4811
rect 28132 4780 29791 4808
rect 28132 4768 28138 4780
rect 29779 4777 29791 4780
rect 29825 4777 29837 4811
rect 30190 4808 30196 4820
rect 30151 4780 30196 4808
rect 29779 4771 29837 4777
rect 30190 4768 30196 4780
rect 30248 4768 30254 4820
rect 2593 4743 2651 4749
rect 2593 4709 2605 4743
rect 2639 4740 2651 4743
rect 2866 4740 2872 4752
rect 2639 4712 2872 4740
rect 2639 4709 2651 4712
rect 2593 4703 2651 4709
rect 2866 4700 2872 4712
rect 2924 4700 2930 4752
rect 4522 4740 4528 4752
rect 4356 4712 4528 4740
rect 1464 4675 1522 4681
rect 1464 4641 1476 4675
rect 1510 4672 1522 4675
rect 1670 4672 1676 4684
rect 1510 4644 1676 4672
rect 1510 4641 1522 4644
rect 1464 4635 1522 4641
rect 1670 4632 1676 4644
rect 1728 4632 1734 4684
rect 4356 4681 4384 4712
rect 4522 4700 4528 4712
rect 4580 4740 4586 4752
rect 5994 4740 6000 4752
rect 4580 4712 6000 4740
rect 4580 4700 4586 4712
rect 5994 4700 6000 4712
rect 6052 4700 6058 4752
rect 6362 4740 6368 4752
rect 6323 4712 6368 4740
rect 6362 4700 6368 4712
rect 6420 4700 6426 4752
rect 10226 4740 10232 4752
rect 9692 4712 10232 4740
rect 4341 4675 4399 4681
rect 4341 4641 4353 4675
rect 4387 4641 4399 4675
rect 4341 4635 4399 4641
rect 4617 4675 4675 4681
rect 4617 4641 4629 4675
rect 4663 4672 4675 4675
rect 4890 4672 4896 4684
rect 4663 4644 4896 4672
rect 4663 4641 4675 4644
rect 4617 4635 4675 4641
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 5258 4632 5264 4684
rect 5316 4672 5322 4684
rect 5629 4675 5687 4681
rect 5629 4672 5641 4675
rect 5316 4644 5641 4672
rect 5316 4632 5322 4644
rect 5629 4641 5641 4644
rect 5675 4641 5687 4675
rect 5902 4672 5908 4684
rect 5863 4644 5908 4672
rect 5629 4635 5687 4641
rect 5902 4632 5908 4644
rect 5960 4632 5966 4684
rect 7190 4672 7196 4684
rect 7151 4644 7196 4672
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 7469 4675 7527 4681
rect 7469 4641 7481 4675
rect 7515 4672 7527 4675
rect 8018 4672 8024 4684
rect 7515 4644 8024 4672
rect 7515 4641 7527 4644
rect 7469 4635 7527 4641
rect 8018 4632 8024 4644
rect 8076 4632 8082 4684
rect 9692 4681 9720 4712
rect 10226 4700 10232 4712
rect 10284 4700 10290 4752
rect 12894 4700 12900 4752
rect 12952 4740 12958 4752
rect 13262 4740 13268 4752
rect 12952 4712 13268 4740
rect 12952 4700 12958 4712
rect 13262 4700 13268 4712
rect 13320 4740 13326 4752
rect 13722 4740 13728 4752
rect 13320 4712 13728 4740
rect 13320 4700 13326 4712
rect 13722 4700 13728 4712
rect 13780 4740 13786 4752
rect 13817 4743 13875 4749
rect 13817 4740 13829 4743
rect 13780 4712 13829 4740
rect 13780 4700 13786 4712
rect 13817 4709 13829 4712
rect 13863 4709 13875 4743
rect 13817 4703 13875 4709
rect 14369 4743 14427 4749
rect 14369 4709 14381 4743
rect 14415 4740 14427 4743
rect 14918 4740 14924 4752
rect 14415 4712 14924 4740
rect 14415 4709 14427 4712
rect 14369 4703 14427 4709
rect 14918 4700 14924 4712
rect 14976 4700 14982 4752
rect 15289 4743 15347 4749
rect 15289 4709 15301 4743
rect 15335 4740 15347 4743
rect 15930 4740 15936 4752
rect 15335 4712 15936 4740
rect 15335 4709 15347 4712
rect 15289 4703 15347 4709
rect 15930 4700 15936 4712
rect 15988 4700 15994 4752
rect 16485 4743 16543 4749
rect 16485 4709 16497 4743
rect 16531 4740 16543 4743
rect 16758 4740 16764 4752
rect 16531 4712 16764 4740
rect 16531 4709 16543 4712
rect 16485 4703 16543 4709
rect 16758 4700 16764 4712
rect 16816 4700 16822 4752
rect 17773 4743 17831 4749
rect 17773 4709 17785 4743
rect 17819 4740 17831 4743
rect 18966 4740 18972 4752
rect 17819 4712 18644 4740
rect 18927 4712 18972 4740
rect 17819 4709 17831 4712
rect 17773 4703 17831 4709
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 9953 4675 10011 4681
rect 9953 4672 9965 4675
rect 9824 4644 9965 4672
rect 9824 4632 9830 4644
rect 9953 4641 9965 4644
rect 9999 4641 10011 4675
rect 12066 4672 12072 4684
rect 12027 4644 12072 4672
rect 9953 4635 10011 4641
rect 12066 4632 12072 4644
rect 12124 4632 12130 4684
rect 12434 4632 12440 4684
rect 12492 4672 12498 4684
rect 12529 4675 12587 4681
rect 12529 4672 12541 4675
rect 12492 4644 12541 4672
rect 12492 4632 12498 4644
rect 12529 4641 12541 4644
rect 12575 4641 12587 4675
rect 12529 4635 12587 4641
rect 15105 4675 15163 4681
rect 15105 4641 15117 4675
rect 15151 4672 15163 4675
rect 15473 4675 15531 4681
rect 15473 4672 15485 4675
rect 15151 4644 15485 4672
rect 15151 4641 15163 4644
rect 15105 4635 15163 4641
rect 15473 4641 15485 4644
rect 15519 4672 15531 4675
rect 16666 4672 16672 4684
rect 15519 4644 16672 4672
rect 15519 4641 15531 4644
rect 15473 4635 15531 4641
rect 16666 4632 16672 4644
rect 16724 4632 16730 4684
rect 16776 4672 16804 4700
rect 18616 4684 18644 4712
rect 18966 4700 18972 4712
rect 19024 4700 19030 4752
rect 21726 4700 21732 4752
rect 21784 4740 21790 4752
rect 25501 4743 25559 4749
rect 21784 4712 23474 4740
rect 21784 4700 21790 4712
rect 16776 4644 17080 4672
rect 2501 4607 2559 4613
rect 2501 4573 2513 4607
rect 2547 4604 2559 4607
rect 2958 4604 2964 4616
rect 2547 4576 2964 4604
rect 2547 4573 2559 4576
rect 2501 4567 2559 4573
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 3142 4604 3148 4616
rect 3103 4576 3148 4604
rect 3142 4564 3148 4576
rect 3200 4604 3206 4616
rect 5350 4604 5356 4616
rect 3200 4576 5356 4604
rect 3200 4564 3206 4576
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 10137 4607 10195 4613
rect 10137 4604 10149 4607
rect 8582 4576 10149 4604
rect 1535 4539 1593 4545
rect 1535 4505 1547 4539
rect 1581 4536 1593 4539
rect 1946 4536 1952 4548
rect 1581 4508 1952 4536
rect 1581 4505 1593 4508
rect 1535 4499 1593 4505
rect 1946 4496 1952 4508
rect 2004 4496 2010 4548
rect 5718 4536 5724 4548
rect 5679 4508 5724 4536
rect 5718 4496 5724 4508
rect 5776 4536 5782 4548
rect 7009 4539 7067 4545
rect 7009 4536 7021 4539
rect 5776 4508 7021 4536
rect 5776 4496 5782 4508
rect 7009 4505 7021 4508
rect 7055 4536 7067 4539
rect 7098 4536 7104 4548
rect 7055 4508 7104 4536
rect 7055 4505 7067 4508
rect 7009 4499 7067 4505
rect 7098 4496 7104 4508
rect 7156 4536 7162 4548
rect 7285 4539 7343 4545
rect 7285 4536 7297 4539
rect 7156 4508 7297 4536
rect 7156 4496 7162 4508
rect 7285 4505 7297 4508
rect 7331 4505 7343 4539
rect 8582 4536 8610 4576
rect 10137 4573 10149 4576
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 13725 4607 13783 4613
rect 13725 4573 13737 4607
rect 13771 4604 13783 4607
rect 13998 4604 14004 4616
rect 13771 4576 14004 4604
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 13998 4564 14004 4576
rect 14056 4564 14062 4616
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4604 15899 4607
rect 16574 4604 16580 4616
rect 15887 4576 16580 4604
rect 15887 4573 15899 4576
rect 15841 4567 15899 4573
rect 16574 4564 16580 4576
rect 16632 4564 16638 4616
rect 16816 4607 16874 4613
rect 16816 4573 16828 4607
rect 16862 4604 16874 4607
rect 16942 4604 16948 4616
rect 16862 4576 16948 4604
rect 16862 4573 16874 4576
rect 16816 4567 16874 4573
rect 16942 4564 16948 4576
rect 17000 4564 17006 4616
rect 17052 4613 17080 4644
rect 17678 4632 17684 4684
rect 17736 4672 17742 4684
rect 18233 4675 18291 4681
rect 18233 4672 18245 4675
rect 17736 4644 18245 4672
rect 17736 4632 17742 4644
rect 18233 4641 18245 4644
rect 18279 4641 18291 4675
rect 18233 4635 18291 4641
rect 18598 4632 18604 4684
rect 18656 4672 18662 4684
rect 18782 4672 18788 4684
rect 18656 4644 18788 4672
rect 18656 4632 18662 4644
rect 18782 4632 18788 4644
rect 18840 4632 18846 4684
rect 18874 4632 18880 4684
rect 18932 4672 18938 4684
rect 19797 4675 19855 4681
rect 19797 4672 19809 4675
rect 18932 4644 19809 4672
rect 18932 4632 18938 4644
rect 19797 4641 19809 4644
rect 19843 4672 19855 4675
rect 20257 4675 20315 4681
rect 20257 4672 20269 4675
rect 19843 4644 20269 4672
rect 19843 4641 19855 4644
rect 19797 4635 19855 4641
rect 20257 4641 20269 4644
rect 20303 4641 20315 4675
rect 22097 4675 22155 4681
rect 22097 4672 22109 4675
rect 20257 4635 20315 4641
rect 21652 4644 22109 4672
rect 17037 4607 17095 4613
rect 17037 4573 17049 4607
rect 17083 4604 17095 4607
rect 18049 4607 18107 4613
rect 18049 4604 18061 4607
rect 17083 4576 18061 4604
rect 17083 4573 17095 4576
rect 17037 4567 17095 4573
rect 18049 4573 18061 4576
rect 18095 4573 18107 4607
rect 18049 4567 18107 4573
rect 18322 4564 18328 4616
rect 18380 4604 18386 4616
rect 21652 4604 21680 4644
rect 22097 4641 22109 4644
rect 22143 4672 22155 4675
rect 22186 4672 22192 4684
rect 22143 4644 22192 4672
rect 22143 4641 22155 4644
rect 22097 4635 22155 4641
rect 22186 4632 22192 4644
rect 22244 4632 22250 4684
rect 22922 4672 22928 4684
rect 22883 4644 22928 4672
rect 22922 4632 22928 4644
rect 22980 4632 22986 4684
rect 23446 4672 23474 4712
rect 25501 4709 25513 4743
rect 25547 4740 25559 4743
rect 26694 4740 26700 4752
rect 25547 4712 26700 4740
rect 25547 4709 25559 4712
rect 25501 4703 25559 4709
rect 26694 4700 26700 4712
rect 26752 4700 26758 4752
rect 28813 4743 28871 4749
rect 28813 4709 28825 4743
rect 28859 4740 28871 4743
rect 29454 4740 29460 4752
rect 28859 4712 29460 4740
rect 28859 4709 28871 4712
rect 28813 4703 28871 4709
rect 29454 4700 29460 4712
rect 29512 4700 29518 4752
rect 24946 4672 24952 4684
rect 23446 4644 24952 4672
rect 24946 4632 24952 4644
rect 25004 4632 25010 4684
rect 25314 4672 25320 4684
rect 25275 4644 25320 4672
rect 25314 4632 25320 4644
rect 25372 4632 25378 4684
rect 27154 4672 27160 4684
rect 27115 4644 27160 4672
rect 27154 4632 27160 4644
rect 27212 4632 27218 4684
rect 28258 4672 28264 4684
rect 28219 4644 28264 4672
rect 28258 4632 28264 4644
rect 28316 4632 28322 4684
rect 28629 4675 28687 4681
rect 28629 4641 28641 4675
rect 28675 4641 28687 4675
rect 29638 4672 29644 4684
rect 29599 4644 29644 4672
rect 28629 4635 28687 4641
rect 18380 4576 21680 4604
rect 21729 4607 21787 4613
rect 18380 4564 18386 4576
rect 21729 4573 21741 4607
rect 21775 4604 21787 4607
rect 22370 4604 22376 4616
rect 21775 4576 22376 4604
rect 21775 4573 21787 4576
rect 21729 4567 21787 4573
rect 22370 4564 22376 4576
rect 22428 4604 22434 4616
rect 22833 4607 22891 4613
rect 22833 4604 22845 4607
rect 22428 4576 22845 4604
rect 22428 4564 22434 4576
rect 22833 4573 22845 4576
rect 22879 4573 22891 4607
rect 22833 4567 22891 4573
rect 23382 4564 23388 4616
rect 23440 4604 23446 4616
rect 25130 4604 25136 4616
rect 23440 4576 25136 4604
rect 23440 4564 23446 4576
rect 25130 4564 25136 4576
rect 25188 4604 25194 4616
rect 25777 4607 25835 4613
rect 25777 4604 25789 4607
rect 25188 4576 25789 4604
rect 25188 4564 25194 4576
rect 25777 4573 25789 4576
rect 25823 4573 25835 4607
rect 26510 4604 26516 4616
rect 26471 4576 26516 4604
rect 25777 4567 25835 4573
rect 26510 4564 26516 4576
rect 26568 4564 26574 4616
rect 27706 4564 27712 4616
rect 27764 4604 27770 4616
rect 28644 4604 28672 4635
rect 29638 4632 29644 4644
rect 29696 4632 29702 4684
rect 30190 4604 30196 4616
rect 27764 4576 30196 4604
rect 27764 4564 27770 4576
rect 30190 4564 30196 4576
rect 30248 4564 30254 4616
rect 7285 4499 7343 4505
rect 7392 4508 8610 4536
rect 9769 4539 9827 4545
rect 5810 4428 5816 4480
rect 5868 4468 5874 4480
rect 7392 4468 7420 4508
rect 9769 4505 9781 4539
rect 9815 4536 9827 4539
rect 9858 4536 9864 4548
rect 9815 4508 9864 4536
rect 9815 4505 9827 4508
rect 9769 4499 9827 4505
rect 9858 4496 9864 4508
rect 9916 4496 9922 4548
rect 10410 4496 10416 4548
rect 10468 4536 10474 4548
rect 10781 4539 10839 4545
rect 10781 4536 10793 4539
rect 10468 4508 10793 4536
rect 10468 4496 10474 4508
rect 10781 4505 10793 4508
rect 10827 4536 10839 4539
rect 16206 4536 16212 4548
rect 10827 4508 16212 4536
rect 10827 4505 10839 4508
rect 10781 4499 10839 4505
rect 16206 4496 16212 4508
rect 16264 4496 16270 4548
rect 16482 4496 16488 4548
rect 16540 4536 16546 4548
rect 19981 4539 20039 4545
rect 19981 4536 19993 4539
rect 16540 4508 19993 4536
rect 16540 4496 16546 4508
rect 19981 4505 19993 4508
rect 20027 4505 20039 4539
rect 19981 4499 20039 4505
rect 23201 4539 23259 4545
rect 23201 4505 23213 4539
rect 23247 4536 23259 4539
rect 27430 4536 27436 4548
rect 23247 4508 27436 4536
rect 23247 4505 23259 4508
rect 23201 4499 23259 4505
rect 27430 4496 27436 4508
rect 27488 4496 27494 4548
rect 8386 4468 8392 4480
rect 5868 4440 7420 4468
rect 8347 4440 8392 4468
rect 5868 4428 5874 4440
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 8846 4468 8852 4480
rect 8759 4440 8852 4468
rect 8846 4428 8852 4440
rect 8904 4468 8910 4480
rect 9306 4468 9312 4480
rect 8904 4440 9312 4468
rect 8904 4428 8910 4440
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 16298 4428 16304 4480
rect 16356 4468 16362 4480
rect 16577 4471 16635 4477
rect 16577 4468 16589 4471
rect 16356 4440 16589 4468
rect 16356 4428 16362 4440
rect 16577 4437 16589 4440
rect 16623 4468 16635 4471
rect 16945 4471 17003 4477
rect 16945 4468 16957 4471
rect 16623 4440 16957 4468
rect 16623 4437 16635 4440
rect 16577 4431 16635 4437
rect 16945 4437 16957 4440
rect 16991 4437 17003 4471
rect 17126 4468 17132 4480
rect 17087 4440 17132 4468
rect 16945 4431 17003 4437
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 19705 4471 19763 4477
rect 19705 4437 19717 4471
rect 19751 4468 19763 4471
rect 19886 4468 19892 4480
rect 19751 4440 19892 4468
rect 19751 4437 19763 4440
rect 19705 4431 19763 4437
rect 19886 4428 19892 4440
rect 19944 4428 19950 4480
rect 24486 4468 24492 4480
rect 24447 4440 24492 4468
rect 24486 4428 24492 4440
rect 24544 4428 24550 4480
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 1670 4264 1676 4276
rect 1631 4236 1676 4264
rect 1670 4224 1676 4236
rect 1728 4224 1734 4276
rect 2866 4264 2872 4276
rect 2827 4236 2872 4264
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 4522 4264 4528 4276
rect 4483 4236 4528 4264
rect 4522 4224 4528 4236
rect 4580 4224 4586 4276
rect 5261 4267 5319 4273
rect 5261 4233 5273 4267
rect 5307 4264 5319 4267
rect 5718 4264 5724 4276
rect 5307 4236 5724 4264
rect 5307 4233 5319 4236
rect 5261 4227 5319 4233
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 7098 4264 7104 4276
rect 7059 4236 7104 4264
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 10226 4264 10232 4276
rect 9876 4236 10232 4264
rect 5629 4199 5687 4205
rect 5629 4165 5641 4199
rect 5675 4196 5687 4199
rect 5902 4196 5908 4208
rect 5675 4168 5908 4196
rect 5675 4165 5687 4168
rect 5629 4159 5687 4165
rect 5902 4156 5908 4168
rect 5960 4196 5966 4208
rect 6365 4199 6423 4205
rect 6365 4196 6377 4199
rect 5960 4168 6377 4196
rect 5960 4156 5966 4168
rect 6365 4165 6377 4168
rect 6411 4165 6423 4199
rect 6638 4196 6644 4208
rect 6365 4159 6423 4165
rect 6564 4168 6644 4196
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 3142 4128 3148 4140
rect 2639 4100 3148 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4128 3387 4131
rect 5994 4128 6000 4140
rect 3375 4100 6000 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 3694 4060 3700 4072
rect 3655 4032 3700 4060
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 3896 4069 3924 4100
rect 5994 4088 6000 4100
rect 6052 4128 6058 4140
rect 6564 4128 6592 4168
rect 6638 4156 6644 4168
rect 6696 4156 6702 4208
rect 9677 4199 9735 4205
rect 9677 4196 9689 4199
rect 8541 4168 9689 4196
rect 6052 4100 6592 4128
rect 6052 4088 6058 4100
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 8541 4128 8569 4168
rect 9677 4165 9689 4168
rect 9723 4196 9735 4199
rect 9876 4196 9904 4236
rect 10226 4224 10232 4236
rect 10284 4264 10290 4276
rect 11974 4264 11980 4276
rect 10284 4236 11980 4264
rect 10284 4224 10290 4236
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 12253 4267 12311 4273
rect 12253 4233 12265 4267
rect 12299 4264 12311 4267
rect 12342 4264 12348 4276
rect 12299 4236 12348 4264
rect 12299 4233 12311 4236
rect 12253 4227 12311 4233
rect 12342 4224 12348 4236
rect 12400 4264 12406 4276
rect 12618 4264 12624 4276
rect 12400 4236 12624 4264
rect 12400 4224 12406 4236
rect 12618 4224 12624 4236
rect 12676 4224 12682 4276
rect 13722 4264 13728 4276
rect 13683 4236 13728 4264
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 16298 4264 16304 4276
rect 16259 4236 16304 4264
rect 16298 4224 16304 4236
rect 16356 4224 16362 4276
rect 16390 4224 16396 4276
rect 16448 4264 16454 4276
rect 19886 4264 19892 4276
rect 16448 4236 16988 4264
rect 16448 4224 16454 4236
rect 9723 4168 9904 4196
rect 9723 4165 9735 4168
rect 9677 4159 9735 4165
rect 9950 4156 9956 4208
rect 10008 4196 10014 4208
rect 11885 4199 11943 4205
rect 10008 4168 10088 4196
rect 10008 4156 10014 4168
rect 7432 4100 8569 4128
rect 10060 4128 10088 4168
rect 11885 4165 11897 4199
rect 11931 4196 11943 4199
rect 12066 4196 12072 4208
rect 11931 4168 12072 4196
rect 11931 4165 11943 4168
rect 11885 4159 11943 4165
rect 12066 4156 12072 4168
rect 12124 4156 12130 4208
rect 16316 4196 16344 4224
rect 16960 4208 16988 4236
rect 19306 4236 19892 4264
rect 15488 4168 16344 4196
rect 16669 4199 16727 4205
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 10060 4100 10517 4128
rect 7432 4088 7438 4100
rect 10505 4097 10517 4100
rect 10551 4097 10563 4131
rect 12986 4128 12992 4140
rect 12947 4100 12992 4128
rect 10505 4091 10563 4097
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 13998 4128 14004 4140
rect 13959 4100 14004 4128
rect 13998 4088 14004 4100
rect 14056 4088 14062 4140
rect 3881 4063 3939 4069
rect 3881 4029 3893 4063
rect 3927 4029 3939 4063
rect 4890 4060 4896 4072
rect 4851 4032 4896 4060
rect 3881 4023 3939 4029
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 5721 4063 5779 4069
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 5810 4060 5816 4072
rect 5767 4032 5816 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 5810 4020 5816 4032
rect 5868 4020 5874 4072
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 7466 4060 7472 4072
rect 6687 4032 7472 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 8386 4060 8392 4072
rect 8347 4032 8392 4060
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8478 4020 8484 4072
rect 8536 4060 8542 4072
rect 8665 4063 8723 4069
rect 8536 4032 8581 4060
rect 8536 4020 8542 4032
rect 8665 4029 8677 4063
rect 8711 4029 8723 4063
rect 9950 4060 9956 4072
rect 8665 4023 8723 4029
rect 9140 4032 9956 4060
rect 1946 3992 1952 4004
rect 1907 3964 1952 3992
rect 1946 3952 1952 3964
rect 2004 3952 2010 4004
rect 2038 3952 2044 4004
rect 2096 3992 2102 4004
rect 2096 3964 2141 3992
rect 2096 3952 2102 3964
rect 4522 3952 4528 4004
rect 4580 3992 4586 4004
rect 6086 3992 6092 4004
rect 4580 3964 6092 3992
rect 4580 3952 4586 3964
rect 3510 3924 3516 3936
rect 3471 3896 3516 3924
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 5920 3933 5948 3964
rect 6086 3952 6092 3964
rect 6144 3952 6150 4004
rect 8680 3992 8708 4023
rect 8220 3964 8708 3992
rect 5905 3927 5963 3933
rect 5905 3893 5917 3927
rect 5951 3893 5963 3927
rect 6178 3924 6184 3936
rect 6139 3896 6184 3924
rect 5905 3887 5963 3893
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 6365 3927 6423 3933
rect 6365 3893 6377 3927
rect 6411 3924 6423 3927
rect 7650 3924 7656 3936
rect 6411 3896 7656 3924
rect 6411 3893 6423 3896
rect 6365 3887 6423 3893
rect 7650 3884 7656 3896
rect 7708 3924 7714 3936
rect 7837 3927 7895 3933
rect 7837 3924 7849 3927
rect 7708 3896 7849 3924
rect 7708 3884 7714 3896
rect 7837 3893 7849 3896
rect 7883 3924 7895 3927
rect 8018 3924 8024 3936
rect 7883 3896 8024 3924
rect 7883 3893 7895 3896
rect 7837 3887 7895 3893
rect 8018 3884 8024 3896
rect 8076 3924 8082 3936
rect 8220 3933 8248 3964
rect 9140 3936 9168 4032
rect 9950 4020 9956 4032
rect 10008 4020 10014 4072
rect 10410 4060 10416 4072
rect 10371 4032 10416 4060
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 12342 4020 12348 4072
rect 12400 4060 12406 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12400 4032 12449 4060
rect 12400 4020 12406 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 12618 4020 12624 4072
rect 12676 4060 12682 4072
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12676 4032 12909 4060
rect 12676 4020 12682 4032
rect 12897 4029 12909 4032
rect 12943 4060 12955 4063
rect 13814 4060 13820 4072
rect 12943 4032 13820 4060
rect 12943 4029 12955 4032
rect 12897 4023 12955 4029
rect 13814 4020 13820 4032
rect 13872 4020 13878 4072
rect 14737 4063 14795 4069
rect 14737 4029 14749 4063
rect 14783 4060 14795 4063
rect 15102 4060 15108 4072
rect 14783 4032 15108 4060
rect 14783 4029 14795 4032
rect 14737 4023 14795 4029
rect 15102 4020 15108 4032
rect 15160 4060 15166 4072
rect 15488 4060 15516 4168
rect 16669 4165 16681 4199
rect 16715 4196 16727 4199
rect 16850 4196 16856 4208
rect 16715 4168 16749 4196
rect 16811 4168 16856 4196
rect 16715 4165 16727 4168
rect 16669 4159 16727 4165
rect 15565 4131 15623 4137
rect 15565 4097 15577 4131
rect 15611 4128 15623 4131
rect 15746 4128 15752 4140
rect 15611 4100 15752 4128
rect 15611 4097 15623 4100
rect 15565 4091 15623 4097
rect 15746 4088 15752 4100
rect 15804 4128 15810 4140
rect 16206 4128 16212 4140
rect 15804 4100 16212 4128
rect 15804 4088 15810 4100
rect 16206 4088 16212 4100
rect 16264 4128 16270 4140
rect 16684 4128 16712 4159
rect 16850 4156 16856 4168
rect 16908 4156 16914 4208
rect 16942 4156 16948 4208
rect 17000 4196 17006 4208
rect 17497 4199 17555 4205
rect 17497 4196 17509 4199
rect 17000 4168 17509 4196
rect 17000 4156 17006 4168
rect 17497 4165 17509 4168
rect 17543 4196 17555 4199
rect 18046 4196 18052 4208
rect 17543 4168 18052 4196
rect 17543 4165 17555 4168
rect 17497 4159 17555 4165
rect 18046 4156 18052 4168
rect 18104 4156 18110 4208
rect 18414 4156 18420 4208
rect 18472 4196 18478 4208
rect 18969 4199 19027 4205
rect 18969 4196 18981 4199
rect 18472 4168 18981 4196
rect 18472 4156 18478 4168
rect 18969 4165 18981 4168
rect 19015 4196 19027 4199
rect 19061 4199 19119 4205
rect 19061 4196 19073 4199
rect 19015 4168 19073 4196
rect 19015 4165 19027 4168
rect 18969 4159 19027 4165
rect 19061 4165 19073 4168
rect 19107 4165 19119 4199
rect 19061 4159 19119 4165
rect 16264 4100 16712 4128
rect 16264 4088 16270 4100
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 17865 4131 17923 4137
rect 16816 4100 16861 4128
rect 16816 4088 16822 4100
rect 17865 4097 17877 4131
rect 17911 4128 17923 4131
rect 19306 4128 19334 4236
rect 19886 4224 19892 4236
rect 19944 4224 19950 4276
rect 24026 4264 24032 4276
rect 23987 4236 24032 4264
rect 24026 4224 24032 4236
rect 24084 4224 24090 4276
rect 25409 4267 25467 4273
rect 25409 4233 25421 4267
rect 25455 4264 25467 4267
rect 26145 4267 26203 4273
rect 26145 4264 26157 4267
rect 25455 4236 26157 4264
rect 25455 4233 25467 4236
rect 25409 4227 25467 4233
rect 26145 4233 26157 4236
rect 26191 4264 26203 4267
rect 26418 4264 26424 4276
rect 26191 4236 26424 4264
rect 26191 4233 26203 4236
rect 26145 4227 26203 4233
rect 26418 4224 26424 4236
rect 26476 4264 26482 4276
rect 27154 4264 27160 4276
rect 26476 4236 27160 4264
rect 26476 4224 26482 4236
rect 27154 4224 27160 4236
rect 27212 4264 27218 4276
rect 27249 4267 27307 4273
rect 27249 4264 27261 4267
rect 27212 4236 27261 4264
rect 27212 4224 27218 4236
rect 27249 4233 27261 4236
rect 27295 4233 27307 4267
rect 29638 4264 29644 4276
rect 27249 4227 27307 4233
rect 27448 4236 29644 4264
rect 19426 4196 19432 4208
rect 19387 4168 19432 4196
rect 19426 4156 19432 4168
rect 19484 4196 19490 4208
rect 19751 4199 19809 4205
rect 19751 4196 19763 4199
rect 19484 4168 19763 4196
rect 19484 4156 19490 4168
rect 19751 4165 19763 4168
rect 19797 4165 19809 4199
rect 19751 4159 19809 4165
rect 24118 4156 24124 4208
rect 24176 4196 24182 4208
rect 27448 4196 27476 4236
rect 29638 4224 29644 4236
rect 29696 4264 29702 4276
rect 30193 4267 30251 4273
rect 30193 4264 30205 4267
rect 29696 4236 30205 4264
rect 29696 4224 29702 4236
rect 30193 4233 30205 4236
rect 30239 4264 30251 4267
rect 35434 4264 35440 4276
rect 30239 4236 35440 4264
rect 30239 4233 30251 4236
rect 30193 4227 30251 4233
rect 35434 4224 35440 4236
rect 35492 4224 35498 4276
rect 27706 4196 27712 4208
rect 24176 4168 27476 4196
rect 27667 4168 27712 4196
rect 24176 4156 24182 4168
rect 27706 4156 27712 4168
rect 27764 4196 27770 4208
rect 27985 4199 28043 4205
rect 27985 4196 27997 4199
rect 27764 4168 27997 4196
rect 27764 4156 27770 4168
rect 27985 4165 27997 4168
rect 28031 4165 28043 4199
rect 28258 4196 28264 4208
rect 28219 4168 28264 4196
rect 27985 4159 28043 4165
rect 28258 4156 28264 4168
rect 28316 4156 28322 4208
rect 19981 4131 20039 4137
rect 19981 4128 19993 4131
rect 17911 4100 19334 4128
rect 19628 4100 19993 4128
rect 17911 4097 17923 4100
rect 17865 4091 17923 4097
rect 18156 4072 18184 4100
rect 15160 4032 15516 4060
rect 16540 4063 16598 4069
rect 15160 4020 15166 4032
rect 16540 4029 16552 4063
rect 16586 4060 16598 4063
rect 17954 4060 17960 4072
rect 16586 4032 17960 4060
rect 16586 4029 16598 4032
rect 16540 4023 16598 4029
rect 17954 4020 17960 4032
rect 18012 4060 18018 4072
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 18012 4032 18061 4060
rect 18012 4020 18018 4032
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 18138 4020 18144 4072
rect 18196 4060 18202 4072
rect 18325 4063 18383 4069
rect 18196 4032 18241 4060
rect 18196 4020 18202 4032
rect 18325 4029 18337 4063
rect 18371 4060 18383 4063
rect 18414 4060 18420 4072
rect 18371 4032 18420 4060
rect 18371 4029 18383 4032
rect 18325 4023 18383 4029
rect 18414 4020 18420 4032
rect 18472 4020 18478 4072
rect 18969 4063 19027 4069
rect 18969 4029 18981 4063
rect 19015 4060 19027 4063
rect 19628 4060 19656 4100
rect 19981 4097 19993 4100
rect 20027 4097 20039 4131
rect 19981 4091 20039 4097
rect 21174 4088 21180 4140
rect 21232 4128 21238 4140
rect 21545 4131 21603 4137
rect 21545 4128 21557 4131
rect 21232 4100 21557 4128
rect 21232 4088 21238 4100
rect 21545 4097 21557 4100
rect 21591 4128 21603 4131
rect 21591 4100 21956 4128
rect 21591 4097 21603 4100
rect 21545 4091 21603 4097
rect 21928 4072 21956 4100
rect 22186 4088 22192 4140
rect 22244 4128 22250 4140
rect 22646 4128 22652 4140
rect 22244 4100 22652 4128
rect 22244 4088 22250 4100
rect 22646 4088 22652 4100
rect 22704 4128 22710 4140
rect 23382 4128 23388 4140
rect 22704 4100 23388 4128
rect 22704 4088 22710 4100
rect 23382 4088 23388 4100
rect 23440 4088 23446 4140
rect 25038 4088 25044 4140
rect 25096 4128 25102 4140
rect 25682 4128 25688 4140
rect 25096 4100 25688 4128
rect 25096 4088 25102 4100
rect 25682 4088 25688 4100
rect 25740 4088 25746 4140
rect 28166 4088 28172 4140
rect 28224 4128 28230 4140
rect 29411 4131 29469 4137
rect 29411 4128 29423 4131
rect 28224 4100 29423 4128
rect 28224 4088 28230 4100
rect 29411 4097 29423 4100
rect 29457 4097 29469 4131
rect 29822 4128 29828 4140
rect 29783 4100 29828 4128
rect 29411 4091 29469 4097
rect 29822 4088 29828 4100
rect 29880 4088 29886 4140
rect 21910 4060 21916 4072
rect 19015 4032 19656 4060
rect 21100 4032 21588 4060
rect 21871 4032 21916 4060
rect 19015 4029 19027 4032
rect 18969 4023 19027 4029
rect 9398 3952 9404 4004
rect 9456 3992 9462 4004
rect 9766 3992 9772 4004
rect 9456 3964 9772 3992
rect 9456 3952 9462 3964
rect 9766 3952 9772 3964
rect 9824 3992 9830 4004
rect 11333 3995 11391 4001
rect 11333 3992 11345 3995
rect 9824 3964 11345 3992
rect 9824 3952 9830 3964
rect 11333 3961 11345 3964
rect 11379 3961 11391 3995
rect 11333 3955 11391 3961
rect 16393 3995 16451 4001
rect 16393 3961 16405 3995
rect 16439 3992 16451 3995
rect 16666 3992 16672 4004
rect 16439 3964 16672 3992
rect 16439 3961 16451 3964
rect 16393 3955 16451 3961
rect 16666 3952 16672 3964
rect 16724 3952 16730 4004
rect 19426 3992 19432 4004
rect 18064 3964 19432 3992
rect 18064 3936 18092 3964
rect 19426 3952 19432 3964
rect 19484 3952 19490 4004
rect 19613 3995 19671 4001
rect 19613 3961 19625 3995
rect 19659 3992 19671 3995
rect 20622 3992 20628 4004
rect 19659 3964 20628 3992
rect 19659 3961 19671 3964
rect 19613 3955 19671 3961
rect 20622 3952 20628 3964
rect 20680 3952 20686 4004
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 8076 3896 8217 3924
rect 8076 3884 8082 3896
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 8846 3924 8852 3936
rect 8807 3896 8852 3924
rect 8205 3887 8263 3893
rect 8846 3884 8852 3896
rect 8904 3884 8910 3936
rect 9122 3884 9128 3936
rect 9180 3884 9186 3936
rect 9858 3884 9864 3936
rect 9916 3924 9922 3936
rect 11057 3927 11115 3933
rect 11057 3924 11069 3927
rect 9916 3896 11069 3924
rect 9916 3884 9922 3896
rect 11057 3893 11069 3896
rect 11103 3924 11115 3927
rect 11698 3924 11704 3936
rect 11103 3896 11704 3924
rect 11103 3893 11115 3896
rect 11057 3887 11115 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 15194 3884 15200 3936
rect 15252 3924 15258 3936
rect 15841 3927 15899 3933
rect 15841 3924 15853 3927
rect 15252 3896 15853 3924
rect 15252 3884 15258 3896
rect 15841 3893 15853 3896
rect 15887 3924 15899 3927
rect 16758 3924 16764 3936
rect 15887 3896 16764 3924
rect 15887 3893 15899 3896
rect 15841 3887 15899 3893
rect 16758 3884 16764 3896
rect 16816 3884 16822 3936
rect 18046 3884 18052 3936
rect 18104 3884 18110 3936
rect 18509 3927 18567 3933
rect 18509 3893 18521 3927
rect 18555 3924 18567 3927
rect 18782 3924 18788 3936
rect 18555 3896 18788 3924
rect 18555 3893 18567 3896
rect 18509 3887 18567 3893
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 19150 3884 19156 3936
rect 19208 3924 19214 3936
rect 20257 3927 20315 3933
rect 20257 3924 20269 3927
rect 19208 3896 20269 3924
rect 19208 3884 19214 3896
rect 20257 3893 20269 3896
rect 20303 3893 20315 3927
rect 20257 3887 20315 3893
rect 20806 3884 20812 3936
rect 20864 3924 20870 3936
rect 21100 3933 21128 4032
rect 21560 3992 21588 4032
rect 21910 4020 21916 4032
rect 21968 4020 21974 4072
rect 22094 4060 22100 4072
rect 22055 4032 22100 4060
rect 22094 4020 22100 4032
rect 22152 4060 22158 4072
rect 22370 4060 22376 4072
rect 22152 4032 22376 4060
rect 22152 4020 22158 4032
rect 22370 4020 22376 4032
rect 22428 4020 22434 4072
rect 22465 4063 22523 4069
rect 22465 4029 22477 4063
rect 22511 4029 22523 4063
rect 24486 4060 24492 4072
rect 24447 4032 24492 4060
rect 22465 4023 22523 4029
rect 22480 3992 22508 4023
rect 24486 4020 24492 4032
rect 24544 4020 24550 4072
rect 27801 4063 27859 4069
rect 27801 4029 27813 4063
rect 27847 4029 27859 4063
rect 27801 4023 27859 4029
rect 22922 3992 22928 4004
rect 21560 3964 22928 3992
rect 22922 3952 22928 3964
rect 22980 3992 22986 4004
rect 23017 3995 23075 4001
rect 23017 3992 23029 3995
rect 22980 3964 23029 3992
rect 22980 3952 22986 3964
rect 23017 3961 23029 3964
rect 23063 3961 23075 3995
rect 23017 3955 23075 3961
rect 23750 3952 23756 4004
rect 23808 3992 23814 4004
rect 24397 3995 24455 4001
rect 24397 3992 24409 3995
rect 23808 3964 24409 3992
rect 23808 3952 23814 3964
rect 24397 3961 24409 3964
rect 24443 3992 24455 3995
rect 24851 3995 24909 4001
rect 24851 3992 24863 3995
rect 24443 3964 24863 3992
rect 24443 3961 24455 3964
rect 24397 3955 24455 3961
rect 24851 3961 24863 3964
rect 24897 3992 24909 3995
rect 24946 3992 24952 4004
rect 24897 3964 24952 3992
rect 24897 3961 24909 3964
rect 24851 3955 24909 3961
rect 24946 3952 24952 3964
rect 25004 3952 25010 4004
rect 26326 3992 26332 4004
rect 26287 3964 26332 3992
rect 26326 3952 26332 3964
rect 26384 3952 26390 4004
rect 26418 3952 26424 4004
rect 26476 3992 26482 4004
rect 26970 3992 26976 4004
rect 26476 3964 26521 3992
rect 26931 3964 26976 3992
rect 26476 3952 26482 3964
rect 26970 3952 26976 3964
rect 27028 3952 27034 4004
rect 27816 3992 27844 4023
rect 28534 4020 28540 4072
rect 28592 4060 28598 4072
rect 29324 4063 29382 4069
rect 29324 4060 29336 4063
rect 28592 4032 29336 4060
rect 28592 4020 28598 4032
rect 29324 4029 29336 4032
rect 29370 4060 29382 4063
rect 29840 4060 29868 4088
rect 30282 4060 30288 4072
rect 29370 4032 29868 4060
rect 30243 4032 30288 4060
rect 29370 4029 29382 4032
rect 29324 4023 29382 4029
rect 30282 4020 30288 4032
rect 30340 4060 30346 4072
rect 30745 4063 30803 4069
rect 30745 4060 30757 4063
rect 30340 4032 30757 4060
rect 30340 4020 30346 4032
rect 30745 4029 30757 4032
rect 30791 4029 30803 4063
rect 30745 4023 30803 4029
rect 28629 3995 28687 4001
rect 28629 3992 28641 3995
rect 27816 3964 28641 3992
rect 21085 3927 21143 3933
rect 21085 3924 21097 3927
rect 20864 3896 21097 3924
rect 20864 3884 20870 3896
rect 21085 3893 21097 3896
rect 21131 3893 21143 3927
rect 22738 3924 22744 3936
rect 22699 3896 22744 3924
rect 21085 3887 21143 3893
rect 22738 3884 22744 3896
rect 22796 3884 22802 3936
rect 25498 3884 25504 3936
rect 25556 3924 25562 3936
rect 27816 3924 27844 3964
rect 28629 3961 28641 3964
rect 28675 3961 28687 3995
rect 28629 3955 28687 3961
rect 30466 3924 30472 3936
rect 25556 3896 27844 3924
rect 30427 3896 30472 3924
rect 25556 3884 25562 3896
rect 30466 3884 30472 3896
rect 30524 3884 30530 3936
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 1762 3720 1768 3732
rect 1723 3692 1768 3720
rect 1762 3680 1768 3692
rect 1820 3680 1826 3732
rect 1946 3680 1952 3732
rect 2004 3720 2010 3732
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 2004 3692 2697 3720
rect 2004 3680 2010 3692
rect 2685 3689 2697 3692
rect 2731 3689 2743 3723
rect 2685 3683 2743 3689
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 3053 3723 3111 3729
rect 3053 3720 3065 3723
rect 3016 3692 3065 3720
rect 3016 3680 3022 3692
rect 3053 3689 3065 3692
rect 3099 3689 3111 3723
rect 3053 3683 3111 3689
rect 4203 3723 4261 3729
rect 4203 3689 4215 3723
rect 4249 3720 4261 3723
rect 5442 3720 5448 3732
rect 4249 3692 5448 3720
rect 4249 3689 4261 3692
rect 4203 3683 4261 3689
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 5810 3720 5816 3732
rect 5771 3692 5816 3720
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 6549 3723 6607 3729
rect 6549 3720 6561 3723
rect 5920 3692 6561 3720
rect 3786 3612 3792 3664
rect 3844 3652 3850 3664
rect 5215 3655 5273 3661
rect 5215 3652 5227 3655
rect 3844 3624 5227 3652
rect 3844 3612 3850 3624
rect 5215 3621 5227 3624
rect 5261 3621 5273 3655
rect 5920 3652 5948 3692
rect 6549 3689 6561 3692
rect 6595 3720 6607 3723
rect 8202 3720 8208 3732
rect 6595 3692 8208 3720
rect 6595 3689 6607 3692
rect 6549 3683 6607 3689
rect 8202 3680 8208 3692
rect 8260 3720 8266 3732
rect 9214 3720 9220 3732
rect 8260 3692 9220 3720
rect 8260 3680 8266 3692
rect 9214 3680 9220 3692
rect 9272 3680 9278 3732
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 9769 3723 9827 3729
rect 9769 3720 9781 3723
rect 9732 3692 9781 3720
rect 9732 3680 9738 3692
rect 9769 3689 9781 3692
rect 9815 3689 9827 3723
rect 9769 3683 9827 3689
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 10008 3692 10701 3720
rect 10008 3680 10014 3692
rect 10689 3689 10701 3692
rect 10735 3720 10747 3723
rect 12434 3720 12440 3732
rect 10735 3692 12440 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 12618 3720 12624 3732
rect 12579 3692 12624 3720
rect 12618 3680 12624 3692
rect 12676 3680 12682 3732
rect 15930 3720 15936 3732
rect 15891 3692 15936 3720
rect 15930 3680 15936 3692
rect 15988 3720 15994 3732
rect 16945 3723 17003 3729
rect 16945 3720 16957 3723
rect 15988 3692 16957 3720
rect 15988 3680 15994 3692
rect 16945 3689 16957 3692
rect 16991 3689 17003 3723
rect 17586 3720 17592 3732
rect 17547 3692 17592 3720
rect 16945 3683 17003 3689
rect 17586 3680 17592 3692
rect 17644 3680 17650 3732
rect 20622 3720 20628 3732
rect 17880 3692 20484 3720
rect 20583 3692 20628 3720
rect 8846 3652 8852 3664
rect 5215 3615 5273 3621
rect 5368 3624 5948 3652
rect 6380 3624 8852 3652
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3584 2007 3587
rect 2130 3584 2136 3596
rect 1995 3556 2136 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 2130 3544 2136 3556
rect 2188 3544 2194 3596
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3553 2283 3587
rect 2225 3547 2283 3553
rect 4132 3587 4190 3593
rect 4132 3553 4144 3587
rect 4178 3584 4190 3587
rect 4246 3584 4252 3596
rect 4178 3556 4252 3584
rect 4178 3553 4190 3556
rect 4132 3547 4190 3553
rect 2240 3516 2268 3547
rect 4246 3544 4252 3556
rect 4304 3544 4310 3596
rect 5074 3584 5080 3596
rect 5035 3556 5080 3584
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 5368 3584 5396 3624
rect 5184 3556 5396 3584
rect 3513 3519 3571 3525
rect 3513 3516 3525 3519
rect 2240 3488 3525 3516
rect 3513 3485 3525 3488
rect 3559 3516 3571 3519
rect 3694 3516 3700 3528
rect 3559 3488 3700 3516
rect 3559 3485 3571 3488
rect 3513 3479 3571 3485
rect 3694 3476 3700 3488
rect 3752 3516 3758 3528
rect 5184 3516 5212 3556
rect 5626 3544 5632 3596
rect 5684 3584 5690 3596
rect 6380 3593 6408 3624
rect 8846 3612 8852 3624
rect 8904 3612 8910 3664
rect 12636 3652 12664 3680
rect 14826 3652 14832 3664
rect 10244 3624 12664 3652
rect 14016 3624 14832 3652
rect 10244 3596 10272 3624
rect 6365 3587 6423 3593
rect 6365 3584 6377 3587
rect 5684 3556 6377 3584
rect 5684 3544 5690 3556
rect 6365 3553 6377 3556
rect 6411 3553 6423 3587
rect 7374 3584 7380 3596
rect 6365 3547 6423 3553
rect 6840 3556 7380 3584
rect 3752 3488 5212 3516
rect 3752 3476 3758 3488
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 6178 3516 6184 3528
rect 5316 3488 6184 3516
rect 5316 3476 5322 3488
rect 6178 3476 6184 3488
rect 6236 3516 6242 3528
rect 6840 3516 6868 3556
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 7650 3584 7656 3596
rect 7611 3556 7656 3584
rect 7650 3544 7656 3556
rect 7708 3544 7714 3596
rect 7760 3556 8524 3584
rect 7466 3516 7472 3528
rect 6236 3488 6868 3516
rect 7379 3488 7472 3516
rect 6236 3476 6242 3488
rect 7466 3476 7472 3488
rect 7524 3516 7530 3528
rect 7760 3516 7788 3556
rect 8496 3528 8524 3556
rect 9030 3544 9036 3596
rect 9088 3584 9094 3596
rect 9950 3584 9956 3596
rect 9088 3556 9956 3584
rect 9088 3544 9094 3556
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 10226 3584 10232 3596
rect 10139 3556 10232 3584
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 11974 3584 11980 3596
rect 11935 3556 11980 3584
rect 11974 3544 11980 3556
rect 12032 3544 12038 3596
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 12897 3587 12955 3593
rect 12897 3584 12909 3587
rect 12492 3556 12909 3584
rect 12492 3544 12498 3556
rect 12897 3553 12909 3556
rect 12943 3553 12955 3587
rect 12897 3547 12955 3553
rect 13814 3544 13820 3596
rect 13872 3584 13878 3596
rect 14016 3593 14044 3624
rect 14826 3612 14832 3624
rect 14884 3652 14890 3664
rect 15565 3655 15623 3661
rect 15565 3652 15577 3655
rect 14884 3624 15577 3652
rect 14884 3612 14890 3624
rect 15565 3621 15577 3624
rect 15611 3652 15623 3655
rect 17770 3652 17776 3664
rect 15611 3624 17776 3652
rect 15611 3621 15623 3624
rect 15565 3615 15623 3621
rect 17770 3612 17776 3624
rect 17828 3612 17834 3664
rect 14001 3587 14059 3593
rect 13872 3556 13917 3584
rect 13872 3544 13878 3556
rect 14001 3553 14013 3587
rect 14047 3553 14059 3587
rect 14366 3584 14372 3596
rect 14327 3556 14372 3584
rect 14001 3547 14059 3553
rect 14366 3544 14372 3556
rect 14424 3544 14430 3596
rect 16390 3584 16396 3596
rect 16351 3556 16396 3584
rect 16390 3544 16396 3556
rect 16448 3544 16454 3596
rect 16945 3587 17003 3593
rect 16945 3553 16957 3587
rect 16991 3584 17003 3587
rect 17880 3584 17908 3692
rect 18509 3655 18567 3661
rect 18509 3621 18521 3655
rect 18555 3652 18567 3655
rect 18690 3652 18696 3664
rect 18555 3624 18696 3652
rect 18555 3621 18567 3624
rect 18509 3615 18567 3621
rect 18690 3612 18696 3624
rect 18748 3612 18754 3664
rect 18874 3612 18880 3664
rect 18932 3652 18938 3664
rect 19337 3655 19395 3661
rect 19337 3652 19349 3655
rect 18932 3624 19349 3652
rect 18932 3612 18938 3624
rect 19337 3621 19349 3624
rect 19383 3652 19395 3655
rect 20254 3652 20260 3664
rect 19383 3624 20260 3652
rect 19383 3621 19395 3624
rect 19337 3615 19395 3621
rect 20254 3612 20260 3624
rect 20312 3612 20318 3664
rect 18785 3587 18843 3593
rect 18785 3584 18797 3587
rect 16991 3556 17908 3584
rect 17972 3556 18797 3584
rect 16991 3553 17003 3556
rect 16945 3547 17003 3553
rect 17972 3528 18000 3556
rect 18785 3553 18797 3556
rect 18831 3553 18843 3587
rect 18785 3547 18843 3553
rect 19242 3544 19248 3596
rect 19300 3584 19306 3596
rect 19521 3587 19579 3593
rect 19521 3584 19533 3587
rect 19300 3556 19533 3584
rect 19300 3544 19306 3556
rect 19521 3553 19533 3556
rect 19567 3553 19579 3587
rect 20456 3584 20484 3692
rect 20622 3680 20628 3692
rect 20680 3680 20686 3732
rect 22646 3720 22652 3732
rect 22607 3692 22652 3720
rect 22646 3680 22652 3692
rect 22704 3680 22710 3732
rect 23937 3723 23995 3729
rect 23937 3689 23949 3723
rect 23983 3720 23995 3723
rect 24486 3720 24492 3732
rect 23983 3692 24492 3720
rect 23983 3689 23995 3692
rect 23937 3683 23995 3689
rect 24486 3680 24492 3692
rect 24544 3680 24550 3732
rect 28629 3723 28687 3729
rect 28629 3689 28641 3723
rect 28675 3720 28687 3723
rect 29086 3720 29092 3732
rect 28675 3692 29092 3720
rect 28675 3689 28687 3692
rect 28629 3683 28687 3689
rect 29086 3680 29092 3692
rect 29144 3720 29150 3732
rect 29144 3692 29684 3720
rect 29144 3680 29150 3692
rect 20640 3652 20668 3680
rect 22094 3652 22100 3664
rect 20640 3624 22100 3652
rect 21174 3584 21180 3596
rect 20456 3556 21180 3584
rect 19521 3547 19579 3553
rect 21174 3544 21180 3556
rect 21232 3544 21238 3596
rect 21376 3593 21404 3624
rect 22094 3612 22100 3624
rect 22152 3652 22158 3664
rect 22281 3655 22339 3661
rect 22281 3652 22293 3655
rect 22152 3624 22293 3652
rect 22152 3612 22158 3624
rect 22281 3621 22293 3624
rect 22327 3621 22339 3655
rect 22281 3615 22339 3621
rect 21361 3587 21419 3593
rect 21361 3553 21373 3587
rect 21407 3553 21419 3587
rect 21361 3547 21419 3553
rect 21729 3587 21787 3593
rect 21729 3553 21741 3587
rect 21775 3584 21787 3587
rect 22554 3584 22560 3596
rect 21775 3556 22560 3584
rect 21775 3553 21787 3556
rect 21729 3547 21787 3553
rect 8110 3516 8116 3528
rect 7524 3488 7788 3516
rect 8071 3488 8116 3516
rect 7524 3476 7530 3488
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 8478 3516 8484 3528
rect 8391 3488 8484 3516
rect 8478 3476 8484 3488
rect 8536 3516 8542 3528
rect 9858 3516 9864 3528
rect 8536 3488 9864 3516
rect 8536 3476 8542 3488
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3516 12311 3519
rect 12342 3516 12348 3528
rect 12299 3488 12348 3516
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 17954 3525 17960 3528
rect 16761 3519 16819 3525
rect 16761 3485 16773 3519
rect 16807 3516 16819 3519
rect 17037 3519 17095 3525
rect 17037 3516 17049 3519
rect 16807 3488 17049 3516
rect 16807 3485 16819 3488
rect 16761 3479 16819 3485
rect 17037 3485 17049 3488
rect 17083 3516 17095 3519
rect 17920 3519 17960 3525
rect 17920 3516 17932 3519
rect 17083 3488 17932 3516
rect 17083 3485 17095 3488
rect 17037 3479 17095 3485
rect 17920 3485 17932 3488
rect 17920 3479 17960 3485
rect 17954 3476 17960 3479
rect 18012 3476 18018 3528
rect 18141 3519 18199 3525
rect 18141 3485 18153 3519
rect 18187 3516 18199 3519
rect 18414 3516 18420 3528
rect 18187 3488 18420 3516
rect 18187 3485 18199 3488
rect 18141 3479 18199 3485
rect 18414 3476 18420 3488
rect 18472 3476 18478 3528
rect 19886 3516 19892 3528
rect 19847 3488 19892 3516
rect 19886 3476 19892 3488
rect 19944 3476 19950 3528
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 21744 3516 21772 3547
rect 22554 3544 22560 3556
rect 22612 3544 22618 3596
rect 22664 3584 22692 3680
rect 24213 3655 24271 3661
rect 24213 3652 24225 3655
rect 22940 3624 24225 3652
rect 22833 3587 22891 3593
rect 22833 3584 22845 3587
rect 22664 3556 22845 3584
rect 22833 3553 22845 3556
rect 22879 3553 22891 3587
rect 22833 3547 22891 3553
rect 20680 3488 21772 3516
rect 20680 3476 20686 3488
rect 21818 3476 21824 3528
rect 21876 3516 21882 3528
rect 22005 3519 22063 3525
rect 22005 3516 22017 3519
rect 21876 3488 22017 3516
rect 21876 3476 21882 3488
rect 22005 3485 22017 3488
rect 22051 3516 22063 3519
rect 22940 3516 22968 3624
rect 24213 3621 24225 3624
rect 24259 3621 24271 3655
rect 24213 3615 24271 3621
rect 24946 3612 24952 3664
rect 25004 3652 25010 3664
rect 28071 3655 28129 3661
rect 28071 3652 28083 3655
rect 25004 3624 28083 3652
rect 25004 3612 25010 3624
rect 28071 3621 28083 3624
rect 28117 3652 28129 3655
rect 28442 3652 28448 3664
rect 28117 3624 28448 3652
rect 28117 3621 28129 3624
rect 28071 3615 28129 3621
rect 28442 3612 28448 3624
rect 28500 3612 28506 3664
rect 29656 3661 29684 3692
rect 29641 3655 29699 3661
rect 29641 3621 29653 3655
rect 29687 3621 29699 3655
rect 29641 3615 29699 3621
rect 23658 3584 23664 3596
rect 23619 3556 23664 3584
rect 23658 3544 23664 3556
rect 23716 3544 23722 3596
rect 24854 3584 24860 3596
rect 24815 3556 24860 3584
rect 24854 3544 24860 3556
rect 24912 3544 24918 3596
rect 26142 3544 26148 3596
rect 26200 3584 26206 3596
rect 26548 3587 26606 3593
rect 26548 3584 26560 3587
rect 26200 3556 26560 3584
rect 26200 3544 26206 3556
rect 26548 3553 26560 3556
rect 26594 3584 26606 3587
rect 27246 3584 27252 3596
rect 26594 3556 27252 3584
rect 26594 3553 26606 3556
rect 26548 3547 26606 3553
rect 27246 3544 27252 3556
rect 27304 3544 27310 3596
rect 27522 3544 27528 3596
rect 27580 3584 27586 3596
rect 27709 3587 27767 3593
rect 27709 3584 27721 3587
rect 27580 3556 27721 3584
rect 27580 3544 27586 3556
rect 27709 3553 27721 3556
rect 27755 3553 27767 3587
rect 27709 3547 27767 3553
rect 23753 3519 23811 3525
rect 23753 3516 23765 3519
rect 22051 3488 22968 3516
rect 23216 3488 23765 3516
rect 22051 3485 22063 3488
rect 22005 3479 22063 3485
rect 16206 3408 16212 3460
rect 16264 3448 16270 3460
rect 18046 3448 18052 3460
rect 16264 3420 18052 3448
rect 16264 3408 16270 3420
rect 18046 3408 18052 3420
rect 18104 3408 18110 3460
rect 18322 3408 18328 3460
rect 18380 3448 18386 3460
rect 20165 3451 20223 3457
rect 20165 3448 20177 3451
rect 18380 3420 20177 3448
rect 18380 3408 18386 3420
rect 20165 3417 20177 3420
rect 20211 3417 20223 3451
rect 20165 3411 20223 3417
rect 22094 3408 22100 3460
rect 22152 3448 22158 3460
rect 23216 3448 23244 3488
rect 23753 3485 23765 3488
rect 23799 3516 23811 3519
rect 23799 3488 24532 3516
rect 23799 3485 23811 3488
rect 23753 3479 23811 3485
rect 22152 3420 23244 3448
rect 24504 3448 24532 3488
rect 26970 3476 26976 3528
rect 27028 3516 27034 3528
rect 29549 3519 29607 3525
rect 29549 3516 29561 3519
rect 27028 3488 29561 3516
rect 27028 3476 27034 3488
rect 29549 3485 29561 3488
rect 29595 3516 29607 3519
rect 30742 3516 30748 3528
rect 29595 3488 30748 3516
rect 29595 3485 29607 3488
rect 29549 3479 29607 3485
rect 30742 3476 30748 3488
rect 30800 3476 30806 3528
rect 27982 3448 27988 3460
rect 24504 3420 27988 3448
rect 22152 3408 22158 3420
rect 27982 3408 27988 3420
rect 28040 3408 28046 3460
rect 30098 3448 30104 3460
rect 30059 3420 30104 3448
rect 30098 3408 30104 3420
rect 30156 3408 30162 3460
rect 7190 3380 7196 3392
rect 7151 3352 7196 3380
rect 7190 3340 7196 3352
rect 7248 3340 7254 3392
rect 14921 3383 14979 3389
rect 14921 3349 14933 3383
rect 14967 3380 14979 3383
rect 15194 3380 15200 3392
rect 14967 3352 15200 3380
rect 14967 3349 14979 3352
rect 14921 3343 14979 3349
rect 15194 3340 15200 3352
rect 15252 3340 15258 3392
rect 18064 3380 18092 3408
rect 19153 3383 19211 3389
rect 19153 3380 19165 3383
rect 18064 3352 19165 3380
rect 19153 3349 19165 3352
rect 19199 3349 19211 3383
rect 24578 3380 24584 3392
rect 24539 3352 24584 3380
rect 19153 3343 19211 3349
rect 24578 3340 24584 3352
rect 24636 3340 24642 3392
rect 25222 3380 25228 3392
rect 25183 3352 25228 3380
rect 25222 3340 25228 3352
rect 25280 3340 25286 3392
rect 26234 3380 26240 3392
rect 26195 3352 26240 3380
rect 26234 3340 26240 3352
rect 26292 3340 26298 3392
rect 26326 3340 26332 3392
rect 26384 3380 26390 3392
rect 26651 3383 26709 3389
rect 26651 3380 26663 3383
rect 26384 3352 26663 3380
rect 26384 3340 26390 3352
rect 26651 3349 26663 3352
rect 26697 3380 26709 3383
rect 26973 3383 27031 3389
rect 26973 3380 26985 3383
rect 26697 3352 26985 3380
rect 26697 3349 26709 3352
rect 26651 3343 26709 3349
rect 26973 3349 26985 3352
rect 27019 3349 27031 3383
rect 26973 3343 27031 3349
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 1765 3179 1823 3185
rect 1765 3145 1777 3179
rect 1811 3176 1823 3179
rect 2130 3176 2136 3188
rect 1811 3148 2136 3176
rect 1811 3145 1823 3148
rect 1765 3139 1823 3145
rect 2130 3136 2136 3148
rect 2188 3136 2194 3188
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 3835 3179 3893 3185
rect 3835 3176 3847 3179
rect 3292 3148 3847 3176
rect 3292 3136 3298 3148
rect 3835 3145 3847 3148
rect 3881 3145 3893 3179
rect 3835 3139 3893 3145
rect 4617 3179 4675 3185
rect 4617 3145 4629 3179
rect 4663 3176 4675 3179
rect 4706 3176 4712 3188
rect 4663 3148 4712 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 3421 3111 3479 3117
rect 3421 3077 3433 3111
rect 3467 3108 3479 3111
rect 3694 3108 3700 3120
rect 3467 3080 3700 3108
rect 3467 3077 3479 3080
rect 3421 3071 3479 3077
rect 3694 3068 3700 3080
rect 3752 3068 3758 3120
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 2682 3040 2688 3052
rect 1544 3012 2452 3040
rect 2643 3012 2688 3040
rect 1544 3000 1550 3012
rect 2130 2972 2136 2984
rect 2091 2944 2136 2972
rect 2130 2932 2136 2944
rect 2188 2932 2194 2984
rect 2424 2981 2452 3012
rect 2682 3000 2688 3012
rect 2740 3000 2746 3052
rect 4522 3040 4528 3052
rect 2976 3012 4528 3040
rect 2976 2981 3004 3012
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2972 2467 2975
rect 2961 2975 3019 2981
rect 2961 2972 2973 2975
rect 2455 2944 2973 2972
rect 2455 2941 2467 2944
rect 2409 2935 2467 2941
rect 2961 2941 2973 2944
rect 3007 2941 3019 2975
rect 2961 2935 3019 2941
rect 3764 2975 3822 2981
rect 3764 2941 3776 2975
rect 3810 2972 3822 2975
rect 4632 2972 4660 3139
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 5074 3176 5080 3188
rect 5035 3148 5080 3176
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 5626 3176 5632 3188
rect 5587 3148 5632 3176
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 5905 3179 5963 3185
rect 5905 3145 5917 3179
rect 5951 3176 5963 3179
rect 5994 3176 6000 3188
rect 5951 3148 6000 3176
rect 5951 3145 5963 3148
rect 5905 3139 5963 3145
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 7374 3176 7380 3188
rect 7335 3148 7380 3176
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 8757 3179 8815 3185
rect 8757 3145 8769 3179
rect 8803 3176 8815 3179
rect 9398 3176 9404 3188
rect 8803 3148 9404 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 6641 3111 6699 3117
rect 6641 3077 6653 3111
rect 6687 3108 6699 3111
rect 7466 3108 7472 3120
rect 6687 3080 7472 3108
rect 6687 3077 6699 3080
rect 6641 3071 6699 3077
rect 7466 3068 7472 3080
rect 7524 3108 7530 3120
rect 7745 3111 7803 3117
rect 7745 3108 7757 3111
rect 7524 3080 7757 3108
rect 7524 3068 7530 3080
rect 7745 3077 7757 3080
rect 7791 3077 7803 3111
rect 7745 3071 7803 3077
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 6512 3012 8125 3040
rect 6512 3000 6518 3012
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 3810 2944 4660 2972
rect 5721 2975 5779 2981
rect 3810 2941 3822 2944
rect 3764 2935 3822 2941
rect 5721 2941 5733 2975
rect 5767 2972 5779 2975
rect 6270 2972 6276 2984
rect 5767 2944 6276 2972
rect 5767 2941 5779 2944
rect 5721 2935 5779 2941
rect 6270 2932 6276 2944
rect 6328 2932 6334 2984
rect 7190 2932 7196 2984
rect 7248 2972 7254 2984
rect 7653 2975 7711 2981
rect 7653 2972 7665 2975
rect 7248 2944 7665 2972
rect 7248 2932 7254 2944
rect 7653 2941 7665 2944
rect 7699 2941 7711 2975
rect 7653 2935 7711 2941
rect 4338 2864 4344 2916
rect 4396 2904 4402 2916
rect 7668 2904 7696 2935
rect 7834 2932 7840 2984
rect 7892 2972 7898 2984
rect 7929 2975 7987 2981
rect 7929 2972 7941 2975
rect 7892 2944 7941 2972
rect 7892 2932 7898 2944
rect 7929 2941 7941 2944
rect 7975 2972 7987 2975
rect 8772 2972 8800 3139
rect 9398 3136 9404 3148
rect 9456 3136 9462 3188
rect 9950 3136 9956 3188
rect 10008 3176 10014 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 10008 3148 10609 3176
rect 10008 3136 10014 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 11471 3179 11529 3185
rect 11471 3145 11483 3179
rect 11517 3176 11529 3179
rect 13078 3176 13084 3188
rect 11517 3148 13084 3176
rect 11517 3145 11529 3148
rect 11471 3139 11529 3145
rect 13078 3136 13084 3148
rect 13136 3136 13142 3188
rect 13403 3179 13461 3185
rect 13403 3145 13415 3179
rect 13449 3176 13461 3179
rect 13998 3176 14004 3188
rect 13449 3148 14004 3176
rect 13449 3145 13461 3148
rect 13403 3139 13461 3145
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 15473 3179 15531 3185
rect 15473 3145 15485 3179
rect 15519 3176 15531 3179
rect 15654 3176 15660 3188
rect 15519 3148 15660 3176
rect 15519 3145 15531 3148
rect 15473 3139 15531 3145
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 17497 3179 17555 3185
rect 17497 3145 17509 3179
rect 17543 3176 17555 3179
rect 17770 3176 17776 3188
rect 17543 3148 17776 3176
rect 17543 3145 17555 3148
rect 17497 3139 17555 3145
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 18230 3176 18236 3188
rect 18191 3148 18236 3176
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 22925 3179 22983 3185
rect 22925 3145 22937 3179
rect 22971 3176 22983 3179
rect 23658 3176 23664 3188
rect 22971 3148 23664 3176
rect 22971 3145 22983 3148
rect 22925 3139 22983 3145
rect 23658 3136 23664 3148
rect 23716 3136 23722 3188
rect 27246 3176 27252 3188
rect 27207 3148 27252 3176
rect 27246 3136 27252 3148
rect 27304 3136 27310 3188
rect 27522 3136 27528 3188
rect 27580 3176 27586 3188
rect 27617 3179 27675 3185
rect 27617 3176 27629 3179
rect 27580 3148 27629 3176
rect 27580 3136 27586 3148
rect 27617 3145 27629 3148
rect 27663 3145 27675 3179
rect 27982 3176 27988 3188
rect 27943 3148 27988 3176
rect 27617 3139 27675 3145
rect 27982 3136 27988 3148
rect 28040 3136 28046 3188
rect 30742 3176 30748 3188
rect 30703 3148 30748 3176
rect 30742 3136 30748 3148
rect 30800 3136 30806 3188
rect 10226 3108 10232 3120
rect 10187 3080 10232 3108
rect 10226 3068 10232 3080
rect 10284 3068 10290 3120
rect 15102 3108 15108 3120
rect 15063 3080 15108 3108
rect 15102 3068 15108 3080
rect 15160 3068 15166 3120
rect 16206 3068 16212 3120
rect 16264 3108 16270 3120
rect 16485 3111 16543 3117
rect 16485 3108 16497 3111
rect 16264 3080 16497 3108
rect 16264 3068 16270 3080
rect 16485 3077 16497 3080
rect 16531 3077 16543 3111
rect 16485 3071 16543 3077
rect 17954 3068 17960 3120
rect 18012 3108 18018 3120
rect 18509 3111 18567 3117
rect 18509 3108 18521 3111
rect 18012 3080 18521 3108
rect 18012 3068 18018 3080
rect 18509 3077 18521 3080
rect 18555 3077 18567 3111
rect 22833 3111 22891 3117
rect 22833 3108 22845 3111
rect 18509 3071 18567 3077
rect 19352 3080 22845 3108
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3040 9183 3043
rect 9171 3012 9812 3040
rect 9171 3009 9183 3012
rect 9125 3003 9183 3009
rect 9214 2972 9220 2984
rect 7975 2944 8800 2972
rect 9175 2944 9220 2972
rect 7975 2941 7987 2944
rect 7929 2935 7987 2941
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 9784 2981 9812 3012
rect 9769 2975 9827 2981
rect 9769 2941 9781 2975
rect 9815 2972 9827 2975
rect 10244 2972 10272 3068
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13814 3040 13820 3052
rect 13219 3012 13820 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 15194 3040 15200 3052
rect 15155 3012 15200 3040
rect 15194 3000 15200 3012
rect 15252 3000 15258 3052
rect 16758 3000 16764 3052
rect 16816 3040 16822 3052
rect 17773 3043 17831 3049
rect 17773 3040 17785 3043
rect 16816 3012 17785 3040
rect 16816 3000 16822 3012
rect 17773 3009 17785 3012
rect 17819 3040 17831 3043
rect 18414 3040 18420 3052
rect 17819 3012 18420 3040
rect 17819 3009 17831 3012
rect 17773 3003 17831 3009
rect 18414 3000 18420 3012
rect 18472 3000 18478 3052
rect 19352 3049 19380 3080
rect 22833 3077 22845 3080
rect 22879 3077 22891 3111
rect 23474 3108 23480 3120
rect 23435 3080 23480 3108
rect 22833 3071 22891 3077
rect 23474 3068 23480 3080
rect 23532 3068 23538 3120
rect 29472 3080 30328 3108
rect 19337 3043 19395 3049
rect 19337 3009 19349 3043
rect 19383 3009 19395 3043
rect 19337 3003 19395 3009
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 20533 3043 20591 3049
rect 20533 3040 20545 3043
rect 19484 3012 20545 3040
rect 19484 3000 19490 3012
rect 20533 3009 20545 3012
rect 20579 3009 20591 3043
rect 20533 3003 20591 3009
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3040 20867 3043
rect 21818 3040 21824 3052
rect 20855 3012 21824 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 22094 3000 22100 3052
rect 22152 3040 22158 3052
rect 22373 3043 22431 3049
rect 22373 3040 22385 3043
rect 22152 3012 22385 3040
rect 22152 3000 22158 3012
rect 22373 3009 22385 3012
rect 22419 3009 22431 3043
rect 23492 3040 23520 3068
rect 29472 3052 29500 3080
rect 22373 3003 22431 3009
rect 22664 3012 23520 3040
rect 23661 3043 23719 3049
rect 11422 2981 11428 2984
rect 9815 2944 10272 2972
rect 11400 2975 11428 2981
rect 9815 2941 9827 2944
rect 9769 2935 9827 2941
rect 11400 2941 11412 2975
rect 11480 2972 11486 2984
rect 13300 2975 13358 2981
rect 13300 2972 13312 2975
rect 11480 2944 12296 2972
rect 11400 2935 11428 2941
rect 11422 2932 11428 2935
rect 11480 2932 11486 2944
rect 12268 2916 12296 2944
rect 12360 2944 13312 2972
rect 8386 2904 8392 2916
rect 4396 2876 7420 2904
rect 7668 2876 8392 2904
rect 4396 2864 4402 2876
rect 4246 2836 4252 2848
rect 4207 2808 4252 2836
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 7098 2836 7104 2848
rect 7059 2808 7104 2836
rect 7098 2796 7104 2808
rect 7156 2796 7162 2848
rect 7392 2836 7420 2876
rect 8386 2864 8392 2876
rect 8444 2864 8450 2916
rect 12250 2904 12256 2916
rect 9140 2876 12112 2904
rect 12211 2876 12256 2904
rect 9140 2836 9168 2876
rect 9306 2836 9312 2848
rect 7392 2808 9168 2836
rect 9267 2808 9312 2836
rect 9306 2796 9312 2808
rect 9364 2796 9370 2848
rect 11885 2839 11943 2845
rect 11885 2805 11897 2839
rect 11931 2836 11943 2839
rect 11974 2836 11980 2848
rect 11931 2808 11980 2836
rect 11931 2805 11943 2808
rect 11885 2799 11943 2805
rect 11974 2796 11980 2808
rect 12032 2796 12038 2848
rect 12084 2836 12112 2876
rect 12250 2864 12256 2876
rect 12308 2864 12314 2916
rect 12360 2836 12388 2944
rect 13300 2941 13312 2944
rect 13346 2972 13358 2975
rect 14093 2975 14151 2981
rect 14093 2972 14105 2975
rect 13346 2944 14105 2972
rect 13346 2941 13358 2944
rect 13300 2935 13358 2941
rect 14093 2941 14105 2944
rect 14139 2941 14151 2975
rect 14093 2935 14151 2941
rect 14737 2975 14795 2981
rect 14737 2941 14749 2975
rect 14783 2972 14795 2975
rect 14918 2972 14924 2984
rect 14783 2944 14924 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 13817 2907 13875 2913
rect 13817 2873 13829 2907
rect 13863 2904 13875 2907
rect 13906 2904 13912 2916
rect 13863 2876 13912 2904
rect 13863 2873 13875 2876
rect 13817 2867 13875 2873
rect 13906 2864 13912 2876
rect 13964 2864 13970 2916
rect 12084 2808 12388 2836
rect 14108 2836 14136 2935
rect 14918 2932 14924 2944
rect 14976 2981 14982 2984
rect 14976 2975 15034 2981
rect 14976 2941 14988 2975
rect 15022 2972 15034 2975
rect 16025 2975 16083 2981
rect 16025 2972 16037 2975
rect 15022 2944 16037 2972
rect 15022 2941 15034 2944
rect 14976 2935 15034 2941
rect 16025 2941 16037 2944
rect 16071 2972 16083 2975
rect 16390 2972 16396 2984
rect 16071 2944 16396 2972
rect 16071 2941 16083 2944
rect 16025 2935 16083 2941
rect 14976 2932 14982 2935
rect 16390 2932 16396 2944
rect 16448 2932 16454 2984
rect 16666 2972 16672 2984
rect 16627 2944 16672 2972
rect 16666 2932 16672 2944
rect 16724 2932 16730 2984
rect 17129 2975 17187 2981
rect 17129 2941 17141 2975
rect 17175 2972 17187 2975
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 17175 2944 18061 2972
rect 17175 2941 17187 2944
rect 17129 2935 17187 2941
rect 18049 2941 18061 2944
rect 18095 2972 18107 2975
rect 18322 2972 18328 2984
rect 18095 2944 18328 2972
rect 18095 2941 18107 2944
rect 18049 2935 18107 2941
rect 18322 2932 18328 2944
rect 18380 2932 18386 2984
rect 22664 2981 22692 3012
rect 23661 3009 23673 3043
rect 23707 3040 23719 3043
rect 24578 3040 24584 3052
rect 23707 3012 24584 3040
rect 23707 3009 23719 3012
rect 23661 3003 23719 3009
rect 22624 2975 22692 2981
rect 22624 2972 22636 2975
rect 20088 2944 22636 2972
rect 14826 2904 14832 2916
rect 14787 2876 14832 2904
rect 14826 2864 14832 2876
rect 14884 2864 14890 2916
rect 17328 2876 19380 2904
rect 17328 2836 17356 2876
rect 14108 2808 17356 2836
rect 19153 2839 19211 2845
rect 19153 2805 19165 2839
rect 19199 2836 19211 2839
rect 19242 2836 19248 2848
rect 19199 2808 19248 2836
rect 19199 2805 19211 2808
rect 19153 2799 19211 2805
rect 19242 2796 19248 2808
rect 19300 2796 19306 2848
rect 19352 2836 19380 2876
rect 19426 2864 19432 2916
rect 19484 2904 19490 2916
rect 19978 2904 19984 2916
rect 19484 2876 19529 2904
rect 19939 2876 19984 2904
rect 19484 2864 19490 2876
rect 19978 2864 19984 2876
rect 20036 2864 20042 2916
rect 20088 2836 20116 2944
rect 22624 2941 22636 2944
rect 22670 2944 22692 2975
rect 22670 2941 22682 2944
rect 22624 2935 22682 2941
rect 22738 2932 22744 2984
rect 22796 2972 22802 2984
rect 23676 2972 23704 3003
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 26326 3040 26332 3052
rect 26287 3012 26332 3040
rect 26326 3000 26332 3012
rect 26384 3000 26390 3052
rect 27706 3000 27712 3052
rect 27764 3040 27770 3052
rect 28629 3043 28687 3049
rect 28629 3040 28641 3043
rect 27764 3012 28641 3040
rect 27764 3000 27770 3012
rect 27816 2981 27844 3012
rect 28629 3009 28641 3012
rect 28675 3009 28687 3043
rect 29454 3040 29460 3052
rect 29367 3012 29460 3040
rect 28629 3003 28687 3009
rect 29454 3000 29460 3012
rect 29512 3000 29518 3052
rect 30098 3040 30104 3052
rect 30059 3012 30104 3040
rect 30098 3000 30104 3012
rect 30156 3000 30162 3052
rect 30300 3040 30328 3080
rect 30929 3043 30987 3049
rect 30929 3040 30941 3043
rect 30300 3012 30941 3040
rect 30929 3009 30941 3012
rect 30975 3009 30987 3043
rect 30929 3003 30987 3009
rect 25593 2975 25651 2981
rect 25593 2972 25605 2975
rect 22796 2944 23704 2972
rect 23860 2944 25605 2972
rect 22796 2932 22802 2944
rect 20254 2904 20260 2916
rect 20215 2876 20260 2904
rect 20254 2864 20260 2876
rect 20312 2864 20318 2916
rect 20533 2907 20591 2913
rect 20533 2873 20545 2907
rect 20579 2904 20591 2907
rect 20579 2876 20852 2904
rect 20579 2873 20591 2876
rect 20533 2867 20591 2873
rect 20622 2836 20628 2848
rect 19352 2808 20116 2836
rect 20583 2808 20628 2836
rect 20622 2796 20628 2808
rect 20680 2796 20686 2848
rect 20824 2836 20852 2876
rect 20898 2864 20904 2916
rect 20956 2904 20962 2916
rect 21130 2907 21188 2913
rect 21130 2904 21142 2907
rect 20956 2876 21142 2904
rect 20956 2864 20962 2876
rect 21130 2873 21142 2876
rect 21176 2873 21188 2907
rect 21130 2867 21188 2873
rect 22833 2907 22891 2913
rect 22833 2873 22845 2907
rect 22879 2904 22891 2907
rect 23860 2904 23888 2944
rect 25593 2941 25605 2944
rect 25639 2941 25651 2975
rect 25593 2935 25651 2941
rect 27801 2975 27859 2981
rect 27801 2941 27813 2975
rect 27847 2941 27859 2975
rect 27801 2935 27859 2941
rect 23979 2904 23985 2916
rect 22879 2876 23888 2904
rect 23940 2876 23985 2904
rect 22879 2873 22891 2876
rect 22833 2867 22891 2873
rect 23979 2864 23985 2876
rect 24037 2864 24043 2916
rect 26145 2907 26203 2913
rect 26145 2873 26157 2907
rect 26191 2904 26203 2907
rect 26421 2907 26479 2913
rect 26421 2904 26433 2907
rect 26191 2876 26433 2904
rect 26191 2873 26203 2876
rect 26145 2867 26203 2873
rect 26421 2873 26433 2876
rect 26467 2904 26479 2907
rect 26510 2904 26516 2916
rect 26467 2876 26516 2904
rect 26467 2873 26479 2876
rect 26421 2867 26479 2873
rect 26510 2864 26516 2876
rect 26568 2864 26574 2916
rect 26970 2904 26976 2916
rect 26931 2876 26976 2904
rect 26970 2864 26976 2876
rect 27028 2864 27034 2916
rect 29546 2864 29552 2916
rect 29604 2904 29610 2916
rect 29604 2876 29649 2904
rect 29604 2864 29610 2876
rect 21450 2836 21456 2848
rect 20824 2808 21456 2836
rect 21450 2796 21456 2808
rect 21508 2836 21514 2848
rect 21729 2839 21787 2845
rect 21729 2836 21741 2839
rect 21508 2808 21741 2836
rect 21508 2796 21514 2808
rect 21729 2805 21741 2808
rect 21775 2836 21787 2839
rect 21910 2836 21916 2848
rect 21775 2808 21916 2836
rect 21775 2805 21787 2808
rect 21729 2799 21787 2805
rect 21910 2796 21916 2808
rect 21968 2796 21974 2848
rect 22094 2836 22100 2848
rect 22055 2808 22100 2836
rect 22094 2796 22100 2808
rect 22152 2796 22158 2848
rect 22554 2796 22560 2848
rect 22612 2836 22618 2848
rect 22925 2839 22983 2845
rect 22925 2836 22937 2839
rect 22612 2808 22937 2836
rect 22612 2796 22618 2808
rect 22925 2805 22937 2808
rect 22971 2836 22983 2839
rect 23017 2839 23075 2845
rect 23017 2836 23029 2839
rect 22971 2808 23029 2836
rect 22971 2805 22983 2808
rect 22925 2799 22983 2805
rect 23017 2805 23029 2808
rect 23063 2805 23075 2839
rect 23017 2799 23075 2805
rect 23566 2796 23572 2848
rect 23624 2836 23630 2848
rect 24581 2839 24639 2845
rect 24581 2836 24593 2839
rect 23624 2808 24593 2836
rect 23624 2796 23630 2808
rect 24581 2805 24593 2808
rect 24627 2836 24639 2839
rect 24854 2836 24860 2848
rect 24627 2808 24860 2836
rect 24627 2805 24639 2808
rect 24581 2799 24639 2805
rect 24854 2796 24860 2808
rect 24912 2836 24918 2848
rect 25225 2839 25283 2845
rect 25225 2836 25237 2839
rect 24912 2808 25237 2836
rect 24912 2796 24918 2808
rect 25225 2805 25237 2808
rect 25271 2805 25283 2839
rect 25225 2799 25283 2805
rect 28353 2839 28411 2845
rect 28353 2805 28365 2839
rect 28399 2836 28411 2839
rect 28442 2836 28448 2848
rect 28399 2808 28448 2836
rect 28399 2805 28411 2808
rect 28353 2799 28411 2805
rect 28442 2796 28448 2808
rect 28500 2796 28506 2848
rect 29089 2839 29147 2845
rect 29089 2805 29101 2839
rect 29135 2836 29147 2839
rect 29564 2836 29592 2864
rect 29135 2808 29592 2836
rect 29135 2805 29147 2808
rect 29089 2799 29147 2805
rect 29822 2796 29828 2848
rect 29880 2836 29886 2848
rect 30377 2839 30435 2845
rect 30377 2836 30389 2839
rect 29880 2808 30389 2836
rect 29880 2796 29886 2808
rect 30377 2805 30389 2808
rect 30423 2805 30435 2839
rect 30377 2799 30435 2805
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 2041 2635 2099 2641
rect 2041 2601 2053 2635
rect 2087 2632 2099 2635
rect 2130 2632 2136 2644
rect 2087 2604 2136 2632
rect 2087 2601 2099 2604
rect 2041 2595 2099 2601
rect 2130 2592 2136 2604
rect 2188 2592 2194 2644
rect 2363 2635 2421 2641
rect 2363 2601 2375 2635
rect 2409 2632 2421 2635
rect 2958 2632 2964 2644
rect 2409 2604 2964 2632
rect 2409 2601 2421 2604
rect 2363 2595 2421 2601
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 7466 2592 7472 2644
rect 7524 2632 7530 2644
rect 8113 2635 8171 2641
rect 8113 2632 8125 2635
rect 7524 2604 8125 2632
rect 7524 2592 7530 2604
rect 8113 2601 8125 2604
rect 8159 2601 8171 2635
rect 10042 2632 10048 2644
rect 10003 2604 10048 2632
rect 8113 2595 8171 2601
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 11655 2635 11713 2641
rect 11655 2601 11667 2635
rect 11701 2632 11713 2635
rect 11882 2632 11888 2644
rect 11701 2604 11888 2632
rect 11701 2601 11713 2604
rect 11655 2595 11713 2601
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12943 2635 13001 2641
rect 12943 2601 12955 2635
rect 12989 2632 13001 2635
rect 14734 2632 14740 2644
rect 12989 2604 14740 2632
rect 12989 2601 13001 2604
rect 12943 2595 13001 2601
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 14921 2635 14979 2641
rect 14921 2601 14933 2635
rect 14967 2632 14979 2635
rect 15102 2632 15108 2644
rect 14967 2604 15108 2632
rect 14967 2601 14979 2604
rect 14921 2595 14979 2601
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 16390 2592 16396 2644
rect 16448 2632 16454 2644
rect 16577 2635 16635 2641
rect 16577 2632 16589 2635
rect 16448 2604 16589 2632
rect 16448 2592 16454 2604
rect 16577 2601 16589 2604
rect 16623 2601 16635 2635
rect 16577 2595 16635 2601
rect 16758 2592 16764 2644
rect 16816 2632 16822 2644
rect 17313 2635 17371 2641
rect 17313 2632 17325 2635
rect 16816 2604 17325 2632
rect 16816 2592 16822 2604
rect 17313 2601 17325 2604
rect 17359 2601 17371 2635
rect 18046 2632 18052 2644
rect 18007 2604 18052 2632
rect 17313 2595 17371 2601
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 18598 2592 18604 2644
rect 18656 2632 18662 2644
rect 18693 2635 18751 2641
rect 18693 2632 18705 2635
rect 18656 2604 18705 2632
rect 18656 2592 18662 2604
rect 18693 2601 18705 2604
rect 18739 2601 18751 2635
rect 18693 2595 18751 2601
rect 19061 2635 19119 2641
rect 19061 2601 19073 2635
rect 19107 2632 19119 2635
rect 19150 2632 19156 2644
rect 19107 2604 19156 2632
rect 19107 2601 19119 2604
rect 19061 2595 19119 2601
rect 7834 2564 7840 2576
rect 7795 2536 7840 2564
rect 7834 2524 7840 2536
rect 7892 2524 7898 2576
rect 9585 2567 9643 2573
rect 9585 2533 9597 2567
rect 9631 2564 9643 2567
rect 9631 2536 10272 2564
rect 9631 2533 9643 2536
rect 9585 2527 9643 2533
rect 10244 2508 10272 2536
rect 13814 2524 13820 2576
rect 13872 2564 13878 2576
rect 14553 2567 14611 2573
rect 14553 2564 14565 2567
rect 13872 2536 14565 2564
rect 13872 2524 13878 2536
rect 14553 2533 14565 2536
rect 14599 2564 14611 2567
rect 18874 2564 18880 2576
rect 14599 2536 18880 2564
rect 14599 2533 14611 2536
rect 14553 2527 14611 2533
rect 18874 2524 18880 2536
rect 18932 2524 18938 2576
rect 106 2456 112 2508
rect 164 2496 170 2508
rect 2260 2499 2318 2505
rect 2260 2496 2272 2499
rect 164 2468 2272 2496
rect 164 2456 170 2468
rect 2260 2465 2272 2468
rect 2306 2496 2318 2499
rect 2685 2499 2743 2505
rect 2685 2496 2697 2499
rect 2306 2468 2697 2496
rect 2306 2465 2318 2468
rect 2260 2459 2318 2465
rect 2685 2465 2697 2468
rect 2731 2496 2743 2499
rect 5534 2496 5540 2508
rect 2731 2468 5540 2496
rect 2731 2465 2743 2468
rect 2685 2459 2743 2465
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7098 2496 7104 2508
rect 6779 2468 7104 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 7098 2456 7104 2468
rect 7156 2496 7162 2508
rect 7745 2499 7803 2505
rect 7745 2496 7757 2499
rect 7156 2468 7757 2496
rect 7156 2456 7162 2468
rect 7745 2465 7757 2468
rect 7791 2496 7803 2499
rect 8018 2496 8024 2508
rect 7791 2468 8024 2496
rect 7791 2465 7803 2468
rect 7745 2459 7803 2465
rect 8018 2456 8024 2468
rect 8076 2456 8082 2508
rect 8110 2456 8116 2508
rect 8168 2496 8174 2508
rect 8665 2499 8723 2505
rect 8665 2496 8677 2499
rect 8168 2468 8677 2496
rect 8168 2456 8174 2468
rect 8665 2465 8677 2468
rect 8711 2496 8723 2499
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8711 2468 9137 2496
rect 8711 2465 8723 2468
rect 8665 2459 8723 2465
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 10042 2496 10048 2508
rect 10003 2468 10048 2496
rect 9125 2459 9183 2465
rect 10042 2456 10048 2468
rect 10100 2456 10106 2508
rect 10226 2496 10232 2508
rect 10187 2468 10232 2496
rect 10226 2456 10232 2468
rect 10284 2456 10290 2508
rect 11584 2499 11642 2505
rect 11584 2465 11596 2499
rect 11630 2496 11642 2499
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11630 2468 11989 2496
rect 11630 2465 11642 2468
rect 11584 2459 11642 2465
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 12872 2499 12930 2505
rect 12872 2465 12884 2499
rect 12918 2496 12930 2499
rect 13354 2496 13360 2508
rect 12918 2468 13360 2496
rect 12918 2465 12930 2468
rect 12872 2459 12930 2465
rect 8294 2388 8300 2440
rect 8352 2428 8358 2440
rect 11599 2428 11627 2459
rect 8352 2400 11627 2428
rect 11992 2428 12020 2459
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 13725 2499 13783 2505
rect 13725 2465 13737 2499
rect 13771 2496 13783 2499
rect 14461 2499 14519 2505
rect 14461 2496 14473 2499
rect 13771 2468 14473 2496
rect 13771 2465 13783 2468
rect 13725 2459 13783 2465
rect 14461 2465 14473 2468
rect 14507 2496 14519 2499
rect 14826 2496 14832 2508
rect 14507 2468 14832 2496
rect 14507 2465 14519 2468
rect 14461 2459 14519 2465
rect 14826 2456 14832 2468
rect 14884 2456 14890 2508
rect 15194 2456 15200 2508
rect 15252 2496 15258 2508
rect 15657 2499 15715 2505
rect 15657 2496 15669 2499
rect 15252 2468 15669 2496
rect 15252 2456 15258 2468
rect 15657 2465 15669 2468
rect 15703 2465 15715 2499
rect 15657 2459 15715 2465
rect 16301 2499 16359 2505
rect 16301 2465 16313 2499
rect 16347 2496 16359 2499
rect 16666 2496 16672 2508
rect 16347 2468 16672 2496
rect 16347 2465 16359 2468
rect 16301 2459 16359 2465
rect 16666 2456 16672 2468
rect 16724 2496 16730 2508
rect 16945 2499 17003 2505
rect 16945 2496 16957 2499
rect 16724 2468 16957 2496
rect 16724 2456 16730 2468
rect 16945 2465 16957 2468
rect 16991 2496 17003 2499
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 16991 2468 17141 2496
rect 16991 2465 17003 2468
rect 16945 2459 17003 2465
rect 17129 2465 17141 2468
rect 17175 2496 17187 2499
rect 17589 2499 17647 2505
rect 17589 2496 17601 2499
rect 17175 2468 17601 2496
rect 17175 2465 17187 2468
rect 17129 2459 17187 2465
rect 17589 2465 17601 2468
rect 17635 2465 17647 2499
rect 17589 2459 17647 2465
rect 18509 2499 18567 2505
rect 18509 2465 18521 2499
rect 18555 2496 18567 2499
rect 19076 2496 19104 2595
rect 19150 2592 19156 2604
rect 19208 2592 19214 2644
rect 20898 2632 20904 2644
rect 20859 2604 20904 2632
rect 20898 2592 20904 2604
rect 20956 2592 20962 2644
rect 21634 2632 21640 2644
rect 21595 2604 21640 2632
rect 21634 2592 21640 2604
rect 21692 2592 21698 2644
rect 21910 2592 21916 2644
rect 21968 2632 21974 2644
rect 22005 2635 22063 2641
rect 22005 2632 22017 2635
rect 21968 2604 22017 2632
rect 21968 2592 21974 2604
rect 22005 2601 22017 2604
rect 22051 2601 22063 2635
rect 23750 2632 23756 2644
rect 23711 2604 23756 2632
rect 22005 2595 22063 2601
rect 23750 2592 23756 2604
rect 23808 2592 23814 2644
rect 25222 2632 25228 2644
rect 24412 2604 25228 2632
rect 19429 2567 19487 2573
rect 19429 2533 19441 2567
rect 19475 2564 19487 2567
rect 19702 2564 19708 2576
rect 19475 2536 19708 2564
rect 19475 2533 19487 2536
rect 19429 2527 19487 2533
rect 19702 2524 19708 2536
rect 19760 2524 19766 2576
rect 19978 2524 19984 2576
rect 20036 2564 20042 2576
rect 20257 2567 20315 2573
rect 20257 2564 20269 2567
rect 20036 2536 20269 2564
rect 20036 2524 20042 2536
rect 20257 2533 20269 2536
rect 20303 2564 20315 2567
rect 21453 2567 21511 2573
rect 21453 2564 21465 2567
rect 20303 2536 21465 2564
rect 20303 2533 20315 2536
rect 20257 2527 20315 2533
rect 21453 2533 21465 2536
rect 21499 2533 21511 2567
rect 21453 2527 21511 2533
rect 18555 2468 19104 2496
rect 21244 2499 21302 2505
rect 18555 2465 18567 2468
rect 18509 2459 18567 2465
rect 21244 2465 21256 2499
rect 21290 2496 21302 2499
rect 21652 2496 21680 2592
rect 22557 2567 22615 2573
rect 22557 2533 22569 2567
rect 22603 2564 22615 2567
rect 23566 2564 23572 2576
rect 22603 2536 23572 2564
rect 22603 2533 22615 2536
rect 22557 2527 22615 2533
rect 23566 2524 23572 2536
rect 23624 2524 23630 2576
rect 24314 2567 24372 2573
rect 24314 2533 24326 2567
rect 24360 2564 24372 2567
rect 24412 2564 24440 2604
rect 25222 2592 25228 2604
rect 25280 2592 25286 2644
rect 26234 2592 26240 2644
rect 26292 2632 26298 2644
rect 27019 2635 27077 2641
rect 27019 2632 27031 2635
rect 26292 2604 27031 2632
rect 26292 2592 26298 2604
rect 27019 2601 27031 2604
rect 27065 2601 27077 2635
rect 29086 2632 29092 2644
rect 29047 2604 29092 2632
rect 27019 2595 27077 2601
rect 29086 2592 29092 2604
rect 29144 2592 29150 2644
rect 29454 2632 29460 2644
rect 29415 2604 29460 2632
rect 29454 2592 29460 2604
rect 29512 2592 29518 2644
rect 24360 2536 24440 2564
rect 24360 2533 24372 2536
rect 24314 2527 24372 2533
rect 24486 2524 24492 2576
rect 24544 2564 24550 2576
rect 26513 2567 26571 2573
rect 26513 2564 26525 2567
rect 24544 2536 26525 2564
rect 24544 2524 24550 2536
rect 26513 2533 26525 2536
rect 26559 2533 26571 2567
rect 26513 2527 26571 2533
rect 26620 2536 27971 2564
rect 21290 2468 21680 2496
rect 23109 2499 23167 2505
rect 21290 2465 21302 2468
rect 21244 2459 21302 2465
rect 23109 2465 23121 2499
rect 23155 2496 23167 2499
rect 24026 2496 24032 2508
rect 23155 2468 24032 2496
rect 23155 2465 23167 2468
rect 23109 2459 23167 2465
rect 24026 2456 24032 2468
rect 24084 2456 24090 2508
rect 24854 2456 24860 2508
rect 24912 2496 24918 2508
rect 26620 2496 26648 2536
rect 24912 2468 26648 2496
rect 26948 2499 27006 2505
rect 24912 2456 24918 2468
rect 26948 2465 26960 2499
rect 26994 2496 27006 2499
rect 27430 2496 27436 2508
rect 26994 2468 27436 2496
rect 26994 2465 27006 2468
rect 26948 2459 27006 2465
rect 27430 2456 27436 2468
rect 27488 2456 27494 2508
rect 27943 2505 27971 2536
rect 27928 2499 27986 2505
rect 27928 2465 27940 2499
rect 27974 2496 27986 2499
rect 28353 2499 28411 2505
rect 28353 2496 28365 2499
rect 27974 2468 28365 2496
rect 27974 2465 27986 2468
rect 27928 2459 27986 2465
rect 28353 2465 28365 2468
rect 28399 2465 28411 2499
rect 29104 2496 29132 2592
rect 29546 2524 29552 2576
rect 29604 2564 29610 2576
rect 29733 2567 29791 2573
rect 29733 2564 29745 2567
rect 29604 2536 29745 2564
rect 29604 2524 29610 2536
rect 29733 2533 29745 2536
rect 29779 2533 29791 2567
rect 29733 2527 29791 2533
rect 29822 2496 29828 2508
rect 29104 2468 29828 2496
rect 28353 2459 28411 2465
rect 29822 2456 29828 2468
rect 29880 2456 29886 2508
rect 30098 2456 30104 2508
rect 30156 2496 30162 2508
rect 31332 2499 31390 2505
rect 31332 2496 31344 2499
rect 30156 2468 31344 2496
rect 30156 2456 30162 2468
rect 31332 2465 31344 2468
rect 31378 2496 31390 2499
rect 31757 2499 31815 2505
rect 31757 2496 31769 2499
rect 31378 2468 31769 2496
rect 31378 2465 31390 2468
rect 31332 2459 31390 2465
rect 31757 2465 31769 2468
rect 31803 2465 31815 2499
rect 31757 2459 31815 2465
rect 18966 2428 18972 2440
rect 11992 2400 18972 2428
rect 8352 2388 8358 2400
rect 18966 2388 18972 2400
rect 19024 2388 19030 2440
rect 19613 2431 19671 2437
rect 19613 2397 19625 2431
rect 19659 2428 19671 2431
rect 21453 2431 21511 2437
rect 19659 2400 21358 2428
rect 19659 2397 19671 2400
rect 19613 2391 19671 2397
rect 7282 2320 7288 2372
rect 7340 2360 7346 2372
rect 8849 2363 8907 2369
rect 8849 2360 8861 2363
rect 7340 2332 8861 2360
rect 7340 2320 7346 2332
rect 8849 2329 8861 2332
rect 8895 2360 8907 2363
rect 10042 2360 10048 2372
rect 8895 2332 10048 2360
rect 8895 2329 8907 2332
rect 8849 2323 8907 2329
rect 10042 2320 10048 2332
rect 10100 2360 10106 2372
rect 21330 2369 21358 2400
rect 21453 2397 21465 2431
rect 21499 2428 21511 2431
rect 22465 2431 22523 2437
rect 22465 2428 22477 2431
rect 21499 2400 22477 2428
rect 21499 2397 21511 2400
rect 21453 2391 21511 2397
rect 22465 2397 22477 2400
rect 22511 2428 22523 2431
rect 23845 2431 23903 2437
rect 23845 2428 23857 2431
rect 22511 2400 23857 2428
rect 22511 2397 22523 2400
rect 22465 2391 22523 2397
rect 23845 2397 23857 2400
rect 23891 2397 23903 2431
rect 23845 2391 23903 2397
rect 24213 2431 24271 2437
rect 24213 2397 24225 2431
rect 24259 2428 24271 2431
rect 25501 2431 25559 2437
rect 25501 2428 25513 2431
rect 24259 2400 25513 2428
rect 24259 2397 24271 2400
rect 24213 2391 24271 2397
rect 25501 2397 25513 2400
rect 25547 2428 25559 2431
rect 25685 2431 25743 2437
rect 25685 2428 25697 2431
rect 25547 2400 25697 2428
rect 25547 2397 25559 2400
rect 25501 2391 25559 2397
rect 25685 2397 25697 2400
rect 25731 2397 25743 2431
rect 25685 2391 25743 2397
rect 10781 2363 10839 2369
rect 10781 2360 10793 2363
rect 10100 2332 10793 2360
rect 10100 2320 10106 2332
rect 10781 2329 10793 2332
rect 10827 2329 10839 2363
rect 10781 2323 10839 2329
rect 21315 2363 21373 2369
rect 21315 2329 21327 2363
rect 21361 2360 21373 2363
rect 26145 2363 26203 2369
rect 26145 2360 26157 2363
rect 21361 2332 24716 2360
rect 21361 2329 21373 2332
rect 21315 2323 21373 2329
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8573 2295 8631 2301
rect 8573 2292 8585 2295
rect 8444 2264 8585 2292
rect 8444 2252 8450 2264
rect 8573 2261 8585 2264
rect 8619 2292 8631 2295
rect 12342 2292 12348 2304
rect 8619 2264 12348 2292
rect 8619 2261 8631 2264
rect 8573 2255 8631 2261
rect 12342 2252 12348 2264
rect 12400 2252 12406 2304
rect 13354 2292 13360 2304
rect 13315 2264 13360 2292
rect 13354 2252 13360 2264
rect 13412 2252 13418 2304
rect 15194 2292 15200 2304
rect 15155 2264 15200 2292
rect 15194 2252 15200 2264
rect 15252 2252 15258 2304
rect 19242 2252 19248 2304
rect 19300 2292 19306 2304
rect 21450 2292 21456 2304
rect 19300 2264 21456 2292
rect 19300 2252 19306 2264
rect 21450 2252 21456 2264
rect 21508 2252 21514 2304
rect 23845 2295 23903 2301
rect 23845 2261 23857 2295
rect 23891 2292 23903 2295
rect 24486 2292 24492 2304
rect 23891 2264 24492 2292
rect 23891 2261 23903 2264
rect 23845 2255 23903 2261
rect 24486 2252 24492 2264
rect 24544 2252 24550 2304
rect 24688 2292 24716 2332
rect 24872 2332 26157 2360
rect 24872 2292 24900 2332
rect 26145 2329 26157 2332
rect 26191 2329 26203 2363
rect 26145 2323 26203 2329
rect 31435 2363 31493 2369
rect 31435 2329 31447 2363
rect 31481 2360 31493 2363
rect 38378 2360 38384 2372
rect 31481 2332 38384 2360
rect 31481 2329 31493 2332
rect 31435 2323 31493 2329
rect 38378 2320 38384 2332
rect 38436 2320 38442 2372
rect 27430 2292 27436 2304
rect 24688 2264 24900 2292
rect 27391 2264 27436 2292
rect 27430 2252 27436 2264
rect 27488 2252 27494 2304
rect 28031 2295 28089 2301
rect 28031 2261 28043 2295
rect 28077 2292 28089 2295
rect 28258 2292 28264 2304
rect 28077 2264 28264 2292
rect 28077 2261 28089 2264
rect 28031 2255 28089 2261
rect 28258 2252 28264 2264
rect 28316 2252 28322 2304
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
rect 25406 76 25412 128
rect 25464 116 25470 128
rect 31662 116 31668 128
rect 25464 88 31668 116
rect 25464 76 25470 88
rect 31662 76 31668 88
rect 31720 76 31726 128
<< via1 >>
rect 5908 15512 5960 15564
rect 7472 15512 7524 15564
rect 31208 15512 31260 15564
rect 32496 15512 32548 15564
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 2412 13336 2464 13388
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 112 12928 164 12980
rect 24124 12656 24176 12708
rect 2136 12588 2188 12640
rect 2412 12631 2464 12640
rect 2412 12597 2421 12631
rect 2421 12597 2455 12631
rect 2455 12597 2464 12631
rect 2412 12588 2464 12597
rect 24584 12588 24636 12640
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 39580 12384 39632 12436
rect 1400 12248 1452 12300
rect 3056 12248 3108 12300
rect 11152 12248 11204 12300
rect 19156 12291 19208 12300
rect 19156 12257 19165 12291
rect 19165 12257 19199 12291
rect 19199 12257 19208 12291
rect 19156 12248 19208 12257
rect 24216 12248 24268 12300
rect 25320 12248 25372 12300
rect 34612 12248 34664 12300
rect 35440 12291 35492 12300
rect 35440 12257 35449 12291
rect 35449 12257 35483 12291
rect 35483 12257 35492 12291
rect 35440 12248 35492 12257
rect 29552 12223 29604 12232
rect 29552 12189 29561 12223
rect 29561 12189 29595 12223
rect 29595 12189 29604 12223
rect 29552 12180 29604 12189
rect 2320 12044 2372 12096
rect 2504 12044 2556 12096
rect 10140 12087 10192 12096
rect 10140 12053 10149 12087
rect 10149 12053 10183 12087
rect 10183 12053 10192 12087
rect 10140 12044 10192 12053
rect 11428 12044 11480 12096
rect 18144 12044 18196 12096
rect 24400 12044 24452 12096
rect 24768 12044 24820 12096
rect 34796 12044 34848 12096
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 112 11840 164 11892
rect 22100 11840 22152 11892
rect 19616 11772 19668 11824
rect 29828 11772 29880 11824
rect 8300 11704 8352 11756
rect 10140 11704 10192 11756
rect 2872 11568 2924 11620
rect 1400 11500 1452 11552
rect 3056 11543 3108 11552
rect 3056 11509 3065 11543
rect 3065 11509 3099 11543
rect 3099 11509 3108 11543
rect 3056 11500 3108 11509
rect 4712 11636 4764 11688
rect 6644 11636 6696 11688
rect 11980 11704 12032 11756
rect 24216 11704 24268 11756
rect 28448 11704 28500 11756
rect 15660 11636 15712 11688
rect 10784 11611 10836 11620
rect 10784 11577 10793 11611
rect 10793 11577 10827 11611
rect 10827 11577 10836 11611
rect 10784 11568 10836 11577
rect 3608 11500 3660 11552
rect 10416 11500 10468 11552
rect 11152 11543 11204 11552
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 11152 11500 11204 11509
rect 15936 11500 15988 11552
rect 16580 11500 16632 11552
rect 19156 11500 19208 11552
rect 19708 11543 19760 11552
rect 19708 11509 19717 11543
rect 19717 11509 19751 11543
rect 19751 11509 19760 11543
rect 19708 11500 19760 11509
rect 21364 11636 21416 11688
rect 25320 11679 25372 11688
rect 25320 11645 25329 11679
rect 25329 11645 25363 11679
rect 25363 11645 25372 11679
rect 25320 11636 25372 11645
rect 22008 11568 22060 11620
rect 33600 11840 33652 11892
rect 35440 11840 35492 11892
rect 35624 11883 35676 11892
rect 35624 11849 35633 11883
rect 35633 11849 35667 11883
rect 35667 11849 35676 11883
rect 35624 11840 35676 11849
rect 37188 11840 37240 11892
rect 34428 11704 34480 11756
rect 32588 11636 32640 11688
rect 35164 11636 35216 11688
rect 33416 11568 33468 11620
rect 34612 11611 34664 11620
rect 21640 11500 21692 11552
rect 24676 11500 24728 11552
rect 25412 11543 25464 11552
rect 25412 11509 25421 11543
rect 25421 11509 25455 11543
rect 25455 11509 25464 11543
rect 25412 11500 25464 11509
rect 30288 11500 30340 11552
rect 31484 11500 31536 11552
rect 31852 11500 31904 11552
rect 34612 11577 34621 11611
rect 34621 11577 34655 11611
rect 34655 11577 34664 11611
rect 34612 11568 34664 11577
rect 34888 11500 34940 11552
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 2688 11339 2740 11348
rect 2688 11305 2697 11339
rect 2697 11305 2731 11339
rect 2731 11305 2740 11339
rect 2688 11296 2740 11305
rect 10140 11339 10192 11348
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 15752 11339 15804 11348
rect 15752 11305 15761 11339
rect 15761 11305 15795 11339
rect 15795 11305 15804 11339
rect 15752 11296 15804 11305
rect 27068 11296 27120 11348
rect 31484 11339 31536 11348
rect 31484 11305 31493 11339
rect 31493 11305 31527 11339
rect 31527 11305 31536 11339
rect 31484 11296 31536 11305
rect 35624 11339 35676 11348
rect 35624 11305 35633 11339
rect 35633 11305 35667 11339
rect 35667 11305 35676 11339
rect 35624 11296 35676 11305
rect 11612 11271 11664 11280
rect 11612 11237 11621 11271
rect 11621 11237 11655 11271
rect 11655 11237 11664 11271
rect 11612 11228 11664 11237
rect 20628 11228 20680 11280
rect 24400 11271 24452 11280
rect 24400 11237 24409 11271
rect 24409 11237 24443 11271
rect 24443 11237 24452 11271
rect 24400 11228 24452 11237
rect 24492 11271 24544 11280
rect 24492 11237 24501 11271
rect 24501 11237 24535 11271
rect 24535 11237 24544 11271
rect 24492 11228 24544 11237
rect 29552 11228 29604 11280
rect 29920 11271 29972 11280
rect 29920 11237 29929 11271
rect 29929 11237 29963 11271
rect 29963 11237 29972 11271
rect 29920 11228 29972 11237
rect 1676 11160 1728 11212
rect 3332 11160 3384 11212
rect 4712 11160 4764 11212
rect 8576 11203 8628 11212
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 10416 11203 10468 11212
rect 10416 11169 10425 11203
rect 10425 11169 10459 11203
rect 10459 11169 10468 11203
rect 10416 11160 10468 11169
rect 12992 11203 13044 11212
rect 12992 11169 13001 11203
rect 13001 11169 13035 11203
rect 13035 11169 13044 11203
rect 12992 11160 13044 11169
rect 15476 11203 15528 11212
rect 15476 11169 15485 11203
rect 15485 11169 15519 11203
rect 15519 11169 15528 11203
rect 15476 11160 15528 11169
rect 15568 11160 15620 11212
rect 16488 11160 16540 11212
rect 18328 11160 18380 11212
rect 19156 11203 19208 11212
rect 19156 11169 19165 11203
rect 19165 11169 19199 11203
rect 19199 11169 19208 11203
rect 19156 11160 19208 11169
rect 19616 11203 19668 11212
rect 19616 11169 19625 11203
rect 19625 11169 19659 11203
rect 19659 11169 19668 11203
rect 19616 11160 19668 11169
rect 23112 11160 23164 11212
rect 27068 11160 27120 11212
rect 27528 11160 27580 11212
rect 28080 11160 28132 11212
rect 31392 11160 31444 11212
rect 32496 11160 32548 11212
rect 34152 11160 34204 11212
rect 35440 11203 35492 11212
rect 35440 11169 35449 11203
rect 35449 11169 35483 11203
rect 35483 11169 35492 11203
rect 35440 11160 35492 11169
rect 37004 11160 37056 11212
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 19892 11135 19944 11144
rect 8116 11024 8168 11076
rect 19892 11101 19901 11135
rect 19901 11101 19935 11135
rect 19935 11101 19944 11135
rect 19892 11092 19944 11101
rect 21456 11092 21508 11144
rect 21640 11135 21692 11144
rect 21640 11101 21649 11135
rect 21649 11101 21683 11135
rect 21683 11101 21692 11135
rect 21640 11092 21692 11101
rect 25228 11092 25280 11144
rect 29644 11092 29696 11144
rect 32680 11135 32732 11144
rect 32680 11101 32689 11135
rect 32689 11101 32723 11135
rect 32723 11101 32732 11135
rect 32680 11092 32732 11101
rect 35072 11092 35124 11144
rect 12072 11067 12124 11076
rect 12072 11033 12081 11067
rect 12081 11033 12115 11067
rect 12115 11033 12124 11067
rect 12072 11024 12124 11033
rect 13176 11067 13228 11076
rect 13176 11033 13185 11067
rect 13185 11033 13219 11067
rect 13219 11033 13228 11067
rect 13176 11024 13228 11033
rect 30564 11024 30616 11076
rect 33692 11024 33744 11076
rect 34428 11024 34480 11076
rect 39580 11024 39632 11076
rect 1584 10999 1636 11008
rect 1584 10965 1593 10999
rect 1593 10965 1627 10999
rect 1627 10965 1636 10999
rect 1584 10956 1636 10965
rect 3792 10956 3844 11008
rect 10048 10956 10100 11008
rect 10232 10956 10284 11008
rect 12440 10999 12492 11008
rect 12440 10965 12449 10999
rect 12449 10965 12483 10999
rect 12483 10965 12492 10999
rect 12440 10956 12492 10965
rect 17592 10956 17644 11008
rect 20168 10999 20220 11008
rect 20168 10965 20177 10999
rect 20177 10965 20211 10999
rect 20211 10965 20220 10999
rect 20168 10956 20220 10965
rect 23020 10956 23072 11008
rect 28080 10956 28132 11008
rect 34980 10956 35032 11008
rect 36728 10999 36780 11008
rect 36728 10965 36737 10999
rect 36737 10965 36771 10999
rect 36771 10965 36780 10999
rect 36728 10956 36780 10965
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 4712 10795 4764 10804
rect 4712 10761 4721 10795
rect 4721 10761 4755 10795
rect 4755 10761 4764 10795
rect 4712 10752 4764 10761
rect 8300 10795 8352 10804
rect 8300 10761 8309 10795
rect 8309 10761 8343 10795
rect 8343 10761 8352 10795
rect 8300 10752 8352 10761
rect 11612 10752 11664 10804
rect 11704 10752 11756 10804
rect 16488 10752 16540 10804
rect 17132 10752 17184 10804
rect 18328 10795 18380 10804
rect 18328 10761 18337 10795
rect 18337 10761 18371 10795
rect 18371 10761 18380 10795
rect 18328 10752 18380 10761
rect 21456 10795 21508 10804
rect 21456 10761 21465 10795
rect 21465 10761 21499 10795
rect 21499 10761 21508 10795
rect 21456 10752 21508 10761
rect 23480 10752 23532 10804
rect 24400 10752 24452 10804
rect 27068 10795 27120 10804
rect 27068 10761 27077 10795
rect 27077 10761 27111 10795
rect 27111 10761 27120 10795
rect 27068 10752 27120 10761
rect 29552 10752 29604 10804
rect 31760 10752 31812 10804
rect 34152 10752 34204 10804
rect 36636 10795 36688 10804
rect 36636 10761 36645 10795
rect 36645 10761 36679 10795
rect 36679 10761 36688 10795
rect 36636 10752 36688 10761
rect 37004 10795 37056 10804
rect 37004 10761 37013 10795
rect 37013 10761 37047 10795
rect 37047 10761 37056 10795
rect 37004 10752 37056 10761
rect 2412 10684 2464 10736
rect 2136 10548 2188 10600
rect 112 10412 164 10464
rect 2044 10455 2096 10464
rect 2044 10421 2053 10455
rect 2053 10421 2087 10455
rect 2087 10421 2096 10455
rect 2044 10412 2096 10421
rect 3424 10480 3476 10532
rect 3148 10412 3200 10464
rect 3332 10455 3384 10464
rect 3332 10421 3341 10455
rect 3341 10421 3375 10455
rect 3375 10421 3384 10455
rect 3332 10412 3384 10421
rect 3884 10412 3936 10464
rect 8208 10548 8260 10600
rect 10416 10684 10468 10736
rect 11520 10616 11572 10668
rect 12992 10684 13044 10736
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 13176 10616 13228 10668
rect 19156 10684 19208 10736
rect 21272 10684 21324 10736
rect 15384 10659 15436 10668
rect 15384 10625 15393 10659
rect 15393 10625 15427 10659
rect 15427 10625 15436 10659
rect 15384 10616 15436 10625
rect 14188 10548 14240 10600
rect 19524 10616 19576 10668
rect 19708 10616 19760 10668
rect 20076 10659 20128 10668
rect 20076 10625 20085 10659
rect 20085 10625 20119 10659
rect 20119 10625 20128 10659
rect 20076 10616 20128 10625
rect 21640 10616 21692 10668
rect 24584 10659 24636 10668
rect 24584 10625 24593 10659
rect 24593 10625 24627 10659
rect 24627 10625 24636 10659
rect 24584 10616 24636 10625
rect 10232 10523 10284 10532
rect 10232 10489 10241 10523
rect 10241 10489 10275 10523
rect 10275 10489 10284 10523
rect 10232 10480 10284 10489
rect 10324 10523 10376 10532
rect 10324 10489 10333 10523
rect 10333 10489 10367 10523
rect 10367 10489 10376 10523
rect 10324 10480 10376 10489
rect 11060 10480 11112 10532
rect 15108 10523 15160 10532
rect 15108 10489 15117 10523
rect 15117 10489 15151 10523
rect 15151 10489 15160 10523
rect 15108 10480 15160 10489
rect 15200 10523 15252 10532
rect 15200 10489 15209 10523
rect 15209 10489 15243 10523
rect 15243 10489 15252 10523
rect 15200 10480 15252 10489
rect 15476 10480 15528 10532
rect 19156 10523 19208 10532
rect 19156 10489 19165 10523
rect 19165 10489 19199 10523
rect 19199 10489 19208 10523
rect 19156 10480 19208 10489
rect 4344 10455 4396 10464
rect 4344 10421 4353 10455
rect 4353 10421 4387 10455
rect 4387 10421 4396 10455
rect 4344 10412 4396 10421
rect 6552 10412 6604 10464
rect 7288 10412 7340 10464
rect 8576 10412 8628 10464
rect 9680 10455 9732 10464
rect 9680 10421 9689 10455
rect 9689 10421 9723 10455
rect 9723 10421 9732 10455
rect 9680 10412 9732 10421
rect 12532 10455 12584 10464
rect 12532 10421 12541 10455
rect 12541 10421 12575 10455
rect 12575 10421 12584 10455
rect 12532 10412 12584 10421
rect 14832 10412 14884 10464
rect 21456 10548 21508 10600
rect 22836 10548 22888 10600
rect 29460 10684 29512 10736
rect 29920 10684 29972 10736
rect 30564 10727 30616 10736
rect 30564 10693 30573 10727
rect 30573 10693 30607 10727
rect 30607 10693 30616 10727
rect 30564 10684 30616 10693
rect 31484 10684 31536 10736
rect 20168 10523 20220 10532
rect 20168 10489 20177 10523
rect 20177 10489 20211 10523
rect 20211 10489 20220 10523
rect 20168 10480 20220 10489
rect 19708 10412 19760 10464
rect 20628 10412 20680 10464
rect 21732 10455 21784 10464
rect 21732 10421 21741 10455
rect 21741 10421 21775 10455
rect 21775 10421 21784 10455
rect 21732 10412 21784 10421
rect 23296 10480 23348 10532
rect 24584 10480 24636 10532
rect 25228 10523 25280 10532
rect 25228 10489 25237 10523
rect 25237 10489 25271 10523
rect 25271 10489 25280 10523
rect 25228 10480 25280 10489
rect 26240 10548 26292 10600
rect 30012 10616 30064 10668
rect 34060 10684 34112 10736
rect 32496 10616 32548 10668
rect 33324 10616 33376 10668
rect 28080 10591 28132 10600
rect 28080 10557 28089 10591
rect 28089 10557 28123 10591
rect 28123 10557 28132 10591
rect 28080 10548 28132 10557
rect 32956 10591 33008 10600
rect 32956 10557 32965 10591
rect 32965 10557 32999 10591
rect 32999 10557 33008 10591
rect 34152 10616 34204 10668
rect 35440 10616 35492 10668
rect 32956 10548 33008 10557
rect 33784 10591 33836 10600
rect 33784 10557 33793 10591
rect 33793 10557 33827 10591
rect 33827 10557 33836 10591
rect 33784 10548 33836 10557
rect 28356 10523 28408 10532
rect 28356 10489 28365 10523
rect 28365 10489 28399 10523
rect 28399 10489 28408 10523
rect 28356 10480 28408 10489
rect 23112 10412 23164 10464
rect 24400 10455 24452 10464
rect 24400 10421 24409 10455
rect 24409 10421 24443 10455
rect 24443 10421 24452 10455
rect 24400 10412 24452 10421
rect 26148 10455 26200 10464
rect 26148 10421 26157 10455
rect 26157 10421 26191 10455
rect 26191 10421 26200 10455
rect 26148 10412 26200 10421
rect 27528 10412 27580 10464
rect 30104 10523 30156 10532
rect 30104 10489 30113 10523
rect 30113 10489 30147 10523
rect 30147 10489 30156 10523
rect 30104 10480 30156 10489
rect 30656 10480 30708 10532
rect 31392 10480 31444 10532
rect 31668 10523 31720 10532
rect 31668 10489 31677 10523
rect 31677 10489 31711 10523
rect 31711 10489 31720 10523
rect 31668 10480 31720 10489
rect 32220 10523 32272 10532
rect 32220 10489 32229 10523
rect 32229 10489 32263 10523
rect 32263 10489 32272 10523
rect 32220 10480 32272 10489
rect 32312 10480 32364 10532
rect 34980 10523 35032 10532
rect 34980 10489 34989 10523
rect 34989 10489 35023 10523
rect 35023 10489 35032 10523
rect 34980 10480 35032 10489
rect 35072 10523 35124 10532
rect 35072 10489 35081 10523
rect 35081 10489 35115 10523
rect 35115 10489 35124 10523
rect 35624 10523 35676 10532
rect 35072 10480 35124 10489
rect 35624 10489 35633 10523
rect 35633 10489 35667 10523
rect 35667 10489 35676 10523
rect 35624 10480 35676 10489
rect 31116 10412 31168 10464
rect 32496 10455 32548 10464
rect 32496 10421 32505 10455
rect 32505 10421 32539 10455
rect 32539 10421 32548 10455
rect 32496 10412 32548 10421
rect 34612 10412 34664 10464
rect 36084 10412 36136 10464
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 1768 10208 1820 10260
rect 2780 10208 2832 10260
rect 10324 10251 10376 10260
rect 10324 10217 10333 10251
rect 10333 10217 10367 10251
rect 10367 10217 10376 10251
rect 10324 10208 10376 10217
rect 11612 10208 11664 10260
rect 10600 10183 10652 10192
rect 10600 10149 10609 10183
rect 10609 10149 10643 10183
rect 10643 10149 10652 10183
rect 10600 10140 10652 10149
rect 11428 10140 11480 10192
rect 13636 10208 13688 10260
rect 1492 10072 1544 10124
rect 2412 10115 2464 10124
rect 2412 10081 2421 10115
rect 2421 10081 2455 10115
rect 2455 10081 2464 10115
rect 2412 10072 2464 10081
rect 5172 10072 5224 10124
rect 8024 10072 8076 10124
rect 8392 10072 8444 10124
rect 13820 10072 13872 10124
rect 15568 10183 15620 10192
rect 15568 10149 15577 10183
rect 15577 10149 15611 10183
rect 15611 10149 15620 10183
rect 16028 10183 16080 10192
rect 15568 10140 15620 10149
rect 14188 10115 14240 10124
rect 14188 10081 14197 10115
rect 14197 10081 14231 10115
rect 14231 10081 14240 10115
rect 16028 10149 16037 10183
rect 16037 10149 16071 10183
rect 16071 10149 16080 10183
rect 16028 10140 16080 10149
rect 19156 10208 19208 10260
rect 19248 10251 19300 10260
rect 19248 10217 19257 10251
rect 19257 10217 19291 10251
rect 19291 10217 19300 10251
rect 19248 10208 19300 10217
rect 20076 10208 20128 10260
rect 17684 10115 17736 10124
rect 14188 10072 14240 10081
rect 17684 10081 17693 10115
rect 17693 10081 17727 10115
rect 17727 10081 17736 10115
rect 17684 10072 17736 10081
rect 18144 10115 18196 10124
rect 18144 10081 18153 10115
rect 18153 10081 18187 10115
rect 18187 10081 18196 10115
rect 18144 10072 18196 10081
rect 21916 10140 21968 10192
rect 19524 10072 19576 10124
rect 19708 10115 19760 10124
rect 19708 10081 19717 10115
rect 19717 10081 19751 10115
rect 19751 10081 19760 10115
rect 19708 10072 19760 10081
rect 21640 10115 21692 10124
rect 21640 10081 21649 10115
rect 21649 10081 21683 10115
rect 21683 10081 21692 10115
rect 21640 10072 21692 10081
rect 9588 10004 9640 10056
rect 10508 10047 10560 10056
rect 10508 10013 10517 10047
rect 10517 10013 10551 10047
rect 10551 10013 10560 10047
rect 10508 10004 10560 10013
rect 12348 10047 12400 10056
rect 12348 10013 12357 10047
rect 12357 10013 12391 10047
rect 12391 10013 12400 10047
rect 12348 10004 12400 10013
rect 15108 10004 15160 10056
rect 15936 10047 15988 10056
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 18328 10047 18380 10056
rect 10968 9936 11020 9988
rect 11060 9979 11112 9988
rect 11060 9945 11069 9979
rect 11069 9945 11103 9979
rect 11103 9945 11112 9979
rect 11060 9936 11112 9945
rect 12072 9936 12124 9988
rect 13176 9936 13228 9988
rect 15384 9936 15436 9988
rect 18328 10013 18337 10047
rect 18337 10013 18371 10047
rect 18371 10013 18380 10047
rect 18328 10004 18380 10013
rect 20720 10004 20772 10056
rect 25228 10208 25280 10260
rect 29460 10251 29512 10260
rect 23204 10140 23256 10192
rect 24584 10140 24636 10192
rect 24768 10183 24820 10192
rect 24768 10149 24777 10183
rect 24777 10149 24811 10183
rect 24811 10149 24820 10183
rect 24768 10140 24820 10149
rect 24860 10183 24912 10192
rect 24860 10149 24869 10183
rect 24869 10149 24903 10183
rect 24903 10149 24912 10183
rect 29460 10217 29469 10251
rect 29469 10217 29503 10251
rect 29503 10217 29512 10251
rect 29460 10208 29512 10217
rect 29644 10208 29696 10260
rect 31668 10208 31720 10260
rect 32680 10251 32732 10260
rect 32680 10217 32689 10251
rect 32689 10217 32723 10251
rect 32723 10217 32732 10251
rect 32680 10208 32732 10217
rect 24860 10140 24912 10149
rect 25964 10140 26016 10192
rect 28632 10140 28684 10192
rect 30288 10140 30340 10192
rect 30564 10183 30616 10192
rect 30564 10149 30573 10183
rect 30573 10149 30607 10183
rect 30607 10149 30616 10183
rect 30564 10140 30616 10149
rect 32220 10140 32272 10192
rect 36268 10251 36320 10260
rect 36268 10217 36277 10251
rect 36277 10217 36311 10251
rect 36311 10217 36320 10251
rect 36268 10208 36320 10217
rect 33140 10183 33192 10192
rect 33140 10149 33149 10183
rect 33149 10149 33183 10183
rect 33183 10149 33192 10183
rect 33692 10183 33744 10192
rect 33140 10140 33192 10149
rect 33692 10149 33701 10183
rect 33701 10149 33735 10183
rect 33735 10149 33744 10183
rect 33692 10140 33744 10149
rect 34704 10183 34756 10192
rect 34704 10149 34713 10183
rect 34713 10149 34747 10183
rect 34747 10149 34756 10183
rect 34704 10140 34756 10149
rect 34888 10140 34940 10192
rect 36544 10140 36596 10192
rect 26240 10072 26292 10124
rect 36084 10115 36136 10124
rect 36084 10081 36093 10115
rect 36093 10081 36127 10115
rect 36127 10081 36136 10115
rect 36084 10072 36136 10081
rect 23020 10004 23072 10056
rect 23480 10047 23532 10056
rect 23480 10013 23489 10047
rect 23489 10013 23523 10047
rect 23523 10013 23532 10047
rect 23480 10004 23532 10013
rect 26332 10004 26384 10056
rect 28540 10047 28592 10056
rect 25780 9936 25832 9988
rect 28540 10013 28549 10047
rect 28549 10013 28583 10047
rect 28583 10013 28592 10047
rect 28540 10004 28592 10013
rect 31116 10047 31168 10056
rect 31116 10013 31125 10047
rect 31125 10013 31159 10047
rect 31159 10013 31168 10047
rect 34612 10047 34664 10056
rect 31116 10004 31168 10013
rect 32496 9936 32548 9988
rect 34612 10013 34621 10047
rect 34621 10013 34655 10047
rect 34655 10013 34664 10047
rect 34612 10004 34664 10013
rect 35256 9936 35308 9988
rect 1676 9911 1728 9920
rect 1676 9877 1685 9911
rect 1685 9877 1719 9911
rect 1719 9877 1728 9911
rect 1676 9868 1728 9877
rect 8852 9868 8904 9920
rect 9036 9911 9088 9920
rect 9036 9877 9045 9911
rect 9045 9877 9079 9911
rect 9079 9877 9088 9911
rect 9036 9868 9088 9877
rect 10048 9868 10100 9920
rect 16120 9868 16172 9920
rect 23664 9868 23716 9920
rect 24400 9868 24452 9920
rect 25964 9868 26016 9920
rect 27068 9868 27120 9920
rect 28080 9868 28132 9920
rect 30104 9911 30156 9920
rect 30104 9877 30113 9911
rect 30113 9877 30147 9911
rect 30147 9877 30156 9911
rect 30104 9868 30156 9877
rect 35624 9868 35676 9920
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 2412 9664 2464 9716
rect 5172 9707 5224 9716
rect 5172 9673 5181 9707
rect 5181 9673 5215 9707
rect 5215 9673 5224 9707
rect 5172 9664 5224 9673
rect 5908 9664 5960 9716
rect 8852 9664 8904 9716
rect 10508 9664 10560 9716
rect 11428 9707 11480 9716
rect 11428 9673 11437 9707
rect 11437 9673 11471 9707
rect 11471 9673 11480 9707
rect 11428 9664 11480 9673
rect 11612 9664 11664 9716
rect 16028 9664 16080 9716
rect 16672 9664 16724 9716
rect 18144 9664 18196 9716
rect 18788 9707 18840 9716
rect 18788 9673 18797 9707
rect 18797 9673 18831 9707
rect 18831 9673 18840 9707
rect 18788 9664 18840 9673
rect 20168 9707 20220 9716
rect 20168 9673 20177 9707
rect 20177 9673 20211 9707
rect 20211 9673 20220 9707
rect 20168 9664 20220 9673
rect 21916 9707 21968 9716
rect 21916 9673 21925 9707
rect 21925 9673 21959 9707
rect 21959 9673 21968 9707
rect 21916 9664 21968 9673
rect 23020 9664 23072 9716
rect 23204 9664 23256 9716
rect 24584 9707 24636 9716
rect 24584 9673 24593 9707
rect 24593 9673 24627 9707
rect 24627 9673 24636 9707
rect 24584 9664 24636 9673
rect 24860 9707 24912 9716
rect 24860 9673 24869 9707
rect 24869 9673 24903 9707
rect 24903 9673 24912 9707
rect 24860 9664 24912 9673
rect 25964 9664 26016 9716
rect 30288 9664 30340 9716
rect 32312 9664 32364 9716
rect 33140 9664 33192 9716
rect 34612 9664 34664 9716
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 7380 9596 7432 9648
rect 12348 9596 12400 9648
rect 8484 9528 8536 9580
rect 9036 9528 9088 9580
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 10968 9528 11020 9580
rect 12256 9528 12308 9580
rect 14188 9596 14240 9648
rect 15936 9596 15988 9648
rect 23296 9596 23348 9648
rect 26332 9596 26384 9648
rect 27068 9639 27120 9648
rect 27068 9605 27077 9639
rect 27077 9605 27111 9639
rect 27111 9605 27120 9639
rect 27068 9596 27120 9605
rect 30564 9639 30616 9648
rect 30564 9605 30573 9639
rect 30573 9605 30607 9639
rect 30607 9605 30616 9639
rect 30564 9596 30616 9605
rect 13636 9528 13688 9580
rect 15016 9571 15068 9580
rect 15016 9537 15025 9571
rect 15025 9537 15059 9571
rect 15059 9537 15068 9571
rect 15016 9528 15068 9537
rect 19156 9528 19208 9580
rect 19892 9528 19944 9580
rect 21824 9528 21876 9580
rect 23664 9571 23716 9580
rect 2412 9435 2464 9444
rect 2412 9401 2421 9435
rect 2421 9401 2455 9435
rect 2455 9401 2464 9435
rect 2412 9392 2464 9401
rect 3056 9392 3108 9444
rect 5908 9460 5960 9512
rect 6000 9460 6052 9512
rect 7380 9503 7432 9512
rect 7380 9469 7389 9503
rect 7389 9469 7423 9503
rect 7423 9469 7432 9503
rect 7380 9460 7432 9469
rect 10324 9460 10376 9512
rect 7196 9392 7248 9444
rect 7472 9392 7524 9444
rect 8392 9435 8444 9444
rect 8392 9401 8401 9435
rect 8401 9401 8435 9435
rect 8435 9401 8444 9435
rect 8392 9392 8444 9401
rect 8760 9435 8812 9444
rect 8760 9401 8769 9435
rect 8769 9401 8803 9435
rect 8803 9401 8812 9435
rect 8760 9392 8812 9401
rect 1492 9324 1544 9376
rect 4068 9324 4120 9376
rect 6736 9324 6788 9376
rect 7840 9367 7892 9376
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 9772 9324 9824 9376
rect 13544 9460 13596 9512
rect 15200 9460 15252 9512
rect 17500 9460 17552 9512
rect 18788 9460 18840 9512
rect 23020 9460 23072 9512
rect 23664 9537 23673 9571
rect 23673 9537 23707 9571
rect 23707 9537 23716 9571
rect 23664 9528 23716 9537
rect 24676 9528 24728 9580
rect 25504 9571 25556 9580
rect 25504 9537 25513 9571
rect 25513 9537 25547 9571
rect 25547 9537 25556 9571
rect 25504 9528 25556 9537
rect 25780 9571 25832 9580
rect 25780 9537 25789 9571
rect 25789 9537 25823 9571
rect 25823 9537 25832 9571
rect 25780 9528 25832 9537
rect 28540 9528 28592 9580
rect 29644 9528 29696 9580
rect 32680 9528 32732 9580
rect 34796 9528 34848 9580
rect 35256 9571 35308 9580
rect 35256 9537 35265 9571
rect 35265 9537 35299 9571
rect 35299 9537 35308 9571
rect 35256 9528 35308 9537
rect 35624 9528 35676 9580
rect 28080 9503 28132 9512
rect 15844 9392 15896 9444
rect 21364 9435 21416 9444
rect 21364 9401 21367 9435
rect 21367 9401 21401 9435
rect 21401 9401 21416 9435
rect 21364 9392 21416 9401
rect 23664 9392 23716 9444
rect 28080 9469 28089 9503
rect 28089 9469 28123 9503
rect 28123 9469 28132 9503
rect 28080 9460 28132 9469
rect 31760 9503 31812 9512
rect 13912 9324 13964 9376
rect 17316 9324 17368 9376
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 18604 9324 18656 9376
rect 19524 9324 19576 9376
rect 21732 9324 21784 9376
rect 24860 9324 24912 9376
rect 28264 9392 28316 9444
rect 28632 9324 28684 9376
rect 28816 9324 28868 9376
rect 30748 9392 30800 9444
rect 31760 9469 31769 9503
rect 31769 9469 31803 9503
rect 31803 9469 31812 9503
rect 31760 9460 31812 9469
rect 32036 9324 32088 9376
rect 35072 9435 35124 9444
rect 35072 9401 35081 9435
rect 35081 9401 35115 9435
rect 35115 9401 35124 9435
rect 35072 9392 35124 9401
rect 36360 9392 36412 9444
rect 36544 9435 36596 9444
rect 36544 9401 36553 9435
rect 36553 9401 36587 9435
rect 36587 9401 36596 9435
rect 36544 9392 36596 9401
rect 36636 9435 36688 9444
rect 36636 9401 36645 9435
rect 36645 9401 36679 9435
rect 36679 9401 36688 9435
rect 36636 9392 36688 9401
rect 34336 9367 34388 9376
rect 34336 9333 34345 9367
rect 34345 9333 34379 9367
rect 34379 9333 34388 9367
rect 34336 9324 34388 9333
rect 36084 9367 36136 9376
rect 36084 9333 36093 9367
rect 36093 9333 36127 9367
rect 36127 9333 36136 9367
rect 36084 9324 36136 9333
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 1676 9120 1728 9172
rect 2596 9095 2648 9104
rect 2596 9061 2605 9095
rect 2605 9061 2639 9095
rect 2639 9061 2648 9095
rect 2596 9052 2648 9061
rect 5080 9095 5132 9104
rect 5080 9061 5089 9095
rect 5089 9061 5123 9095
rect 5123 9061 5132 9095
rect 5080 9052 5132 9061
rect 6552 9095 6604 9104
rect 6552 9061 6561 9095
rect 6561 9061 6595 9095
rect 6595 9061 6604 9095
rect 6552 9052 6604 9061
rect 6644 9095 6696 9104
rect 6644 9061 6653 9095
rect 6653 9061 6687 9095
rect 6687 9061 6696 9095
rect 6920 9120 6972 9172
rect 10140 9163 10192 9172
rect 10140 9129 10149 9163
rect 10149 9129 10183 9163
rect 10183 9129 10192 9163
rect 10140 9120 10192 9129
rect 10784 9120 10836 9172
rect 11428 9163 11480 9172
rect 11428 9129 11437 9163
rect 11437 9129 11471 9163
rect 11471 9129 11480 9163
rect 11428 9120 11480 9129
rect 11612 9120 11664 9172
rect 12256 9120 12308 9172
rect 15016 9163 15068 9172
rect 15016 9129 15025 9163
rect 15025 9129 15059 9163
rect 15059 9129 15068 9163
rect 15016 9120 15068 9129
rect 16672 9163 16724 9172
rect 16672 9129 16681 9163
rect 16681 9129 16715 9163
rect 16715 9129 16724 9163
rect 16672 9120 16724 9129
rect 17684 9163 17736 9172
rect 17684 9129 17693 9163
rect 17693 9129 17727 9163
rect 17727 9129 17736 9163
rect 17684 9120 17736 9129
rect 18604 9120 18656 9172
rect 20720 9163 20772 9172
rect 6644 9052 6696 9061
rect 1676 8984 1728 9036
rect 8116 9027 8168 9036
rect 8116 8993 8125 9027
rect 8125 8993 8159 9027
rect 8159 8993 8168 9027
rect 8116 8984 8168 8993
rect 8484 9027 8536 9036
rect 8484 8993 8493 9027
rect 8493 8993 8527 9027
rect 8527 8993 8536 9027
rect 8484 8984 8536 8993
rect 10232 9052 10284 9104
rect 13820 9095 13872 9104
rect 13820 9061 13829 9095
rect 13829 9061 13863 9095
rect 13863 9061 13872 9095
rect 13820 9052 13872 9061
rect 15384 9052 15436 9104
rect 15844 9052 15896 9104
rect 20720 9129 20729 9163
rect 20729 9129 20763 9163
rect 20763 9129 20772 9163
rect 20720 9120 20772 9129
rect 21824 9163 21876 9172
rect 21824 9129 21833 9163
rect 21833 9129 21867 9163
rect 21867 9129 21876 9163
rect 21824 9120 21876 9129
rect 24768 9120 24820 9172
rect 25136 9120 25188 9172
rect 28540 9163 28592 9172
rect 28540 9129 28549 9163
rect 28549 9129 28583 9163
rect 28583 9129 28592 9163
rect 28540 9120 28592 9129
rect 30104 9120 30156 9172
rect 34060 9163 34112 9172
rect 34060 9129 34069 9163
rect 34069 9129 34103 9163
rect 34103 9129 34112 9163
rect 34060 9120 34112 9129
rect 34796 9120 34848 9172
rect 35808 9163 35860 9172
rect 35808 9129 35817 9163
rect 35817 9129 35851 9163
rect 35851 9129 35860 9163
rect 35808 9120 35860 9129
rect 36360 9163 36412 9172
rect 36360 9129 36369 9163
rect 36369 9129 36403 9163
rect 36403 9129 36412 9163
rect 36360 9120 36412 9129
rect 36636 9163 36688 9172
rect 36636 9129 36645 9163
rect 36645 9129 36679 9163
rect 36679 9129 36688 9163
rect 36636 9120 36688 9129
rect 19064 9095 19116 9104
rect 19064 9061 19073 9095
rect 19073 9061 19107 9095
rect 19107 9061 19116 9095
rect 19064 9052 19116 9061
rect 19708 9052 19760 9104
rect 23020 9095 23072 9104
rect 9956 8984 10008 9036
rect 11704 8984 11756 9036
rect 15752 9027 15804 9036
rect 15752 8993 15761 9027
rect 15761 8993 15795 9027
rect 15795 8993 15804 9027
rect 15752 8984 15804 8993
rect 17960 8984 18012 9036
rect 20812 8984 20864 9036
rect 22468 9027 22520 9036
rect 22468 8993 22477 9027
rect 22477 8993 22511 9027
rect 22511 8993 22520 9027
rect 22468 8984 22520 8993
rect 23020 9061 23029 9095
rect 23029 9061 23063 9095
rect 23063 9061 23072 9095
rect 23020 9052 23072 9061
rect 23664 9052 23716 9104
rect 25504 9095 25556 9104
rect 25504 9061 25513 9095
rect 25513 9061 25547 9095
rect 25547 9061 25556 9095
rect 25504 9052 25556 9061
rect 26332 9095 26384 9104
rect 26332 9061 26341 9095
rect 26341 9061 26375 9095
rect 26375 9061 26384 9095
rect 26332 9052 26384 9061
rect 28816 9052 28868 9104
rect 32772 9052 32824 9104
rect 22928 8984 22980 9036
rect 24860 8984 24912 9036
rect 26516 9027 26568 9036
rect 26516 8993 26525 9027
rect 26525 8993 26559 9027
rect 26559 8993 26568 9027
rect 26516 8984 26568 8993
rect 27068 9027 27120 9036
rect 27068 8993 27077 9027
rect 27077 8993 27111 9027
rect 27111 8993 27120 9027
rect 27068 8984 27120 8993
rect 28356 8984 28408 9036
rect 30564 9027 30616 9036
rect 30564 8993 30573 9027
rect 30573 8993 30607 9027
rect 30607 8993 30616 9027
rect 30564 8984 30616 8993
rect 30932 9027 30984 9036
rect 30932 8993 30941 9027
rect 30941 8993 30975 9027
rect 30975 8993 30984 9027
rect 30932 8984 30984 8993
rect 32128 9027 32180 9036
rect 32128 8993 32137 9027
rect 32137 8993 32171 9027
rect 32171 8993 32180 9027
rect 32128 8984 32180 8993
rect 32404 8984 32456 9036
rect 33324 8984 33376 9036
rect 34336 8984 34388 9036
rect 34704 8984 34756 9036
rect 2504 8959 2556 8968
rect 2504 8925 2513 8959
rect 2513 8925 2547 8959
rect 2547 8925 2556 8959
rect 2504 8916 2556 8925
rect 2964 8916 3016 8968
rect 4804 8916 4856 8968
rect 5172 8916 5224 8968
rect 11060 8959 11112 8968
rect 11060 8925 11069 8959
rect 11069 8925 11103 8959
rect 11103 8925 11112 8959
rect 11060 8916 11112 8925
rect 13176 8916 13228 8968
rect 25136 8916 25188 8968
rect 33784 8916 33836 8968
rect 36268 8916 36320 8968
rect 2044 8848 2096 8900
rect 1860 8823 1912 8832
rect 1860 8789 1869 8823
rect 1869 8789 1903 8823
rect 1903 8789 1912 8823
rect 1860 8780 1912 8789
rect 2320 8823 2372 8832
rect 2320 8789 2329 8823
rect 2329 8789 2363 8823
rect 2363 8789 2372 8823
rect 2320 8780 2372 8789
rect 5540 8848 5592 8900
rect 7840 8848 7892 8900
rect 19524 8891 19576 8900
rect 19524 8857 19533 8891
rect 19533 8857 19567 8891
rect 19567 8857 19576 8891
rect 19524 8848 19576 8857
rect 33416 8848 33468 8900
rect 39580 8848 39632 8900
rect 4712 8780 4764 8832
rect 8760 8780 8812 8832
rect 10600 8823 10652 8832
rect 10600 8789 10609 8823
rect 10609 8789 10643 8823
rect 10643 8789 10652 8823
rect 10600 8780 10652 8789
rect 12808 8823 12860 8832
rect 12808 8789 12817 8823
rect 12817 8789 12851 8823
rect 12851 8789 12860 8823
rect 12808 8780 12860 8789
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 13728 8780 13780 8832
rect 18236 8780 18288 8832
rect 18420 8823 18472 8832
rect 18420 8789 18429 8823
rect 18429 8789 18463 8823
rect 18463 8789 18472 8823
rect 18420 8780 18472 8789
rect 20720 8780 20772 8832
rect 21548 8823 21600 8832
rect 21548 8789 21557 8823
rect 21557 8789 21591 8823
rect 21591 8789 21600 8823
rect 21548 8780 21600 8789
rect 23664 8823 23716 8832
rect 23664 8789 23673 8823
rect 23673 8789 23707 8823
rect 23707 8789 23716 8823
rect 23664 8780 23716 8789
rect 27712 8823 27764 8832
rect 27712 8789 27721 8823
rect 27721 8789 27755 8823
rect 27755 8789 27764 8823
rect 27712 8780 27764 8789
rect 30196 8780 30248 8832
rect 34980 8823 35032 8832
rect 34980 8789 34989 8823
rect 34989 8789 35023 8823
rect 35023 8789 35032 8823
rect 34980 8780 35032 8789
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 1676 8619 1728 8628
rect 1676 8585 1685 8619
rect 1685 8585 1719 8619
rect 1719 8585 1728 8619
rect 1676 8576 1728 8585
rect 2596 8576 2648 8628
rect 3148 8576 3200 8628
rect 3976 8619 4028 8628
rect 3976 8585 3985 8619
rect 3985 8585 4019 8619
rect 4019 8585 4028 8619
rect 3976 8576 4028 8585
rect 6552 8576 6604 8628
rect 8116 8619 8168 8628
rect 8116 8585 8125 8619
rect 8125 8585 8159 8619
rect 8159 8585 8168 8619
rect 8116 8576 8168 8585
rect 8484 8619 8536 8628
rect 8484 8585 8493 8619
rect 8493 8585 8527 8619
rect 8527 8585 8536 8619
rect 8484 8576 8536 8585
rect 9036 8576 9088 8628
rect 9956 8619 10008 8628
rect 9956 8585 9965 8619
rect 9965 8585 9999 8619
rect 9999 8585 10008 8619
rect 9956 8576 10008 8585
rect 10600 8576 10652 8628
rect 11060 8576 11112 8628
rect 12532 8576 12584 8628
rect 13820 8576 13872 8628
rect 15752 8576 15804 8628
rect 19248 8619 19300 8628
rect 19248 8585 19257 8619
rect 19257 8585 19291 8619
rect 19291 8585 19300 8619
rect 19248 8576 19300 8585
rect 20628 8619 20680 8628
rect 20628 8585 20637 8619
rect 20637 8585 20671 8619
rect 20671 8585 20680 8619
rect 20628 8576 20680 8585
rect 20812 8576 20864 8628
rect 21272 8619 21324 8628
rect 21272 8585 21281 8619
rect 21281 8585 21315 8619
rect 21315 8585 21324 8619
rect 21272 8576 21324 8585
rect 24400 8576 24452 8628
rect 25136 8576 25188 8628
rect 25412 8576 25464 8628
rect 27068 8619 27120 8628
rect 2504 8508 2556 8560
rect 5172 8508 5224 8560
rect 1860 8440 1912 8492
rect 2964 8483 3016 8492
rect 2964 8449 2973 8483
rect 2973 8449 3007 8483
rect 3007 8449 3016 8483
rect 2964 8440 3016 8449
rect 5448 8440 5500 8492
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 10784 8440 10836 8492
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 4620 8372 4672 8424
rect 2320 8304 2372 8356
rect 2688 8304 2740 8356
rect 5356 8347 5408 8356
rect 5356 8313 5365 8347
rect 5365 8313 5399 8347
rect 5399 8313 5408 8347
rect 5356 8304 5408 8313
rect 9496 8415 9548 8424
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 11244 8372 11296 8424
rect 12808 8415 12860 8424
rect 12808 8381 12817 8415
rect 12817 8381 12851 8415
rect 12851 8381 12860 8415
rect 12808 8372 12860 8381
rect 14648 8372 14700 8424
rect 17132 8440 17184 8492
rect 16856 8415 16908 8424
rect 16856 8381 16865 8415
rect 16865 8381 16899 8415
rect 16899 8381 16908 8415
rect 16856 8372 16908 8381
rect 4712 8236 4764 8288
rect 7196 8304 7248 8356
rect 9772 8304 9824 8356
rect 11428 8304 11480 8356
rect 6828 8236 6880 8288
rect 17040 8347 17092 8356
rect 17040 8313 17049 8347
rect 17049 8313 17083 8347
rect 17083 8313 17092 8347
rect 17040 8304 17092 8313
rect 17316 8440 17368 8492
rect 18512 8440 18564 8492
rect 18604 8483 18656 8492
rect 18604 8449 18613 8483
rect 18613 8449 18647 8483
rect 18647 8449 18656 8483
rect 18604 8440 18656 8449
rect 27068 8585 27077 8619
rect 27077 8585 27111 8619
rect 27111 8585 27120 8619
rect 27068 8576 27120 8585
rect 28356 8576 28408 8628
rect 31208 8576 31260 8628
rect 34060 8619 34112 8628
rect 34060 8585 34069 8619
rect 34069 8585 34103 8619
rect 34103 8585 34112 8619
rect 34060 8576 34112 8585
rect 35808 8576 35860 8628
rect 36268 8619 36320 8628
rect 36268 8585 36277 8619
rect 36277 8585 36311 8619
rect 36311 8585 36320 8619
rect 36268 8576 36320 8585
rect 36636 8619 36688 8628
rect 36636 8585 36645 8619
rect 36645 8585 36679 8619
rect 36679 8585 36688 8619
rect 36636 8576 36688 8585
rect 26976 8440 27028 8492
rect 17960 8372 18012 8424
rect 21272 8372 21324 8424
rect 21548 8372 21600 8424
rect 24216 8372 24268 8424
rect 18420 8304 18472 8356
rect 19248 8304 19300 8356
rect 15752 8279 15804 8288
rect 15752 8245 15761 8279
rect 15761 8245 15795 8279
rect 15795 8245 15804 8279
rect 15752 8236 15804 8245
rect 17868 8236 17920 8288
rect 19064 8236 19116 8288
rect 20536 8304 20588 8356
rect 23756 8304 23808 8356
rect 21364 8236 21416 8288
rect 21548 8279 21600 8288
rect 21548 8245 21557 8279
rect 21557 8245 21591 8279
rect 21591 8245 21600 8279
rect 21548 8236 21600 8245
rect 22468 8279 22520 8288
rect 22468 8245 22477 8279
rect 22477 8245 22511 8279
rect 22511 8245 22520 8279
rect 22468 8236 22520 8245
rect 22928 8279 22980 8288
rect 22928 8245 22937 8279
rect 22937 8245 22971 8279
rect 22971 8245 22980 8279
rect 22928 8236 22980 8245
rect 23664 8236 23716 8288
rect 25872 8347 25924 8356
rect 25872 8313 25881 8347
rect 25881 8313 25915 8347
rect 25915 8313 25924 8347
rect 25872 8304 25924 8313
rect 24676 8236 24728 8288
rect 25136 8236 25188 8288
rect 26516 8236 26568 8288
rect 27528 8372 27580 8424
rect 27712 8372 27764 8424
rect 30288 8508 30340 8560
rect 30932 8508 30984 8560
rect 35624 8440 35676 8492
rect 32772 8415 32824 8424
rect 32772 8381 32781 8415
rect 32781 8381 32815 8415
rect 32815 8381 32824 8415
rect 32772 8372 32824 8381
rect 29644 8304 29696 8356
rect 30104 8347 30156 8356
rect 30104 8313 30113 8347
rect 30113 8313 30147 8347
rect 30147 8313 30156 8347
rect 30104 8304 30156 8313
rect 30196 8347 30248 8356
rect 30196 8313 30205 8347
rect 30205 8313 30239 8347
rect 30239 8313 30248 8347
rect 30196 8304 30248 8313
rect 32036 8304 32088 8356
rect 34060 8304 34112 8356
rect 28816 8236 28868 8288
rect 30472 8236 30524 8288
rect 32128 8279 32180 8288
rect 32128 8245 32137 8279
rect 32137 8245 32171 8279
rect 32171 8245 32180 8279
rect 32128 8236 32180 8245
rect 36268 8372 36320 8424
rect 34980 8347 35032 8356
rect 34980 8313 34989 8347
rect 34989 8313 35023 8347
rect 35023 8313 35032 8347
rect 34980 8304 35032 8313
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 2136 8075 2188 8084
rect 2136 8041 2145 8075
rect 2145 8041 2179 8075
rect 2179 8041 2188 8075
rect 2136 8032 2188 8041
rect 2688 8075 2740 8084
rect 2688 8041 2697 8075
rect 2697 8041 2731 8075
rect 2731 8041 2740 8075
rect 2688 8032 2740 8041
rect 4068 8032 4120 8084
rect 5816 8075 5868 8084
rect 5816 8041 5825 8075
rect 5825 8041 5859 8075
rect 5859 8041 5868 8075
rect 5816 8032 5868 8041
rect 6644 8032 6696 8084
rect 12164 8032 12216 8084
rect 3792 7964 3844 8016
rect 4252 8007 4304 8016
rect 4252 7973 4261 8007
rect 4261 7973 4295 8007
rect 4295 7973 4304 8007
rect 4804 8007 4856 8016
rect 4252 7964 4304 7973
rect 4804 7973 4813 8007
rect 4813 7973 4847 8007
rect 4847 7973 4856 8007
rect 4804 7964 4856 7973
rect 5080 7964 5132 8016
rect 6828 7964 6880 8016
rect 7196 8007 7248 8016
rect 7196 7973 7199 8007
rect 7199 7973 7233 8007
rect 7233 7973 7248 8007
rect 7196 7964 7248 7973
rect 11244 8007 11296 8016
rect 11244 7973 11253 8007
rect 11253 7973 11287 8007
rect 11287 7973 11296 8007
rect 11244 7964 11296 7973
rect 12624 8032 12676 8084
rect 12992 8032 13044 8084
rect 13176 8075 13228 8084
rect 13176 8041 13185 8075
rect 13185 8041 13219 8075
rect 13219 8041 13228 8075
rect 13176 8032 13228 8041
rect 17040 8032 17092 8084
rect 18512 8075 18564 8084
rect 18512 8041 18521 8075
rect 18521 8041 18555 8075
rect 18555 8041 18564 8075
rect 18512 8032 18564 8041
rect 19064 8032 19116 8084
rect 1768 7939 1820 7948
rect 1768 7905 1777 7939
rect 1777 7905 1811 7939
rect 1811 7905 1820 7939
rect 1768 7896 1820 7905
rect 5632 7939 5684 7948
rect 5632 7905 5641 7939
rect 5641 7905 5675 7939
rect 5675 7905 5684 7939
rect 5632 7896 5684 7905
rect 9036 7896 9088 7948
rect 10784 7939 10836 7948
rect 10784 7905 10793 7939
rect 10793 7905 10827 7939
rect 10827 7905 10836 7939
rect 10784 7896 10836 7905
rect 12072 7939 12124 7948
rect 6920 7828 6972 7880
rect 7380 7828 7432 7880
rect 10048 7828 10100 7880
rect 12072 7905 12081 7939
rect 12081 7905 12115 7939
rect 12115 7905 12124 7939
rect 12072 7896 12124 7905
rect 12164 7896 12216 7948
rect 13636 7939 13688 7948
rect 13636 7905 13645 7939
rect 13645 7905 13679 7939
rect 13679 7905 13688 7939
rect 13636 7896 13688 7905
rect 14648 8007 14700 8016
rect 14648 7973 14657 8007
rect 14657 7973 14691 8007
rect 14691 7973 14700 8007
rect 14648 7964 14700 7973
rect 15752 7964 15804 8016
rect 17592 8007 17644 8016
rect 17592 7973 17601 8007
rect 17601 7973 17635 8007
rect 17635 7973 17644 8007
rect 17592 7964 17644 7973
rect 17868 7964 17920 8016
rect 18236 7964 18288 8016
rect 22928 8032 22980 8084
rect 19248 8007 19300 8016
rect 19248 7973 19257 8007
rect 19257 7973 19291 8007
rect 19291 7973 19300 8007
rect 21640 8007 21692 8016
rect 19248 7964 19300 7973
rect 21640 7973 21649 8007
rect 21649 7973 21683 8007
rect 21683 7973 21692 8007
rect 21640 7964 21692 7973
rect 14096 7896 14148 7948
rect 14556 7828 14608 7880
rect 3516 7692 3568 7744
rect 5448 7735 5500 7744
rect 5448 7701 5457 7735
rect 5457 7701 5491 7735
rect 5491 7701 5500 7735
rect 5448 7692 5500 7701
rect 9772 7692 9824 7744
rect 13820 7692 13872 7744
rect 22652 7896 22704 7948
rect 23112 7896 23164 7948
rect 25872 8032 25924 8084
rect 30104 8032 30156 8084
rect 32404 8075 32456 8084
rect 32404 8041 32413 8075
rect 32413 8041 32447 8075
rect 32447 8041 32456 8075
rect 32404 8032 32456 8041
rect 24676 7964 24728 8016
rect 27344 7964 27396 8016
rect 28816 7964 28868 8016
rect 34060 7964 34112 8016
rect 35440 8007 35492 8016
rect 35440 7973 35449 8007
rect 35449 7973 35483 8007
rect 35483 7973 35492 8007
rect 35440 7964 35492 7973
rect 24124 7896 24176 7948
rect 27068 7896 27120 7948
rect 30196 7896 30248 7948
rect 32680 7896 32732 7948
rect 35164 7896 35216 7948
rect 18604 7828 18656 7880
rect 19524 7871 19576 7880
rect 19524 7837 19533 7871
rect 19533 7837 19567 7871
rect 19567 7837 19576 7871
rect 19524 7828 19576 7837
rect 21824 7871 21876 7880
rect 21824 7837 21833 7871
rect 21833 7837 21867 7871
rect 21867 7837 21876 7871
rect 21824 7828 21876 7837
rect 24400 7828 24452 7880
rect 25044 7828 25096 7880
rect 26700 7828 26752 7880
rect 29460 7828 29512 7880
rect 29644 7828 29696 7880
rect 30104 7871 30156 7880
rect 30104 7837 30113 7871
rect 30113 7837 30147 7871
rect 30147 7837 30156 7871
rect 30104 7828 30156 7837
rect 33508 7871 33560 7880
rect 33508 7837 33517 7871
rect 33517 7837 33551 7871
rect 33551 7837 33560 7871
rect 33508 7828 33560 7837
rect 35348 7871 35400 7880
rect 35348 7837 35357 7871
rect 35357 7837 35391 7871
rect 35391 7837 35400 7871
rect 35348 7828 35400 7837
rect 35624 7871 35676 7880
rect 35624 7837 35633 7871
rect 35633 7837 35667 7871
rect 35667 7837 35676 7871
rect 35624 7828 35676 7837
rect 17868 7760 17920 7812
rect 25688 7760 25740 7812
rect 30564 7760 30616 7812
rect 16856 7692 16908 7744
rect 20536 7692 20588 7744
rect 24216 7735 24268 7744
rect 24216 7701 24225 7735
rect 24225 7701 24259 7735
rect 24259 7701 24268 7735
rect 24216 7692 24268 7701
rect 27436 7735 27488 7744
rect 27436 7701 27445 7735
rect 27445 7701 27479 7735
rect 27479 7701 27488 7735
rect 27436 7692 27488 7701
rect 27712 7735 27764 7744
rect 27712 7701 27721 7735
rect 27721 7701 27755 7735
rect 27755 7701 27764 7735
rect 27712 7692 27764 7701
rect 33324 7760 33376 7812
rect 33416 7692 33468 7744
rect 34888 7735 34940 7744
rect 34888 7701 34897 7735
rect 34897 7701 34931 7735
rect 34931 7701 34940 7735
rect 34888 7692 34940 7701
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 3148 7531 3200 7540
rect 3148 7497 3157 7531
rect 3157 7497 3191 7531
rect 3191 7497 3200 7531
rect 3148 7488 3200 7497
rect 5356 7488 5408 7540
rect 9588 7531 9640 7540
rect 9588 7497 9597 7531
rect 9597 7497 9631 7531
rect 9631 7497 9640 7531
rect 9588 7488 9640 7497
rect 10232 7488 10284 7540
rect 12164 7488 12216 7540
rect 5908 7420 5960 7472
rect 10140 7420 10192 7472
rect 10784 7420 10836 7472
rect 14188 7488 14240 7540
rect 14556 7531 14608 7540
rect 14556 7497 14565 7531
rect 14565 7497 14599 7531
rect 14599 7497 14608 7531
rect 14556 7488 14608 7497
rect 15476 7488 15528 7540
rect 17868 7488 17920 7540
rect 19248 7488 19300 7540
rect 4068 7352 4120 7404
rect 5632 7352 5684 7404
rect 8300 7352 8352 7404
rect 9036 7352 9088 7404
rect 9864 7352 9916 7404
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 10416 7352 10468 7404
rect 13820 7352 13872 7404
rect 16120 7420 16172 7472
rect 20720 7488 20772 7540
rect 21640 7488 21692 7540
rect 23480 7531 23532 7540
rect 23480 7497 23489 7531
rect 23489 7497 23523 7531
rect 23523 7497 23532 7531
rect 23480 7488 23532 7497
rect 17040 7352 17092 7404
rect 19524 7352 19576 7404
rect 21548 7352 21600 7404
rect 3516 7284 3568 7336
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 8024 7284 8076 7336
rect 10048 7327 10100 7336
rect 10048 7293 10057 7327
rect 10057 7293 10091 7327
rect 10091 7293 10100 7327
rect 10048 7284 10100 7293
rect 12348 7284 12400 7336
rect 2136 7216 2188 7268
rect 3700 7216 3752 7268
rect 7196 7216 7248 7268
rect 8116 7216 8168 7268
rect 5080 7191 5132 7200
rect 5080 7157 5089 7191
rect 5089 7157 5123 7191
rect 5123 7157 5132 7191
rect 5080 7148 5132 7157
rect 6920 7148 6972 7200
rect 7104 7148 7156 7200
rect 10048 7148 10100 7200
rect 10140 7148 10192 7200
rect 10416 7216 10468 7268
rect 12440 7216 12492 7268
rect 13636 7216 13688 7268
rect 14004 7216 14056 7268
rect 15292 7284 15344 7336
rect 15752 7284 15804 7336
rect 16212 7216 16264 7268
rect 20628 7327 20680 7336
rect 16672 7216 16724 7268
rect 10968 7191 11020 7200
rect 10968 7157 10977 7191
rect 10977 7157 11011 7191
rect 11011 7157 11020 7191
rect 10968 7148 11020 7157
rect 12164 7191 12216 7200
rect 12164 7157 12173 7191
rect 12173 7157 12207 7191
rect 12207 7157 12216 7191
rect 12164 7148 12216 7157
rect 12900 7148 12952 7200
rect 20628 7293 20637 7327
rect 20637 7293 20671 7327
rect 20671 7293 20680 7327
rect 20628 7284 20680 7293
rect 22836 7284 22888 7336
rect 28908 7488 28960 7540
rect 32680 7531 32732 7540
rect 32680 7497 32689 7531
rect 32689 7497 32723 7531
rect 32723 7497 32732 7531
rect 32680 7488 32732 7497
rect 34060 7488 34112 7540
rect 35440 7488 35492 7540
rect 36636 7531 36688 7540
rect 36636 7497 36645 7531
rect 36645 7497 36679 7531
rect 36679 7497 36688 7531
rect 36636 7488 36688 7497
rect 26976 7420 27028 7472
rect 27528 7420 27580 7472
rect 34888 7420 34940 7472
rect 24216 7395 24268 7404
rect 24216 7361 24225 7395
rect 24225 7361 24259 7395
rect 24259 7361 24268 7395
rect 24216 7352 24268 7361
rect 26148 7352 26200 7404
rect 27712 7395 27764 7404
rect 27712 7361 27721 7395
rect 27721 7361 27755 7395
rect 27755 7361 27764 7395
rect 27712 7352 27764 7361
rect 27988 7352 28040 7404
rect 28816 7352 28868 7404
rect 30104 7395 30156 7404
rect 24124 7327 24176 7336
rect 24124 7293 24133 7327
rect 24133 7293 24167 7327
rect 24167 7293 24176 7327
rect 24124 7284 24176 7293
rect 18604 7148 18656 7200
rect 19432 7216 19484 7268
rect 21364 7259 21416 7268
rect 21364 7225 21373 7259
rect 21373 7225 21407 7259
rect 21407 7225 21416 7259
rect 21364 7216 21416 7225
rect 27344 7216 27396 7268
rect 22008 7148 22060 7200
rect 22652 7191 22704 7200
rect 22652 7157 22661 7191
rect 22661 7157 22695 7191
rect 22695 7157 22704 7191
rect 22652 7148 22704 7157
rect 23020 7191 23072 7200
rect 23020 7157 23029 7191
rect 23029 7157 23063 7191
rect 23063 7157 23072 7191
rect 23020 7148 23072 7157
rect 24676 7191 24728 7200
rect 24676 7157 24685 7191
rect 24685 7157 24719 7191
rect 24719 7157 24728 7191
rect 24676 7148 24728 7157
rect 25044 7191 25096 7200
rect 25044 7157 25053 7191
rect 25053 7157 25087 7191
rect 25087 7157 25096 7191
rect 25044 7148 25096 7157
rect 30104 7361 30113 7395
rect 30113 7361 30147 7395
rect 30147 7361 30156 7395
rect 30104 7352 30156 7361
rect 31760 7284 31812 7336
rect 32036 7216 32088 7268
rect 33416 7352 33468 7404
rect 35348 7395 35400 7404
rect 33324 7259 33376 7268
rect 29460 7191 29512 7200
rect 29460 7157 29469 7191
rect 29469 7157 29503 7191
rect 29503 7157 29512 7191
rect 29460 7148 29512 7157
rect 33324 7225 33333 7259
rect 33333 7225 33367 7259
rect 33367 7225 33376 7259
rect 33324 7216 33376 7225
rect 33416 7259 33468 7268
rect 33416 7225 33425 7259
rect 33425 7225 33459 7259
rect 33459 7225 33468 7259
rect 33416 7216 33468 7225
rect 35348 7361 35357 7395
rect 35357 7361 35391 7395
rect 35391 7361 35400 7395
rect 35348 7352 35400 7361
rect 34060 7148 34112 7200
rect 35164 7216 35216 7268
rect 34980 7148 35032 7200
rect 36360 7148 36412 7200
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 1768 6987 1820 6996
rect 1768 6953 1777 6987
rect 1777 6953 1811 6987
rect 1811 6953 1820 6987
rect 1768 6944 1820 6953
rect 2872 6944 2924 6996
rect 10416 6944 10468 6996
rect 14004 6987 14056 6996
rect 14004 6953 14013 6987
rect 14013 6953 14047 6987
rect 14047 6953 14056 6987
rect 14004 6944 14056 6953
rect 14188 6944 14240 6996
rect 17592 6944 17644 6996
rect 18512 6987 18564 6996
rect 18512 6953 18521 6987
rect 18521 6953 18555 6987
rect 18555 6953 18564 6987
rect 18512 6944 18564 6953
rect 19432 6944 19484 6996
rect 2136 6876 2188 6928
rect 4160 6876 4212 6928
rect 5080 6876 5132 6928
rect 7196 6876 7248 6928
rect 9772 6876 9824 6928
rect 12164 6876 12216 6928
rect 14096 6876 14148 6928
rect 16304 6876 16356 6928
rect 16672 6876 16724 6928
rect 19340 6876 19392 6928
rect 21548 6944 21600 6996
rect 21640 6944 21692 6996
rect 6736 6808 6788 6860
rect 8576 6851 8628 6860
rect 8576 6817 8585 6851
rect 8585 6817 8619 6851
rect 8619 6817 8628 6851
rect 8576 6808 8628 6817
rect 10140 6808 10192 6860
rect 14740 6808 14792 6860
rect 17592 6851 17644 6860
rect 17592 6817 17601 6851
rect 17601 6817 17635 6851
rect 17635 6817 17644 6851
rect 17592 6808 17644 6817
rect 17776 6851 17828 6860
rect 17776 6817 17785 6851
rect 17785 6817 17819 6851
rect 17819 6817 17828 6851
rect 17776 6808 17828 6817
rect 18696 6808 18748 6860
rect 21272 6876 21324 6928
rect 21824 6808 21876 6860
rect 22468 6851 22520 6860
rect 22468 6817 22512 6851
rect 22512 6817 22520 6851
rect 22468 6808 22520 6817
rect 23112 6808 23164 6860
rect 25044 6876 25096 6928
rect 26148 6944 26200 6996
rect 28264 6944 28316 6996
rect 30288 6987 30340 6996
rect 30288 6953 30297 6987
rect 30297 6953 30331 6987
rect 30331 6953 30340 6987
rect 30288 6944 30340 6953
rect 33324 6944 33376 6996
rect 27436 6876 27488 6928
rect 28816 6919 28868 6928
rect 28816 6885 28825 6919
rect 28825 6885 28859 6919
rect 28859 6885 28868 6919
rect 28816 6876 28868 6885
rect 3240 6740 3292 6792
rect 3884 6740 3936 6792
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 3056 6672 3108 6724
rect 5448 6740 5500 6792
rect 9680 6783 9732 6792
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 9680 6740 9732 6749
rect 11980 6783 12032 6792
rect 11980 6749 11989 6783
rect 11989 6749 12023 6783
rect 12023 6749 12032 6783
rect 11980 6740 12032 6749
rect 14832 6740 14884 6792
rect 16028 6783 16080 6792
rect 16028 6749 16037 6783
rect 16037 6749 16071 6783
rect 16071 6749 16080 6783
rect 16028 6740 16080 6749
rect 16120 6740 16172 6792
rect 18880 6740 18932 6792
rect 24400 6808 24452 6860
rect 25320 6851 25372 6860
rect 25320 6817 25329 6851
rect 25329 6817 25363 6851
rect 25363 6817 25372 6851
rect 25320 6808 25372 6817
rect 30472 6851 30524 6860
rect 30472 6817 30481 6851
rect 30481 6817 30515 6851
rect 30515 6817 30524 6851
rect 30472 6808 30524 6817
rect 32036 6876 32088 6928
rect 34612 6919 34664 6928
rect 34612 6885 34621 6919
rect 34621 6885 34655 6919
rect 34655 6885 34664 6919
rect 34612 6876 34664 6885
rect 35348 6944 35400 6996
rect 36176 6919 36228 6928
rect 36176 6885 36185 6919
rect 36185 6885 36219 6919
rect 36219 6885 36228 6919
rect 36176 6876 36228 6885
rect 31116 6808 31168 6860
rect 26332 6740 26384 6792
rect 27528 6783 27580 6792
rect 27528 6749 27537 6783
rect 27537 6749 27571 6783
rect 27571 6749 27580 6783
rect 27528 6740 27580 6749
rect 28724 6783 28776 6792
rect 28724 6749 28733 6783
rect 28733 6749 28767 6783
rect 28767 6749 28776 6783
rect 28724 6740 28776 6749
rect 29644 6740 29696 6792
rect 33876 6740 33928 6792
rect 34152 6740 34204 6792
rect 36084 6783 36136 6792
rect 36084 6749 36093 6783
rect 36093 6749 36127 6783
rect 36127 6749 36136 6783
rect 36084 6740 36136 6749
rect 36360 6783 36412 6792
rect 36360 6749 36369 6783
rect 36369 6749 36403 6783
rect 36403 6749 36412 6783
rect 36360 6740 36412 6749
rect 24952 6672 25004 6724
rect 26240 6672 26292 6724
rect 2964 6604 3016 6656
rect 7012 6604 7064 6656
rect 8024 6604 8076 6656
rect 8484 6604 8536 6656
rect 9036 6647 9088 6656
rect 9036 6613 9045 6647
rect 9045 6613 9079 6647
rect 9079 6613 9088 6647
rect 9036 6604 9088 6613
rect 10876 6604 10928 6656
rect 16948 6647 17000 6656
rect 16948 6613 16957 6647
rect 16957 6613 16991 6647
rect 16991 6613 17000 6647
rect 16948 6604 17000 6613
rect 18972 6604 19024 6656
rect 25412 6604 25464 6656
rect 26700 6647 26752 6656
rect 26700 6613 26709 6647
rect 26709 6613 26743 6647
rect 26743 6613 26752 6647
rect 26700 6604 26752 6613
rect 33048 6647 33100 6656
rect 33048 6613 33057 6647
rect 33057 6613 33091 6647
rect 33091 6613 33100 6647
rect 33048 6604 33100 6613
rect 33324 6604 33376 6656
rect 33508 6647 33560 6656
rect 33508 6613 33517 6647
rect 33517 6613 33551 6647
rect 33551 6613 33560 6647
rect 33508 6604 33560 6613
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 2136 6400 2188 6452
rect 4160 6443 4212 6452
rect 4160 6409 4169 6443
rect 4169 6409 4203 6443
rect 4203 6409 4212 6443
rect 4160 6400 4212 6409
rect 4436 6400 4488 6452
rect 7196 6400 7248 6452
rect 8392 6400 8444 6452
rect 9680 6400 9732 6452
rect 9956 6400 10008 6452
rect 14004 6400 14056 6452
rect 15292 6443 15344 6452
rect 15292 6409 15301 6443
rect 15301 6409 15335 6443
rect 15335 6409 15344 6443
rect 15292 6400 15344 6409
rect 16304 6443 16356 6452
rect 16304 6409 16313 6443
rect 16313 6409 16347 6443
rect 16347 6409 16356 6443
rect 16304 6400 16356 6409
rect 17776 6400 17828 6452
rect 21272 6443 21324 6452
rect 21272 6409 21281 6443
rect 21281 6409 21315 6443
rect 21315 6409 21324 6443
rect 21272 6400 21324 6409
rect 23112 6443 23164 6452
rect 23112 6409 23121 6443
rect 23121 6409 23155 6443
rect 23155 6409 23164 6443
rect 23112 6400 23164 6409
rect 24952 6443 25004 6452
rect 24952 6409 24961 6443
rect 24961 6409 24995 6443
rect 24995 6409 25004 6443
rect 24952 6400 25004 6409
rect 25320 6443 25372 6452
rect 25320 6409 25329 6443
rect 25329 6409 25363 6443
rect 25363 6409 25372 6443
rect 25320 6400 25372 6409
rect 27436 6400 27488 6452
rect 9772 6332 9824 6384
rect 12164 6332 12216 6384
rect 12256 6332 12308 6384
rect 13452 6332 13504 6384
rect 16028 6332 16080 6384
rect 17592 6332 17644 6384
rect 18236 6375 18288 6384
rect 18236 6341 18245 6375
rect 18245 6341 18279 6375
rect 18279 6341 18288 6375
rect 18236 6332 18288 6341
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 2872 6264 2924 6316
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 3148 6128 3200 6180
rect 2964 6060 3016 6112
rect 4436 6264 4488 6316
rect 7012 6264 7064 6316
rect 9036 6264 9088 6316
rect 14740 6307 14792 6316
rect 14740 6273 14749 6307
rect 14749 6273 14783 6307
rect 14783 6273 14792 6307
rect 14740 6264 14792 6273
rect 16856 6264 16908 6316
rect 17132 6264 17184 6316
rect 18512 6307 18564 6316
rect 18512 6273 18521 6307
rect 18521 6273 18555 6307
rect 18555 6273 18564 6307
rect 18512 6264 18564 6273
rect 18696 6264 18748 6316
rect 23756 6332 23808 6384
rect 8668 6239 8720 6248
rect 8668 6205 8677 6239
rect 8677 6205 8711 6239
rect 8711 6205 8720 6239
rect 8668 6196 8720 6205
rect 4344 6171 4396 6180
rect 4344 6137 4353 6171
rect 4353 6137 4387 6171
rect 4387 6137 4396 6171
rect 4344 6128 4396 6137
rect 4436 6171 4488 6180
rect 4436 6137 4445 6171
rect 4445 6137 4479 6171
rect 4479 6137 4488 6171
rect 4436 6128 4488 6137
rect 4804 6128 4856 6180
rect 7012 6171 7064 6180
rect 7012 6137 7021 6171
rect 7021 6137 7055 6171
rect 7055 6137 7064 6171
rect 7012 6128 7064 6137
rect 8392 6128 8444 6180
rect 12992 6196 13044 6248
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 15384 6239 15436 6248
rect 10784 6171 10836 6180
rect 10784 6137 10793 6171
rect 10793 6137 10827 6171
rect 10827 6137 10836 6171
rect 10784 6128 10836 6137
rect 10876 6171 10928 6180
rect 10876 6137 10885 6171
rect 10885 6137 10919 6171
rect 10919 6137 10928 6171
rect 10876 6128 10928 6137
rect 13084 6128 13136 6180
rect 15384 6205 15393 6239
rect 15393 6205 15427 6239
rect 15427 6205 15436 6239
rect 15384 6196 15436 6205
rect 17684 6196 17736 6248
rect 20168 6196 20220 6248
rect 23480 6264 23532 6316
rect 28080 6332 28132 6384
rect 28816 6400 28868 6452
rect 28908 6400 28960 6452
rect 30472 6375 30524 6384
rect 30472 6341 30481 6375
rect 30481 6341 30515 6375
rect 30515 6341 30524 6375
rect 30472 6332 30524 6341
rect 27988 6307 28040 6316
rect 27988 6273 27997 6307
rect 27997 6273 28031 6307
rect 28031 6273 28040 6307
rect 27988 6264 28040 6273
rect 29184 6264 29236 6316
rect 29644 6307 29696 6316
rect 29644 6273 29653 6307
rect 29653 6273 29687 6307
rect 29687 6273 29696 6307
rect 29644 6264 29696 6273
rect 22100 6196 22152 6248
rect 23664 6239 23716 6248
rect 23664 6205 23673 6239
rect 23673 6205 23707 6239
rect 23707 6205 23716 6239
rect 23664 6196 23716 6205
rect 25872 6239 25924 6248
rect 25872 6205 25881 6239
rect 25881 6205 25915 6239
rect 25915 6205 25924 6239
rect 25872 6196 25924 6205
rect 32956 6400 33008 6452
rect 33876 6443 33928 6452
rect 33876 6409 33885 6443
rect 33885 6409 33919 6443
rect 33919 6409 33928 6443
rect 33876 6400 33928 6409
rect 36084 6400 36136 6452
rect 36452 6400 36504 6452
rect 32036 6332 32088 6384
rect 33048 6332 33100 6384
rect 34612 6332 34664 6384
rect 36176 6332 36228 6384
rect 32128 6264 32180 6316
rect 35164 6264 35216 6316
rect 35348 6307 35400 6316
rect 35348 6273 35357 6307
rect 35357 6273 35391 6307
rect 35391 6273 35400 6307
rect 35348 6264 35400 6273
rect 31208 6196 31260 6248
rect 32680 6239 32732 6248
rect 32680 6205 32689 6239
rect 32689 6205 32723 6239
rect 32723 6205 32732 6239
rect 32680 6196 32732 6205
rect 34612 6239 34664 6248
rect 34612 6205 34621 6239
rect 34621 6205 34655 6239
rect 34655 6205 34664 6239
rect 34612 6196 34664 6205
rect 8484 6103 8536 6112
rect 8484 6069 8493 6103
rect 8493 6069 8527 6103
rect 8527 6069 8536 6103
rect 8484 6060 8536 6069
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 18604 6171 18656 6180
rect 15292 6060 15344 6112
rect 18604 6137 18613 6171
rect 18613 6137 18647 6171
rect 18647 6137 18656 6171
rect 18604 6128 18656 6137
rect 19340 6128 19392 6180
rect 21364 6128 21416 6180
rect 24676 6128 24728 6180
rect 16212 6060 16264 6112
rect 20628 6060 20680 6112
rect 22284 6103 22336 6112
rect 22284 6069 22293 6103
rect 22293 6069 22327 6103
rect 22327 6069 22336 6103
rect 22284 6060 22336 6069
rect 23572 6060 23624 6112
rect 24584 6103 24636 6112
rect 24584 6069 24593 6103
rect 24593 6069 24627 6103
rect 24627 6069 24636 6103
rect 24584 6060 24636 6069
rect 28816 6128 28868 6180
rect 29368 6171 29420 6180
rect 29368 6137 29377 6171
rect 29377 6137 29411 6171
rect 29411 6137 29420 6171
rect 29368 6128 29420 6137
rect 34980 6171 35032 6180
rect 29000 6103 29052 6112
rect 29000 6069 29009 6103
rect 29009 6069 29043 6103
rect 29043 6069 29052 6103
rect 34980 6137 34989 6171
rect 34989 6137 35023 6171
rect 35023 6137 35032 6171
rect 34980 6128 35032 6137
rect 29000 6060 29052 6069
rect 34612 6060 34664 6112
rect 36912 6103 36964 6112
rect 36912 6069 36921 6103
rect 36921 6069 36955 6103
rect 36955 6069 36964 6103
rect 36912 6060 36964 6069
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 2136 5856 2188 5908
rect 3148 5856 3200 5908
rect 3240 5899 3292 5908
rect 3240 5865 3249 5899
rect 3249 5865 3283 5899
rect 3283 5865 3292 5899
rect 3240 5856 3292 5865
rect 3424 5856 3476 5908
rect 4344 5856 4396 5908
rect 6736 5899 6788 5908
rect 6736 5865 6745 5899
rect 6745 5865 6779 5899
rect 6779 5865 6788 5899
rect 6736 5856 6788 5865
rect 6920 5856 6972 5908
rect 8668 5856 8720 5908
rect 12072 5856 12124 5908
rect 13084 5899 13136 5908
rect 2044 5831 2096 5840
rect 2044 5797 2053 5831
rect 2053 5797 2087 5831
rect 2087 5797 2096 5831
rect 2044 5788 2096 5797
rect 2688 5788 2740 5840
rect 5816 5831 5868 5840
rect 5816 5797 5825 5831
rect 5825 5797 5859 5831
rect 5859 5797 5868 5831
rect 5816 5788 5868 5797
rect 3792 5720 3844 5772
rect 4804 5763 4856 5772
rect 4804 5729 4813 5763
rect 4813 5729 4847 5763
rect 4847 5729 4856 5763
rect 7104 5763 7156 5772
rect 4804 5720 4856 5729
rect 7104 5729 7113 5763
rect 7113 5729 7147 5763
rect 7147 5729 7156 5763
rect 7104 5720 7156 5729
rect 3240 5652 3292 5704
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 5356 5584 5408 5636
rect 6644 5652 6696 5704
rect 8392 5720 8444 5772
rect 9772 5788 9824 5840
rect 13084 5865 13093 5899
rect 13093 5865 13127 5899
rect 13127 5865 13136 5899
rect 13084 5856 13136 5865
rect 13912 5856 13964 5908
rect 18604 5856 18656 5908
rect 18696 5856 18748 5908
rect 21456 5856 21508 5908
rect 22468 5899 22520 5908
rect 12900 5788 12952 5840
rect 13452 5788 13504 5840
rect 14556 5788 14608 5840
rect 16948 5831 17000 5840
rect 16948 5797 16957 5831
rect 16957 5797 16991 5831
rect 16991 5797 17000 5831
rect 16948 5788 17000 5797
rect 10416 5720 10468 5772
rect 9680 5695 9732 5704
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 9680 5652 9732 5661
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 14832 5652 14884 5704
rect 10784 5584 10836 5636
rect 13820 5584 13872 5636
rect 16120 5652 16172 5704
rect 19340 5788 19392 5840
rect 20628 5788 20680 5840
rect 22468 5865 22477 5899
rect 22477 5865 22511 5899
rect 22511 5865 22520 5899
rect 22468 5856 22520 5865
rect 23572 5899 23624 5908
rect 23572 5865 23581 5899
rect 23581 5865 23615 5899
rect 23615 5865 23624 5899
rect 23572 5856 23624 5865
rect 23664 5856 23716 5908
rect 26332 5899 26384 5908
rect 26332 5865 26341 5899
rect 26341 5865 26375 5899
rect 26375 5865 26384 5899
rect 26332 5856 26384 5865
rect 29184 5856 29236 5908
rect 31116 5899 31168 5908
rect 24584 5788 24636 5840
rect 27528 5788 27580 5840
rect 27988 5788 28040 5840
rect 28448 5788 28500 5840
rect 18328 5720 18380 5772
rect 24676 5720 24728 5772
rect 25136 5763 25188 5772
rect 25136 5729 25145 5763
rect 25145 5729 25179 5763
rect 25179 5729 25188 5763
rect 25136 5720 25188 5729
rect 30104 5763 30156 5772
rect 30104 5729 30113 5763
rect 30113 5729 30147 5763
rect 30147 5729 30156 5763
rect 30104 5720 30156 5729
rect 30196 5720 30248 5772
rect 31116 5865 31125 5899
rect 31125 5865 31159 5899
rect 31159 5865 31168 5899
rect 31116 5856 31168 5865
rect 32680 5899 32732 5908
rect 32680 5865 32689 5899
rect 32689 5865 32723 5899
rect 32723 5865 32732 5899
rect 32680 5856 32732 5865
rect 34152 5856 34204 5908
rect 34980 5856 35032 5908
rect 36452 5899 36504 5908
rect 36452 5865 36461 5899
rect 36461 5865 36495 5899
rect 36495 5865 36504 5899
rect 36452 5856 36504 5865
rect 33324 5788 33376 5840
rect 34612 5831 34664 5840
rect 34612 5797 34621 5831
rect 34621 5797 34655 5831
rect 34655 5797 34664 5831
rect 34612 5788 34664 5797
rect 36360 5788 36412 5840
rect 32128 5720 32180 5772
rect 33600 5720 33652 5772
rect 36268 5720 36320 5772
rect 20812 5652 20864 5704
rect 22284 5652 22336 5704
rect 25504 5695 25556 5704
rect 25504 5661 25513 5695
rect 25513 5661 25547 5695
rect 25547 5661 25556 5695
rect 25504 5652 25556 5661
rect 27068 5695 27120 5704
rect 27068 5661 27077 5695
rect 27077 5661 27111 5695
rect 27111 5661 27120 5695
rect 27068 5652 27120 5661
rect 28632 5695 28684 5704
rect 28632 5661 28641 5695
rect 28641 5661 28675 5695
rect 28675 5661 28684 5695
rect 28632 5652 28684 5661
rect 29368 5652 29420 5704
rect 34152 5652 34204 5704
rect 19616 5584 19668 5636
rect 23112 5584 23164 5636
rect 29184 5627 29236 5636
rect 29184 5593 29193 5627
rect 29193 5593 29227 5627
rect 29227 5593 29236 5627
rect 29184 5584 29236 5593
rect 8576 5516 8628 5568
rect 9036 5516 9088 5568
rect 11980 5559 12032 5568
rect 11980 5525 11989 5559
rect 11989 5525 12023 5559
rect 12023 5525 12032 5559
rect 11980 5516 12032 5525
rect 12348 5516 12400 5568
rect 14740 5559 14792 5568
rect 14740 5525 14749 5559
rect 14749 5525 14783 5559
rect 14783 5525 14792 5559
rect 14740 5516 14792 5525
rect 15384 5516 15436 5568
rect 16304 5516 16356 5568
rect 16672 5516 16724 5568
rect 17776 5516 17828 5568
rect 20168 5559 20220 5568
rect 20168 5525 20177 5559
rect 20177 5525 20211 5559
rect 20211 5525 20220 5559
rect 20168 5516 20220 5525
rect 20720 5559 20772 5568
rect 20720 5525 20729 5559
rect 20729 5525 20763 5559
rect 20763 5525 20772 5559
rect 20720 5516 20772 5525
rect 22100 5559 22152 5568
rect 22100 5525 22109 5559
rect 22109 5525 22143 5559
rect 22143 5525 22152 5559
rect 22100 5516 22152 5525
rect 24124 5559 24176 5568
rect 24124 5525 24133 5559
rect 24133 5525 24167 5559
rect 24167 5525 24176 5559
rect 24124 5516 24176 5525
rect 25872 5559 25924 5568
rect 25872 5525 25881 5559
rect 25881 5525 25915 5559
rect 25915 5525 25924 5559
rect 25872 5516 25924 5525
rect 28080 5559 28132 5568
rect 28080 5525 28089 5559
rect 28089 5525 28123 5559
rect 28123 5525 28132 5559
rect 28080 5516 28132 5525
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 2044 5312 2096 5364
rect 3700 5312 3752 5364
rect 5816 5312 5868 5364
rect 8668 5312 8720 5364
rect 9772 5312 9824 5364
rect 12072 5355 12124 5364
rect 12072 5321 12081 5355
rect 12081 5321 12115 5355
rect 12115 5321 12124 5355
rect 12072 5312 12124 5321
rect 6644 5287 6696 5296
rect 6644 5253 6653 5287
rect 6653 5253 6687 5287
rect 6687 5253 6696 5287
rect 6644 5244 6696 5253
rect 7380 5244 7432 5296
rect 11428 5244 11480 5296
rect 14556 5355 14608 5364
rect 14556 5321 14565 5355
rect 14565 5321 14599 5355
rect 14599 5321 14608 5355
rect 14556 5312 14608 5321
rect 17776 5312 17828 5364
rect 19340 5355 19392 5364
rect 19340 5321 19349 5355
rect 19349 5321 19383 5355
rect 19383 5321 19392 5355
rect 20536 5355 20588 5364
rect 19340 5312 19392 5321
rect 20536 5321 20545 5355
rect 20545 5321 20579 5355
rect 20579 5321 20588 5355
rect 20536 5312 20588 5321
rect 20812 5312 20864 5364
rect 22284 5312 22336 5364
rect 24124 5312 24176 5364
rect 27252 5312 27304 5364
rect 27528 5312 27580 5364
rect 28448 5312 28500 5364
rect 28724 5312 28776 5364
rect 29828 5355 29880 5364
rect 29828 5321 29837 5355
rect 29837 5321 29871 5355
rect 29871 5321 29880 5355
rect 29828 5312 29880 5321
rect 30104 5355 30156 5364
rect 30104 5321 30113 5355
rect 30113 5321 30147 5355
rect 30147 5321 30156 5355
rect 30104 5312 30156 5321
rect 30748 5355 30800 5364
rect 30748 5321 30757 5355
rect 30757 5321 30791 5355
rect 30791 5321 30800 5355
rect 30748 5312 30800 5321
rect 33600 5312 33652 5364
rect 34152 5355 34204 5364
rect 34152 5321 34161 5355
rect 34161 5321 34195 5355
rect 34195 5321 34204 5355
rect 34152 5312 34204 5321
rect 34612 5312 34664 5364
rect 34980 5312 35032 5364
rect 35992 5312 36044 5364
rect 36268 5312 36320 5364
rect 25044 5287 25096 5296
rect 25044 5253 25053 5287
rect 25053 5253 25087 5287
rect 25087 5253 25096 5287
rect 25044 5244 25096 5253
rect 26240 5287 26292 5296
rect 26240 5253 26249 5287
rect 26249 5253 26283 5287
rect 26283 5253 26292 5287
rect 26240 5244 26292 5253
rect 27068 5244 27120 5296
rect 14740 5219 14792 5228
rect 1768 5108 1820 5160
rect 3700 5151 3752 5160
rect 3700 5117 3709 5151
rect 3709 5117 3743 5151
rect 3743 5117 3752 5151
rect 3700 5108 3752 5117
rect 3240 5015 3292 5024
rect 3240 4981 3249 5015
rect 3249 4981 3283 5015
rect 3283 4981 3292 5015
rect 3240 4972 3292 4981
rect 6368 5108 6420 5160
rect 8852 5108 8904 5160
rect 8116 5083 8168 5092
rect 8116 5049 8125 5083
rect 8125 5049 8159 5083
rect 8159 5049 8168 5083
rect 8116 5040 8168 5049
rect 9772 5040 9824 5092
rect 13820 5151 13872 5160
rect 13820 5117 13829 5151
rect 13829 5117 13863 5151
rect 13863 5117 13872 5151
rect 13820 5108 13872 5117
rect 13176 5083 13228 5092
rect 13176 5049 13185 5083
rect 13185 5049 13219 5083
rect 13219 5049 13228 5083
rect 13176 5040 13228 5049
rect 13268 5083 13320 5092
rect 13268 5049 13277 5083
rect 13277 5049 13311 5083
rect 13311 5049 13320 5083
rect 14740 5185 14749 5219
rect 14749 5185 14783 5219
rect 14783 5185 14792 5219
rect 14740 5176 14792 5185
rect 14832 5176 14884 5228
rect 16948 5176 17000 5228
rect 18788 5176 18840 5228
rect 20168 5219 20220 5228
rect 16212 5151 16264 5160
rect 16212 5117 16221 5151
rect 16221 5117 16255 5151
rect 16255 5117 16264 5151
rect 16212 5108 16264 5117
rect 14832 5083 14884 5092
rect 13268 5040 13320 5049
rect 14832 5049 14841 5083
rect 14841 5049 14875 5083
rect 14875 5049 14884 5083
rect 14832 5040 14884 5049
rect 6460 4972 6512 5024
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 12900 5015 12952 5024
rect 12900 4981 12909 5015
rect 12909 4981 12943 5015
rect 12943 4981 12952 5015
rect 12900 4972 12952 4981
rect 13820 4972 13872 5024
rect 18144 5108 18196 5160
rect 19248 5108 19300 5160
rect 19616 5151 19668 5160
rect 19616 5117 19625 5151
rect 19625 5117 19659 5151
rect 19659 5117 19668 5151
rect 19616 5108 19668 5117
rect 20168 5185 20177 5219
rect 20177 5185 20211 5219
rect 20211 5185 20220 5219
rect 20168 5176 20220 5185
rect 20536 5108 20588 5160
rect 20720 5108 20772 5160
rect 21456 5108 21508 5160
rect 23756 5151 23808 5160
rect 23756 5117 23765 5151
rect 23765 5117 23799 5151
rect 23799 5117 23808 5151
rect 23756 5108 23808 5117
rect 25872 5219 25924 5228
rect 25872 5185 25881 5219
rect 25881 5185 25915 5219
rect 25915 5185 25924 5219
rect 25872 5176 25924 5185
rect 27988 5176 28040 5228
rect 28632 5176 28684 5228
rect 31760 5219 31812 5228
rect 31760 5185 31769 5219
rect 31769 5185 31803 5219
rect 31803 5185 31812 5219
rect 31760 5176 31812 5185
rect 18512 5040 18564 5092
rect 19708 5040 19760 5092
rect 22100 5040 22152 5092
rect 24032 5040 24084 5092
rect 25320 5040 25372 5092
rect 29828 5108 29880 5160
rect 30748 5108 30800 5160
rect 15752 5015 15804 5024
rect 15752 4981 15761 5015
rect 15761 4981 15795 5015
rect 15795 4981 15804 5015
rect 15752 4972 15804 4981
rect 16304 5015 16356 5024
rect 16304 4981 16313 5015
rect 16313 4981 16347 5015
rect 16347 4981 16356 5015
rect 16304 4972 16356 4981
rect 23572 4972 23624 5024
rect 23664 4972 23716 5024
rect 24676 5015 24728 5024
rect 24676 4981 24685 5015
rect 24685 4981 24719 5015
rect 24719 4981 24728 5015
rect 24676 4972 24728 4981
rect 27252 5083 27304 5092
rect 27252 5049 27261 5083
rect 27261 5049 27295 5083
rect 27295 5049 27304 5083
rect 27252 5040 27304 5049
rect 29000 5040 29052 5092
rect 28172 5015 28224 5024
rect 28172 4981 28181 5015
rect 28181 4981 28215 5015
rect 28215 4981 28224 5015
rect 28172 4972 28224 4981
rect 32128 5015 32180 5024
rect 32128 4981 32137 5015
rect 32137 4981 32171 5015
rect 32171 4981 32180 5015
rect 32128 4972 32180 4981
rect 35440 5015 35492 5024
rect 35440 4981 35449 5015
rect 35449 4981 35483 5015
rect 35483 4981 35492 5015
rect 35440 4972 35492 4981
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 2044 4768 2096 4820
rect 3700 4811 3752 4820
rect 3700 4777 3709 4811
rect 3709 4777 3743 4811
rect 3743 4777 3752 4811
rect 3700 4768 3752 4777
rect 5448 4768 5500 4820
rect 5724 4768 5776 4820
rect 6828 4768 6880 4820
rect 9680 4768 9732 4820
rect 11888 4768 11940 4820
rect 12164 4768 12216 4820
rect 12348 4811 12400 4820
rect 12348 4777 12357 4811
rect 12357 4777 12391 4811
rect 12391 4777 12400 4811
rect 12348 4768 12400 4777
rect 13176 4811 13228 4820
rect 13176 4777 13185 4811
rect 13185 4777 13219 4811
rect 13219 4777 13228 4811
rect 13176 4768 13228 4777
rect 13452 4811 13504 4820
rect 13452 4777 13461 4811
rect 13461 4777 13495 4811
rect 13495 4777 13504 4811
rect 13452 4768 13504 4777
rect 14832 4768 14884 4820
rect 18144 4768 18196 4820
rect 18328 4768 18380 4820
rect 20628 4811 20680 4820
rect 20628 4777 20637 4811
rect 20637 4777 20671 4811
rect 20671 4777 20680 4811
rect 20628 4768 20680 4777
rect 20812 4768 20864 4820
rect 23756 4811 23808 4820
rect 23756 4777 23765 4811
rect 23765 4777 23799 4811
rect 23799 4777 23808 4811
rect 23756 4768 23808 4777
rect 27528 4811 27580 4820
rect 27528 4777 27537 4811
rect 27537 4777 27571 4811
rect 27571 4777 27580 4811
rect 27528 4768 27580 4777
rect 28080 4768 28132 4820
rect 30196 4811 30248 4820
rect 30196 4777 30205 4811
rect 30205 4777 30239 4811
rect 30239 4777 30248 4811
rect 30196 4768 30248 4777
rect 2872 4700 2924 4752
rect 1676 4632 1728 4684
rect 4528 4700 4580 4752
rect 6000 4700 6052 4752
rect 6368 4743 6420 4752
rect 6368 4709 6377 4743
rect 6377 4709 6411 4743
rect 6411 4709 6420 4743
rect 6368 4700 6420 4709
rect 4896 4632 4948 4684
rect 5264 4632 5316 4684
rect 5908 4675 5960 4684
rect 5908 4641 5917 4675
rect 5917 4641 5951 4675
rect 5951 4641 5960 4675
rect 5908 4632 5960 4641
rect 7196 4675 7248 4684
rect 7196 4641 7205 4675
rect 7205 4641 7239 4675
rect 7239 4641 7248 4675
rect 7196 4632 7248 4641
rect 8024 4632 8076 4684
rect 10232 4700 10284 4752
rect 12900 4700 12952 4752
rect 13268 4700 13320 4752
rect 13728 4700 13780 4752
rect 14924 4700 14976 4752
rect 15936 4700 15988 4752
rect 16764 4700 16816 4752
rect 18972 4743 19024 4752
rect 9772 4632 9824 4684
rect 12072 4675 12124 4684
rect 12072 4641 12081 4675
rect 12081 4641 12115 4675
rect 12115 4641 12124 4675
rect 12072 4632 12124 4641
rect 12440 4632 12492 4684
rect 16672 4675 16724 4684
rect 16672 4641 16681 4675
rect 16681 4641 16715 4675
rect 16715 4641 16724 4675
rect 16672 4632 16724 4641
rect 18972 4709 18981 4743
rect 18981 4709 19015 4743
rect 19015 4709 19024 4743
rect 18972 4700 19024 4709
rect 21732 4700 21784 4752
rect 2964 4564 3016 4616
rect 3148 4607 3200 4616
rect 3148 4573 3157 4607
rect 3157 4573 3191 4607
rect 3191 4573 3200 4607
rect 3148 4564 3200 4573
rect 5356 4564 5408 4616
rect 1952 4496 2004 4548
rect 5724 4539 5776 4548
rect 5724 4505 5733 4539
rect 5733 4505 5767 4539
rect 5767 4505 5776 4539
rect 5724 4496 5776 4505
rect 7104 4496 7156 4548
rect 14004 4564 14056 4616
rect 16580 4564 16632 4616
rect 16948 4564 17000 4616
rect 17684 4632 17736 4684
rect 18604 4632 18656 4684
rect 18788 4675 18840 4684
rect 18788 4641 18797 4675
rect 18797 4641 18831 4675
rect 18831 4641 18840 4675
rect 18788 4632 18840 4641
rect 18880 4632 18932 4684
rect 18328 4564 18380 4616
rect 22192 4632 22244 4684
rect 22928 4675 22980 4684
rect 22928 4641 22937 4675
rect 22937 4641 22971 4675
rect 22971 4641 22980 4675
rect 22928 4632 22980 4641
rect 26700 4700 26752 4752
rect 29460 4700 29512 4752
rect 24952 4675 25004 4684
rect 24952 4641 24961 4675
rect 24961 4641 24995 4675
rect 24995 4641 25004 4675
rect 24952 4632 25004 4641
rect 25320 4675 25372 4684
rect 25320 4641 25329 4675
rect 25329 4641 25363 4675
rect 25363 4641 25372 4675
rect 25320 4632 25372 4641
rect 27160 4675 27212 4684
rect 27160 4641 27169 4675
rect 27169 4641 27203 4675
rect 27203 4641 27212 4675
rect 27160 4632 27212 4641
rect 28264 4675 28316 4684
rect 28264 4641 28273 4675
rect 28273 4641 28307 4675
rect 28307 4641 28316 4675
rect 28264 4632 28316 4641
rect 29644 4675 29696 4684
rect 22376 4564 22428 4616
rect 23388 4564 23440 4616
rect 25136 4564 25188 4616
rect 26516 4607 26568 4616
rect 26516 4573 26525 4607
rect 26525 4573 26559 4607
rect 26559 4573 26568 4607
rect 26516 4564 26568 4573
rect 27712 4564 27764 4616
rect 29644 4641 29653 4675
rect 29653 4641 29687 4675
rect 29687 4641 29696 4675
rect 29644 4632 29696 4641
rect 30196 4564 30248 4616
rect 5816 4428 5868 4480
rect 9864 4496 9916 4548
rect 10416 4496 10468 4548
rect 16212 4496 16264 4548
rect 16488 4496 16540 4548
rect 27436 4496 27488 4548
rect 8392 4471 8444 4480
rect 8392 4437 8401 4471
rect 8401 4437 8435 4471
rect 8435 4437 8444 4471
rect 8392 4428 8444 4437
rect 8852 4471 8904 4480
rect 8852 4437 8861 4471
rect 8861 4437 8895 4471
rect 8895 4437 8904 4471
rect 8852 4428 8904 4437
rect 9312 4428 9364 4480
rect 16304 4428 16356 4480
rect 17132 4471 17184 4480
rect 17132 4437 17141 4471
rect 17141 4437 17175 4471
rect 17175 4437 17184 4471
rect 17132 4428 17184 4437
rect 19892 4428 19944 4480
rect 24492 4471 24544 4480
rect 24492 4437 24501 4471
rect 24501 4437 24535 4471
rect 24535 4437 24544 4471
rect 24492 4428 24544 4437
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 1676 4267 1728 4276
rect 1676 4233 1685 4267
rect 1685 4233 1719 4267
rect 1719 4233 1728 4267
rect 1676 4224 1728 4233
rect 2872 4267 2924 4276
rect 2872 4233 2881 4267
rect 2881 4233 2915 4267
rect 2915 4233 2924 4267
rect 2872 4224 2924 4233
rect 4528 4267 4580 4276
rect 4528 4233 4537 4267
rect 4537 4233 4571 4267
rect 4571 4233 4580 4267
rect 4528 4224 4580 4233
rect 5724 4224 5776 4276
rect 7104 4267 7156 4276
rect 7104 4233 7113 4267
rect 7113 4233 7147 4267
rect 7147 4233 7156 4267
rect 7104 4224 7156 4233
rect 5908 4156 5960 4208
rect 3148 4088 3200 4140
rect 3700 4063 3752 4072
rect 3700 4029 3709 4063
rect 3709 4029 3743 4063
rect 3743 4029 3752 4063
rect 3700 4020 3752 4029
rect 6000 4088 6052 4140
rect 6644 4156 6696 4208
rect 7380 4088 7432 4140
rect 10232 4224 10284 4276
rect 11980 4224 12032 4276
rect 12348 4224 12400 4276
rect 12624 4224 12676 4276
rect 13728 4267 13780 4276
rect 13728 4233 13737 4267
rect 13737 4233 13771 4267
rect 13771 4233 13780 4267
rect 13728 4224 13780 4233
rect 16304 4267 16356 4276
rect 16304 4233 16313 4267
rect 16313 4233 16347 4267
rect 16347 4233 16356 4267
rect 16304 4224 16356 4233
rect 16396 4224 16448 4276
rect 19892 4267 19944 4276
rect 9956 4156 10008 4208
rect 12072 4156 12124 4208
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 14004 4131 14056 4140
rect 14004 4097 14013 4131
rect 14013 4097 14047 4131
rect 14047 4097 14056 4131
rect 14004 4088 14056 4097
rect 4896 4063 4948 4072
rect 4896 4029 4905 4063
rect 4905 4029 4939 4063
rect 4939 4029 4948 4063
rect 4896 4020 4948 4029
rect 5816 4020 5868 4072
rect 7472 4063 7524 4072
rect 7472 4029 7481 4063
rect 7481 4029 7515 4063
rect 7515 4029 7524 4063
rect 7472 4020 7524 4029
rect 8392 4063 8444 4072
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 8484 4063 8536 4072
rect 8484 4029 8493 4063
rect 8493 4029 8527 4063
rect 8527 4029 8536 4063
rect 8484 4020 8536 4029
rect 9956 4063 10008 4072
rect 1952 3995 2004 4004
rect 1952 3961 1961 3995
rect 1961 3961 1995 3995
rect 1995 3961 2004 3995
rect 1952 3952 2004 3961
rect 2044 3995 2096 4004
rect 2044 3961 2053 3995
rect 2053 3961 2087 3995
rect 2087 3961 2096 3995
rect 2044 3952 2096 3961
rect 4528 3952 4580 4004
rect 3516 3927 3568 3936
rect 3516 3893 3525 3927
rect 3525 3893 3559 3927
rect 3559 3893 3568 3927
rect 3516 3884 3568 3893
rect 6092 3952 6144 4004
rect 6184 3927 6236 3936
rect 6184 3893 6193 3927
rect 6193 3893 6227 3927
rect 6227 3893 6236 3927
rect 6184 3884 6236 3893
rect 7656 3884 7708 3936
rect 8024 3884 8076 3936
rect 9956 4029 9965 4063
rect 9965 4029 9999 4063
rect 9999 4029 10008 4063
rect 9956 4020 10008 4029
rect 10416 4063 10468 4072
rect 10416 4029 10425 4063
rect 10425 4029 10459 4063
rect 10459 4029 10468 4063
rect 10416 4020 10468 4029
rect 12348 4020 12400 4072
rect 12624 4020 12676 4072
rect 13820 4020 13872 4072
rect 15108 4063 15160 4072
rect 15108 4029 15117 4063
rect 15117 4029 15151 4063
rect 15151 4029 15160 4063
rect 16856 4199 16908 4208
rect 15752 4088 15804 4140
rect 16212 4088 16264 4140
rect 16856 4165 16865 4199
rect 16865 4165 16899 4199
rect 16899 4165 16908 4199
rect 16856 4156 16908 4165
rect 16948 4156 17000 4208
rect 18052 4156 18104 4208
rect 18420 4156 18472 4208
rect 16764 4131 16816 4140
rect 16764 4097 16773 4131
rect 16773 4097 16807 4131
rect 16807 4097 16816 4131
rect 16764 4088 16816 4097
rect 19892 4233 19901 4267
rect 19901 4233 19935 4267
rect 19935 4233 19944 4267
rect 19892 4224 19944 4233
rect 24032 4267 24084 4276
rect 24032 4233 24041 4267
rect 24041 4233 24075 4267
rect 24075 4233 24084 4267
rect 24032 4224 24084 4233
rect 26424 4224 26476 4276
rect 27160 4224 27212 4276
rect 19432 4199 19484 4208
rect 19432 4165 19441 4199
rect 19441 4165 19475 4199
rect 19475 4165 19484 4199
rect 19432 4156 19484 4165
rect 24124 4156 24176 4208
rect 29644 4224 29696 4276
rect 35440 4224 35492 4276
rect 27712 4199 27764 4208
rect 27712 4165 27721 4199
rect 27721 4165 27755 4199
rect 27755 4165 27764 4199
rect 27712 4156 27764 4165
rect 28264 4199 28316 4208
rect 28264 4165 28273 4199
rect 28273 4165 28307 4199
rect 28307 4165 28316 4199
rect 28264 4156 28316 4165
rect 15108 4020 15160 4029
rect 17960 4020 18012 4072
rect 18144 4063 18196 4072
rect 18144 4029 18153 4063
rect 18153 4029 18187 4063
rect 18187 4029 18196 4063
rect 18144 4020 18196 4029
rect 18420 4020 18472 4072
rect 21180 4088 21232 4140
rect 22192 4088 22244 4140
rect 22652 4088 22704 4140
rect 23388 4131 23440 4140
rect 23388 4097 23397 4131
rect 23397 4097 23431 4131
rect 23431 4097 23440 4131
rect 23388 4088 23440 4097
rect 25044 4088 25096 4140
rect 25688 4131 25740 4140
rect 25688 4097 25697 4131
rect 25697 4097 25731 4131
rect 25731 4097 25740 4131
rect 25688 4088 25740 4097
rect 28172 4088 28224 4140
rect 29828 4131 29880 4140
rect 29828 4097 29837 4131
rect 29837 4097 29871 4131
rect 29871 4097 29880 4131
rect 29828 4088 29880 4097
rect 21916 4063 21968 4072
rect 9404 3952 9456 4004
rect 9772 3952 9824 4004
rect 16672 3952 16724 4004
rect 19432 3952 19484 4004
rect 20628 3995 20680 4004
rect 20628 3961 20637 3995
rect 20637 3961 20671 3995
rect 20671 3961 20680 3995
rect 20628 3952 20680 3961
rect 8852 3927 8904 3936
rect 8852 3893 8861 3927
rect 8861 3893 8895 3927
rect 8895 3893 8904 3927
rect 8852 3884 8904 3893
rect 9128 3884 9180 3936
rect 9864 3884 9916 3936
rect 11704 3884 11756 3936
rect 15200 3884 15252 3936
rect 16764 3884 16816 3936
rect 18052 3884 18104 3936
rect 18788 3884 18840 3936
rect 19156 3884 19208 3936
rect 20812 3884 20864 3936
rect 21916 4029 21925 4063
rect 21925 4029 21959 4063
rect 21959 4029 21968 4063
rect 21916 4020 21968 4029
rect 22100 4063 22152 4072
rect 22100 4029 22109 4063
rect 22109 4029 22143 4063
rect 22143 4029 22152 4063
rect 22100 4020 22152 4029
rect 22376 4020 22428 4072
rect 24492 4063 24544 4072
rect 24492 4029 24501 4063
rect 24501 4029 24535 4063
rect 24535 4029 24544 4063
rect 24492 4020 24544 4029
rect 22928 3952 22980 4004
rect 23756 3952 23808 4004
rect 24952 3952 25004 4004
rect 26332 3995 26384 4004
rect 26332 3961 26341 3995
rect 26341 3961 26375 3995
rect 26375 3961 26384 3995
rect 26332 3952 26384 3961
rect 26424 3995 26476 4004
rect 26424 3961 26433 3995
rect 26433 3961 26467 3995
rect 26467 3961 26476 3995
rect 26976 3995 27028 4004
rect 26424 3952 26476 3961
rect 26976 3961 26985 3995
rect 26985 3961 27019 3995
rect 27019 3961 27028 3995
rect 26976 3952 27028 3961
rect 28540 4020 28592 4072
rect 30288 4063 30340 4072
rect 30288 4029 30297 4063
rect 30297 4029 30331 4063
rect 30331 4029 30340 4063
rect 30288 4020 30340 4029
rect 22744 3927 22796 3936
rect 22744 3893 22753 3927
rect 22753 3893 22787 3927
rect 22787 3893 22796 3927
rect 22744 3884 22796 3893
rect 25504 3884 25556 3936
rect 30472 3927 30524 3936
rect 30472 3893 30481 3927
rect 30481 3893 30515 3927
rect 30515 3893 30524 3927
rect 30472 3884 30524 3893
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 1768 3723 1820 3732
rect 1768 3689 1777 3723
rect 1777 3689 1811 3723
rect 1811 3689 1820 3723
rect 1768 3680 1820 3689
rect 1952 3680 2004 3732
rect 2964 3680 3016 3732
rect 5448 3680 5500 3732
rect 5816 3723 5868 3732
rect 5816 3689 5825 3723
rect 5825 3689 5859 3723
rect 5859 3689 5868 3723
rect 5816 3680 5868 3689
rect 3792 3612 3844 3664
rect 8208 3680 8260 3732
rect 9220 3723 9272 3732
rect 9220 3689 9229 3723
rect 9229 3689 9263 3723
rect 9263 3689 9272 3723
rect 9220 3680 9272 3689
rect 9680 3680 9732 3732
rect 9956 3680 10008 3732
rect 12440 3680 12492 3732
rect 12624 3723 12676 3732
rect 12624 3689 12633 3723
rect 12633 3689 12667 3723
rect 12667 3689 12676 3723
rect 12624 3680 12676 3689
rect 15936 3723 15988 3732
rect 15936 3689 15945 3723
rect 15945 3689 15979 3723
rect 15979 3689 15988 3723
rect 15936 3680 15988 3689
rect 17592 3723 17644 3732
rect 17592 3689 17601 3723
rect 17601 3689 17635 3723
rect 17635 3689 17644 3723
rect 17592 3680 17644 3689
rect 20628 3723 20680 3732
rect 2136 3544 2188 3596
rect 4252 3544 4304 3596
rect 5080 3587 5132 3596
rect 5080 3553 5089 3587
rect 5089 3553 5123 3587
rect 5123 3553 5132 3587
rect 5080 3544 5132 3553
rect 3700 3476 3752 3528
rect 5632 3544 5684 3596
rect 8852 3612 8904 3664
rect 7380 3587 7432 3596
rect 5264 3476 5316 3528
rect 6184 3476 6236 3528
rect 7380 3553 7389 3587
rect 7389 3553 7423 3587
rect 7423 3553 7432 3587
rect 7380 3544 7432 3553
rect 7656 3587 7708 3596
rect 7656 3553 7665 3587
rect 7665 3553 7699 3587
rect 7699 3553 7708 3587
rect 7656 3544 7708 3553
rect 7472 3519 7524 3528
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 9036 3544 9088 3596
rect 9956 3587 10008 3596
rect 9956 3553 9965 3587
rect 9965 3553 9999 3587
rect 9999 3553 10008 3587
rect 9956 3544 10008 3553
rect 10232 3587 10284 3596
rect 10232 3553 10241 3587
rect 10241 3553 10275 3587
rect 10275 3553 10284 3587
rect 10232 3544 10284 3553
rect 11980 3587 12032 3596
rect 11980 3553 11989 3587
rect 11989 3553 12023 3587
rect 12023 3553 12032 3587
rect 11980 3544 12032 3553
rect 12440 3544 12492 3596
rect 13820 3587 13872 3596
rect 13820 3553 13829 3587
rect 13829 3553 13863 3587
rect 13863 3553 13872 3587
rect 14832 3612 14884 3664
rect 17776 3655 17828 3664
rect 17776 3621 17785 3655
rect 17785 3621 17819 3655
rect 17819 3621 17828 3655
rect 17776 3612 17828 3621
rect 13820 3544 13872 3553
rect 14372 3587 14424 3596
rect 14372 3553 14381 3587
rect 14381 3553 14415 3587
rect 14415 3553 14424 3587
rect 14372 3544 14424 3553
rect 16396 3587 16448 3596
rect 16396 3553 16405 3587
rect 16405 3553 16439 3587
rect 16439 3553 16448 3587
rect 16396 3544 16448 3553
rect 18696 3612 18748 3664
rect 18880 3612 18932 3664
rect 20260 3612 20312 3664
rect 19248 3544 19300 3596
rect 20628 3689 20637 3723
rect 20637 3689 20671 3723
rect 20671 3689 20680 3723
rect 20628 3680 20680 3689
rect 22652 3723 22704 3732
rect 22652 3689 22661 3723
rect 22661 3689 22695 3723
rect 22695 3689 22704 3723
rect 22652 3680 22704 3689
rect 24492 3680 24544 3732
rect 29092 3680 29144 3732
rect 21180 3587 21232 3596
rect 21180 3553 21189 3587
rect 21189 3553 21223 3587
rect 21223 3553 21232 3587
rect 21180 3544 21232 3553
rect 22100 3612 22152 3664
rect 8116 3519 8168 3528
rect 7472 3476 7524 3485
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 9864 3476 9916 3528
rect 12348 3476 12400 3528
rect 17960 3519 18012 3528
rect 17960 3485 17966 3519
rect 17966 3485 18012 3519
rect 17960 3476 18012 3485
rect 18420 3476 18472 3528
rect 19892 3519 19944 3528
rect 19892 3485 19901 3519
rect 19901 3485 19935 3519
rect 19935 3485 19944 3519
rect 19892 3476 19944 3485
rect 20628 3476 20680 3528
rect 22560 3544 22612 3596
rect 21824 3476 21876 3528
rect 24952 3612 25004 3664
rect 28448 3612 28500 3664
rect 23664 3587 23716 3596
rect 23664 3553 23673 3587
rect 23673 3553 23707 3587
rect 23707 3553 23716 3587
rect 23664 3544 23716 3553
rect 24860 3587 24912 3596
rect 24860 3553 24869 3587
rect 24869 3553 24903 3587
rect 24903 3553 24912 3587
rect 24860 3544 24912 3553
rect 26148 3544 26200 3596
rect 27252 3544 27304 3596
rect 27528 3544 27580 3596
rect 16212 3408 16264 3460
rect 18052 3451 18104 3460
rect 18052 3417 18061 3451
rect 18061 3417 18095 3451
rect 18095 3417 18104 3451
rect 18052 3408 18104 3417
rect 18328 3408 18380 3460
rect 22100 3408 22152 3460
rect 26976 3476 27028 3528
rect 30748 3476 30800 3528
rect 27988 3408 28040 3460
rect 30104 3451 30156 3460
rect 30104 3417 30113 3451
rect 30113 3417 30147 3451
rect 30147 3417 30156 3451
rect 30104 3408 30156 3417
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 15200 3340 15252 3392
rect 24584 3383 24636 3392
rect 24584 3349 24593 3383
rect 24593 3349 24627 3383
rect 24627 3349 24636 3383
rect 24584 3340 24636 3349
rect 25228 3383 25280 3392
rect 25228 3349 25237 3383
rect 25237 3349 25271 3383
rect 25271 3349 25280 3383
rect 25228 3340 25280 3349
rect 26240 3383 26292 3392
rect 26240 3349 26249 3383
rect 26249 3349 26283 3383
rect 26283 3349 26292 3383
rect 26240 3340 26292 3349
rect 26332 3340 26384 3392
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 2136 3136 2188 3188
rect 3240 3136 3292 3188
rect 3700 3068 3752 3120
rect 1492 3000 1544 3052
rect 2688 3043 2740 3052
rect 2136 2975 2188 2984
rect 2136 2941 2145 2975
rect 2145 2941 2179 2975
rect 2179 2941 2188 2975
rect 2136 2932 2188 2941
rect 2688 3009 2697 3043
rect 2697 3009 2731 3043
rect 2731 3009 2740 3043
rect 2688 3000 2740 3009
rect 4528 3000 4580 3052
rect 4712 3136 4764 3188
rect 5080 3179 5132 3188
rect 5080 3145 5089 3179
rect 5089 3145 5123 3179
rect 5123 3145 5132 3179
rect 5080 3136 5132 3145
rect 5632 3179 5684 3188
rect 5632 3145 5641 3179
rect 5641 3145 5675 3179
rect 5675 3145 5684 3179
rect 5632 3136 5684 3145
rect 6000 3136 6052 3188
rect 7380 3179 7432 3188
rect 7380 3145 7389 3179
rect 7389 3145 7423 3179
rect 7423 3145 7432 3179
rect 7380 3136 7432 3145
rect 7472 3068 7524 3120
rect 6460 3000 6512 3052
rect 6276 2975 6328 2984
rect 6276 2941 6285 2975
rect 6285 2941 6319 2975
rect 6319 2941 6328 2975
rect 6276 2932 6328 2941
rect 7196 2932 7248 2984
rect 4344 2864 4396 2916
rect 7840 2932 7892 2984
rect 9404 3136 9456 3188
rect 9956 3136 10008 3188
rect 13084 3136 13136 3188
rect 14004 3136 14056 3188
rect 15660 3136 15712 3188
rect 17776 3136 17828 3188
rect 18236 3179 18288 3188
rect 18236 3145 18245 3179
rect 18245 3145 18279 3179
rect 18279 3145 18288 3179
rect 18236 3136 18288 3145
rect 23664 3136 23716 3188
rect 27252 3179 27304 3188
rect 27252 3145 27261 3179
rect 27261 3145 27295 3179
rect 27295 3145 27304 3179
rect 27252 3136 27304 3145
rect 27528 3136 27580 3188
rect 27988 3179 28040 3188
rect 27988 3145 27997 3179
rect 27997 3145 28031 3179
rect 28031 3145 28040 3179
rect 27988 3136 28040 3145
rect 30748 3179 30800 3188
rect 30748 3145 30757 3179
rect 30757 3145 30791 3179
rect 30791 3145 30800 3179
rect 30748 3136 30800 3145
rect 10232 3111 10284 3120
rect 10232 3077 10241 3111
rect 10241 3077 10275 3111
rect 10275 3077 10284 3111
rect 10232 3068 10284 3077
rect 15108 3111 15160 3120
rect 15108 3077 15117 3111
rect 15117 3077 15151 3111
rect 15151 3077 15160 3111
rect 15108 3068 15160 3077
rect 16212 3068 16264 3120
rect 17960 3068 18012 3120
rect 9220 2975 9272 2984
rect 9220 2941 9229 2975
rect 9229 2941 9263 2975
rect 9263 2941 9272 2975
rect 9220 2932 9272 2941
rect 13820 3000 13872 3052
rect 15200 3043 15252 3052
rect 15200 3009 15209 3043
rect 15209 3009 15243 3043
rect 15243 3009 15252 3043
rect 15200 3000 15252 3009
rect 16764 3000 16816 3052
rect 18420 3000 18472 3052
rect 23480 3111 23532 3120
rect 23480 3077 23489 3111
rect 23489 3077 23523 3111
rect 23523 3077 23532 3111
rect 23480 3068 23532 3077
rect 19432 3000 19484 3052
rect 21824 3000 21876 3052
rect 22100 3000 22152 3052
rect 11428 2975 11480 2984
rect 11428 2941 11446 2975
rect 11446 2941 11480 2975
rect 11428 2932 11480 2941
rect 4252 2839 4304 2848
rect 4252 2805 4261 2839
rect 4261 2805 4295 2839
rect 4295 2805 4304 2839
rect 4252 2796 4304 2805
rect 7104 2839 7156 2848
rect 7104 2805 7113 2839
rect 7113 2805 7147 2839
rect 7147 2805 7156 2839
rect 7104 2796 7156 2805
rect 8392 2864 8444 2916
rect 12256 2907 12308 2916
rect 9312 2839 9364 2848
rect 9312 2805 9321 2839
rect 9321 2805 9355 2839
rect 9355 2805 9364 2839
rect 9312 2796 9364 2805
rect 11980 2796 12032 2848
rect 12256 2873 12265 2907
rect 12265 2873 12299 2907
rect 12299 2873 12308 2907
rect 12256 2864 12308 2873
rect 13912 2864 13964 2916
rect 14924 2932 14976 2984
rect 16396 2975 16448 2984
rect 16396 2941 16405 2975
rect 16405 2941 16439 2975
rect 16439 2941 16448 2975
rect 16396 2932 16448 2941
rect 16672 2975 16724 2984
rect 16672 2941 16681 2975
rect 16681 2941 16715 2975
rect 16715 2941 16724 2975
rect 16672 2932 16724 2941
rect 18328 2932 18380 2984
rect 14832 2907 14884 2916
rect 14832 2873 14841 2907
rect 14841 2873 14875 2907
rect 14875 2873 14884 2907
rect 14832 2864 14884 2873
rect 19248 2796 19300 2848
rect 19432 2907 19484 2916
rect 19432 2873 19441 2907
rect 19441 2873 19475 2907
rect 19475 2873 19484 2907
rect 19984 2907 20036 2916
rect 19432 2864 19484 2873
rect 19984 2873 19993 2907
rect 19993 2873 20027 2907
rect 20027 2873 20036 2907
rect 19984 2864 20036 2873
rect 22744 2932 22796 2984
rect 24584 3000 24636 3052
rect 26332 3043 26384 3052
rect 26332 3009 26341 3043
rect 26341 3009 26375 3043
rect 26375 3009 26384 3043
rect 26332 3000 26384 3009
rect 27712 3000 27764 3052
rect 29460 3043 29512 3052
rect 29460 3009 29469 3043
rect 29469 3009 29503 3043
rect 29503 3009 29512 3043
rect 29460 3000 29512 3009
rect 30104 3043 30156 3052
rect 30104 3009 30113 3043
rect 30113 3009 30147 3043
rect 30147 3009 30156 3043
rect 30104 3000 30156 3009
rect 20260 2907 20312 2916
rect 20260 2873 20269 2907
rect 20269 2873 20303 2907
rect 20303 2873 20312 2907
rect 20260 2864 20312 2873
rect 20628 2839 20680 2848
rect 20628 2805 20637 2839
rect 20637 2805 20671 2839
rect 20671 2805 20680 2839
rect 20628 2796 20680 2805
rect 20904 2864 20956 2916
rect 23985 2907 24037 2916
rect 23985 2873 23994 2907
rect 23994 2873 24028 2907
rect 24028 2873 24037 2907
rect 23985 2864 24037 2873
rect 26516 2864 26568 2916
rect 26976 2907 27028 2916
rect 26976 2873 26985 2907
rect 26985 2873 27019 2907
rect 27019 2873 27028 2907
rect 26976 2864 27028 2873
rect 29552 2907 29604 2916
rect 29552 2873 29561 2907
rect 29561 2873 29595 2907
rect 29595 2873 29604 2907
rect 29552 2864 29604 2873
rect 21456 2796 21508 2848
rect 21916 2796 21968 2848
rect 22100 2839 22152 2848
rect 22100 2805 22109 2839
rect 22109 2805 22143 2839
rect 22143 2805 22152 2839
rect 22100 2796 22152 2805
rect 22560 2796 22612 2848
rect 23572 2796 23624 2848
rect 24860 2839 24912 2848
rect 24860 2805 24869 2839
rect 24869 2805 24903 2839
rect 24903 2805 24912 2839
rect 24860 2796 24912 2805
rect 28448 2796 28500 2848
rect 29828 2796 29880 2848
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 2136 2592 2188 2644
rect 2964 2592 3016 2644
rect 7472 2592 7524 2644
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 11888 2592 11940 2644
rect 14740 2592 14792 2644
rect 15108 2592 15160 2644
rect 16396 2592 16448 2644
rect 16764 2592 16816 2644
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 18604 2592 18656 2644
rect 7840 2567 7892 2576
rect 7840 2533 7849 2567
rect 7849 2533 7883 2567
rect 7883 2533 7892 2567
rect 7840 2524 7892 2533
rect 13820 2524 13872 2576
rect 18880 2524 18932 2576
rect 112 2456 164 2508
rect 5540 2456 5592 2508
rect 7104 2456 7156 2508
rect 8024 2456 8076 2508
rect 8116 2456 8168 2508
rect 10048 2499 10100 2508
rect 10048 2465 10057 2499
rect 10057 2465 10091 2499
rect 10091 2465 10100 2499
rect 10048 2456 10100 2465
rect 10232 2499 10284 2508
rect 10232 2465 10241 2499
rect 10241 2465 10275 2499
rect 10275 2465 10284 2499
rect 10232 2456 10284 2465
rect 8300 2388 8352 2440
rect 13360 2456 13412 2508
rect 14832 2456 14884 2508
rect 15200 2456 15252 2508
rect 16672 2456 16724 2508
rect 19156 2592 19208 2644
rect 20904 2635 20956 2644
rect 20904 2601 20913 2635
rect 20913 2601 20947 2635
rect 20947 2601 20956 2635
rect 20904 2592 20956 2601
rect 21640 2635 21692 2644
rect 21640 2601 21649 2635
rect 21649 2601 21683 2635
rect 21683 2601 21692 2635
rect 21640 2592 21692 2601
rect 21916 2592 21968 2644
rect 23756 2635 23808 2644
rect 23756 2601 23765 2635
rect 23765 2601 23799 2635
rect 23799 2601 23808 2635
rect 23756 2592 23808 2601
rect 25228 2635 25280 2644
rect 19708 2567 19760 2576
rect 19708 2533 19717 2567
rect 19717 2533 19751 2567
rect 19751 2533 19760 2567
rect 19708 2524 19760 2533
rect 19984 2524 20036 2576
rect 23572 2524 23624 2576
rect 25228 2601 25237 2635
rect 25237 2601 25271 2635
rect 25271 2601 25280 2635
rect 25228 2592 25280 2601
rect 26240 2592 26292 2644
rect 29092 2635 29144 2644
rect 29092 2601 29101 2635
rect 29101 2601 29135 2635
rect 29135 2601 29144 2635
rect 29092 2592 29144 2601
rect 29460 2635 29512 2644
rect 29460 2601 29469 2635
rect 29469 2601 29503 2635
rect 29503 2601 29512 2635
rect 29460 2592 29512 2601
rect 24492 2524 24544 2576
rect 24032 2456 24084 2508
rect 24860 2499 24912 2508
rect 24860 2465 24869 2499
rect 24869 2465 24903 2499
rect 24903 2465 24912 2499
rect 24860 2456 24912 2465
rect 27436 2456 27488 2508
rect 29552 2524 29604 2576
rect 29828 2499 29880 2508
rect 29828 2465 29837 2499
rect 29837 2465 29871 2499
rect 29871 2465 29880 2499
rect 29828 2456 29880 2465
rect 30104 2456 30156 2508
rect 18972 2388 19024 2440
rect 7288 2320 7340 2372
rect 10048 2320 10100 2372
rect 8392 2252 8444 2304
rect 12348 2252 12400 2304
rect 13360 2295 13412 2304
rect 13360 2261 13369 2295
rect 13369 2261 13403 2295
rect 13403 2261 13412 2295
rect 13360 2252 13412 2261
rect 15200 2295 15252 2304
rect 15200 2261 15209 2295
rect 15209 2261 15243 2295
rect 15243 2261 15252 2295
rect 15200 2252 15252 2261
rect 19248 2252 19300 2304
rect 21456 2252 21508 2304
rect 24492 2252 24544 2304
rect 38384 2320 38436 2372
rect 27436 2295 27488 2304
rect 27436 2261 27445 2295
rect 27445 2261 27479 2295
rect 27479 2261 27488 2295
rect 27436 2252 27488 2261
rect 28264 2252 28316 2304
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
rect 25412 76 25464 128
rect 31668 76 31720 128
<< metal2 >>
rect 2502 15586 2558 16000
rect 2502 15558 2820 15586
rect 2502 15520 2558 15558
rect 2686 15056 2742 15065
rect 2686 14991 2742 15000
rect 1582 14240 1638 14249
rect 1582 14175 1638 14184
rect 110 13800 166 13809
rect 110 13735 166 13744
rect 124 12986 152 13735
rect 1596 13530 1624 14175
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 112 12980 164 12986
rect 112 12922 164 12928
rect 2424 12646 2452 13330
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 110 12064 166 12073
rect 110 11999 166 12008
rect 124 11898 152 11999
rect 112 11892 164 11898
rect 112 11834 164 11840
rect 1412 11558 1440 12242
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1412 10713 1440 11494
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1584 11008 1636 11014
rect 1584 10950 1636 10956
rect 1596 10849 1624 10950
rect 1582 10840 1638 10849
rect 1582 10775 1638 10784
rect 1398 10704 1454 10713
rect 1398 10639 1454 10648
rect 112 10464 164 10470
rect 112 10406 164 10412
rect 124 10305 152 10406
rect 110 10296 166 10305
rect 110 10231 166 10240
rect 754 6760 810 6769
rect 754 6695 810 6704
rect 768 3641 796 6695
rect 1412 4593 1440 10639
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1504 9382 1532 10066
rect 1688 9926 1716 11154
rect 2148 10606 2176 12582
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1398 4584 1454 4593
rect 1398 4519 1454 4528
rect 754 3632 810 3641
rect 754 3567 810 3576
rect 1504 3058 1532 9318
rect 1688 9178 1716 9862
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1688 8634 1716 8978
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1688 8537 1716 8570
rect 1674 8528 1730 8537
rect 1674 8463 1730 8472
rect 1582 7984 1638 7993
rect 1780 7954 1808 10202
rect 2056 8906 2084 10406
rect 2226 10024 2282 10033
rect 2226 9959 2282 9968
rect 2044 8900 2096 8906
rect 2044 8842 2096 8848
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1872 8498 1900 8774
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 1582 7919 1638 7928
rect 1768 7948 1820 7954
rect 1596 6458 1624 7919
rect 1768 7890 1820 7896
rect 1780 7002 1808 7890
rect 2148 7274 2176 8026
rect 2240 7857 2268 9959
rect 2332 9586 2360 12038
rect 2424 10742 2452 12582
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 2412 10736 2464 10742
rect 2412 10678 2464 10684
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2424 9722 2452 10066
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2412 9444 2464 9450
rect 2332 9404 2412 9432
rect 2332 8838 2360 9404
rect 2412 9386 2464 9392
rect 2516 8974 2544 12038
rect 2700 11354 2728 14991
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2792 10266 2820 15558
rect 5908 15564 5960 15570
rect 7470 15564 7526 16000
rect 12438 15586 12494 16000
rect 17498 15586 17554 16000
rect 22466 15586 22522 16000
rect 27434 15586 27490 16000
rect 7470 15520 7472 15564
rect 5908 15506 5960 15512
rect 7524 15520 7526 15564
rect 12176 15558 12494 15586
rect 7472 15506 7524 15512
rect 5814 12336 5870 12345
rect 3056 12300 3108 12306
rect 5814 12271 5870 12280
rect 3056 12242 3108 12248
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2596 9104 2648 9110
rect 2596 9046 2648 9052
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2332 8362 2360 8774
rect 2516 8566 2544 8910
rect 2608 8634 2636 9046
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2504 8560 2556 8566
rect 2504 8502 2556 8508
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2700 8090 2728 8298
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2226 7848 2282 7857
rect 2226 7783 2282 7792
rect 2136 7268 2188 7274
rect 2136 7210 2188 7216
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 2148 6934 2176 7210
rect 2884 7002 2912 11562
rect 3068 11558 3096 12242
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3068 10033 3096 11494
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3344 10470 3372 11154
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3054 10024 3110 10033
rect 3054 9959 3110 9968
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2976 8498 3004 8910
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2136 6928 2188 6934
rect 2136 6870 2188 6876
rect 2148 6458 2176 6870
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2056 6225 2084 6258
rect 2042 6216 2098 6225
rect 2042 6151 2098 6160
rect 2148 5914 2176 6394
rect 2884 6322 2912 6938
rect 3068 6730 3096 9386
rect 3160 8945 3188 10406
rect 3146 8936 3202 8945
rect 3146 8871 3202 8880
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3160 7546 3188 8570
rect 3344 8537 3372 10406
rect 3330 8528 3386 8537
rect 3330 8463 3386 8472
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2976 6118 3004 6598
rect 3068 6322 3096 6666
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3160 6186 3188 7482
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2044 5840 2096 5846
rect 2044 5782 2096 5788
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2056 5370 2084 5782
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1688 4282 1716 4626
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1688 4185 1716 4218
rect 1674 4176 1730 4185
rect 1674 4111 1730 4120
rect 1780 3738 1808 5102
rect 2056 4826 2084 5306
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 1952 4548 2004 4554
rect 1952 4490 2004 4496
rect 1964 4010 1992 4490
rect 2056 4010 2084 4762
rect 2134 4040 2190 4049
rect 1952 4004 2004 4010
rect 1952 3946 2004 3952
rect 2044 4004 2096 4010
rect 2134 3975 2190 3984
rect 2044 3946 2096 3952
rect 1964 3738 1992 3946
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 2148 3602 2176 3975
rect 2136 3596 2188 3602
rect 2136 3538 2188 3544
rect 2148 3194 2176 3538
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 2148 2990 2176 3130
rect 2700 3058 2728 5782
rect 2872 4752 2924 4758
rect 2976 4740 3004 6054
rect 3160 5914 3188 6122
rect 3252 5914 3280 6734
rect 3436 5914 3464 10474
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3528 7342 3556 7686
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3252 5030 3280 5646
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 2924 4712 3004 4740
rect 2872 4694 2924 4700
rect 2884 4282 2912 4694
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2976 3738 3004 4558
rect 3160 4146 3188 4558
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 2148 2650 2176 2926
rect 2976 2650 3004 3674
rect 3252 3194 3280 4966
rect 3528 3942 3556 7278
rect 3620 6225 3648 11494
rect 4724 11218 4752 11630
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 8022 3832 10950
rect 4724 10810 4752 11154
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 3700 7268 3752 7274
rect 3700 7210 3752 7216
rect 3606 6216 3662 6225
rect 3606 6151 3662 6160
rect 3712 5370 3740 7210
rect 3896 6798 3924 10406
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3974 8800 4030 8809
rect 3974 8735 4030 8744
rect 3988 8634 4016 8735
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4080 8090 4108 9318
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4080 7410 4108 8026
rect 4252 8016 4304 8022
rect 4172 7976 4252 8004
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4172 6934 4200 7976
rect 4252 7958 4304 7964
rect 4356 7868 4384 10406
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5184 9722 5212 10066
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4264 7840 4384 7868
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 4172 6458 4200 6870
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 3792 5772 3844 5778
rect 3792 5714 3844 5720
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3712 4826 3740 5102
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3712 3534 3740 4014
rect 3804 3670 3832 5714
rect 4264 4154 4292 7840
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4448 6458 4476 6734
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4448 6186 4476 6258
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 4356 5914 4384 6122
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4528 4752 4580 4758
rect 4528 4694 4580 4700
rect 4540 4282 4568 4694
rect 4632 4593 4660 8366
rect 4724 8294 4752 8774
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4618 4584 4674 4593
rect 4618 4519 4674 4528
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4540 4154 4568 4218
rect 4264 4126 4384 4154
rect 4540 4126 4660 4154
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3712 3126 3740 3470
rect 3700 3120 3752 3126
rect 3700 3062 3752 3068
rect 4264 2854 4292 3538
rect 4356 2922 4384 4126
rect 4632 4049 4660 4126
rect 4618 4040 4674 4049
rect 4528 4004 4580 4010
rect 4618 3975 4674 3984
rect 4528 3946 4580 3952
rect 4540 3058 4568 3946
rect 4724 3194 4752 8230
rect 4816 8022 4844 8910
rect 5092 8022 5120 9046
rect 5184 8974 5212 9658
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5184 8566 5212 8910
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 5368 7546 5396 8298
rect 5460 7750 5488 8434
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 5092 6934 5120 7142
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 5460 6798 5488 7686
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 4804 6180 4856 6186
rect 4804 6122 4856 6128
rect 4816 5778 4844 6122
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 5078 5672 5134 5681
rect 5078 5607 5134 5616
rect 5356 5636 5408 5642
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4908 4078 4936 4626
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4908 3913 4936 4014
rect 4894 3904 4950 3913
rect 4894 3839 4950 3848
rect 5092 3602 5120 5607
rect 5356 5578 5408 5584
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 5092 3194 5120 3538
rect 5276 3534 5304 4626
rect 5368 4622 5396 5578
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5460 3738 5488 4762
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 112 2508 164 2514
rect 112 2450 164 2456
rect 124 2281 152 2450
rect 110 2272 166 2281
rect 110 2207 166 2216
rect 4264 2009 4292 2790
rect 4250 2000 4306 2009
rect 4250 1935 4306 1944
rect 4356 1057 4384 2858
rect 4342 1048 4398 1057
rect 4342 983 4398 992
rect 1674 82 1730 480
rect 1950 368 2006 377
rect 1950 303 2006 312
rect 1964 82 1992 303
rect 1674 54 1992 82
rect 4986 82 5042 480
rect 5276 82 5304 3470
rect 5552 2514 5580 8842
rect 5828 8090 5856 12271
rect 5920 9722 5948 15506
rect 7484 15475 7512 15506
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 6642 11792 6698 11801
rect 10152 11762 10180 12038
rect 6642 11727 6698 11736
rect 8300 11756 8352 11762
rect 6656 11694 6684 11727
rect 8300 11698 8352 11704
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 7622 10908 7918 10928
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5644 7410 5672 7890
rect 5920 7478 5948 9454
rect 5908 7472 5960 7478
rect 5908 7414 5960 7420
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5736 4826 5764 5646
rect 5828 5370 5856 5782
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 6012 4758 6040 9454
rect 6564 9110 6592 10406
rect 7196 9444 7248 9450
rect 7300 9432 7328 10406
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 8036 9674 8064 10066
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7852 9646 8064 9674
rect 7392 9518 7420 9590
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7248 9404 7328 9432
rect 7196 9386 7248 9392
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6552 9104 6604 9110
rect 6552 9046 6604 9052
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6564 8634 6592 9046
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6656 8090 6684 9046
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6748 6866 6776 9318
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6932 8498 6960 9114
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6840 8022 6868 8230
rect 7208 8022 7236 8298
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6748 5914 6776 6802
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6656 5302 6684 5646
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6380 4758 6408 5102
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 6368 4752 6420 4758
rect 6368 4694 6420 4700
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5736 4282 5764 4490
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5828 4078 5856 4422
rect 5920 4214 5948 4626
rect 5908 4208 5960 4214
rect 5908 4150 5960 4156
rect 6090 4176 6146 4185
rect 6000 4140 6052 4146
rect 6090 4111 6146 4120
rect 6000 4082 6052 4088
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5828 3738 5856 4014
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5644 3194 5672 3538
rect 6012 3194 6040 4082
rect 6104 4010 6132 4111
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6196 3534 6224 3878
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6274 3088 6330 3097
rect 6472 3058 6500 4966
rect 6656 4214 6684 5238
rect 6840 4826 6868 7278
rect 6932 7206 6960 7822
rect 7208 7274 7236 7958
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 6932 5914 6960 7142
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7024 6322 7052 6598
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7024 6186 7052 6258
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7116 5778 7144 7142
rect 7208 6934 7236 7210
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7208 6458 7236 6870
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7116 4282 7144 4490
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 7208 3398 7236 4626
rect 7300 3913 7328 9404
rect 7392 7886 7420 9454
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7392 5302 7420 7822
rect 7484 6361 7512 9386
rect 7852 9382 7880 9646
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7852 8906 7880 9318
rect 8128 9042 8156 11018
rect 8312 10810 8340 11698
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 7840 8900 7892 8906
rect 7892 8860 8064 8888
rect 7840 8842 7892 8848
rect 8036 8809 8064 8860
rect 8022 8800 8078 8809
rect 7622 8732 7918 8752
rect 8022 8735 8078 8744
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 8128 8634 8156 8978
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 8036 6662 8064 7278
rect 8116 7268 8168 7274
rect 8116 7210 8168 7216
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7622 6480 7918 6500
rect 7470 6352 7526 6361
rect 7470 6287 7526 6296
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 8128 5098 8156 7210
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7286 3904 7342 3913
rect 7286 3839 7342 3848
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 6274 3023 6330 3032
rect 6460 3052 6512 3058
rect 6288 2990 6316 3023
rect 6460 2994 6512 3000
rect 7208 2990 7236 3334
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7116 2514 7144 2790
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7300 2378 7328 3839
rect 7392 3602 7420 4082
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7392 3194 7420 3538
rect 7484 3534 7512 4014
rect 8036 3942 8064 4626
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7668 3602 7696 3878
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7484 3126 7512 3470
rect 7622 3292 7918 3312
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7484 2650 7512 3062
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7852 2582 7880 2926
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 8036 2514 8064 3878
rect 8220 3738 8248 10542
rect 8588 10470 8616 11154
rect 10060 11014 10088 11154
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8404 9489 8432 10066
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 8864 9722 8892 9862
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 9048 9586 9076 9862
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 8390 9480 8446 9489
rect 8390 9415 8392 9424
rect 8444 9415 8446 9424
rect 8392 9386 8444 9392
rect 8404 9355 8432 9386
rect 8496 9042 8524 9522
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8496 8634 8524 8978
rect 8772 8838 8800 9386
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 9048 8634 9076 9522
rect 8484 8628 8536 8634
rect 8404 8588 8484 8616
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8128 2514 8156 3470
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7622 2128 7918 2148
rect 4986 54 5304 82
rect 8036 82 8064 2450
rect 8312 2446 8340 7346
rect 8404 6458 8432 8588
rect 8484 8570 8536 8576
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 9048 7410 9076 7890
rect 9508 7857 9536 8366
rect 9494 7848 9550 7857
rect 9494 7783 9550 7792
rect 9600 7546 9628 9998
rect 9692 9625 9720 10406
rect 10060 9926 10088 10950
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9678 9616 9734 9625
rect 10152 9586 10180 11290
rect 10428 11218 10456 11494
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10244 10538 10272 10950
rect 10428 10742 10456 11154
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 9678 9551 9734 9560
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9784 8362 9812 9318
rect 10152 9178 10180 9522
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10244 9110 10272 10474
rect 10336 10266 10364 10474
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10336 9518 10364 10202
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10520 9722 10548 9998
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9968 8634 9996 8978
rect 10612 8838 10640 10134
rect 10796 9178 10824 11562
rect 11164 11558 11192 12242
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11072 9994 11100 10474
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 10980 9586 11008 9930
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10612 8634 10640 8774
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10796 8498 10824 9114
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 8634 11100 8910
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9784 7750 9812 8298
rect 10506 7984 10562 7993
rect 10506 7919 10562 7928
rect 10784 7948 10836 7954
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8404 6186 8432 6394
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8404 5778 8432 6122
rect 8496 6118 8524 6598
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8588 5574 8616 6802
rect 9048 6662 9076 7346
rect 9784 6934 9812 7686
rect 9954 7440 10010 7449
rect 9864 7404 9916 7410
rect 9954 7375 10010 7384
rect 9864 7346 9916 7352
rect 9876 7313 9904 7346
rect 9862 7304 9918 7313
rect 9862 7239 9918 7248
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 6322 9076 6598
rect 9692 6458 9720 6734
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9784 6390 9812 6870
rect 9968 6769 9996 7375
rect 10060 7342 10088 7822
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10152 7290 10180 7414
rect 10244 7410 10272 7482
rect 10232 7404 10284 7410
rect 10416 7404 10468 7410
rect 10232 7346 10284 7352
rect 10336 7364 10416 7392
rect 10336 7290 10364 7364
rect 10416 7346 10468 7352
rect 10152 7262 10364 7290
rect 10416 7268 10468 7274
rect 10416 7210 10468 7216
rect 10048 7200 10100 7206
rect 10140 7200 10192 7206
rect 10100 7160 10140 7188
rect 10048 7142 10100 7148
rect 10140 7142 10192 7148
rect 10152 6866 10180 7142
rect 10428 7002 10456 7210
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 9954 6760 10010 6769
rect 9954 6695 10010 6704
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8680 6089 8708 6190
rect 9784 6118 9812 6326
rect 9772 6112 9824 6118
rect 8666 6080 8722 6089
rect 9772 6054 9824 6060
rect 8666 6015 8722 6024
rect 8680 5914 8708 6015
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8680 5370 8708 5850
rect 9784 5846 9812 6054
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8864 4486 8892 5102
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8404 4078 8432 4422
rect 9048 4185 9076 5510
rect 9692 4826 9720 5646
rect 9784 5370 9812 5782
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9784 5098 9812 5306
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9034 4176 9090 4185
rect 9034 4111 9090 4120
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8404 2922 8432 4014
rect 8496 3534 8524 4014
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8864 3670 8892 3878
rect 8852 3664 8904 3670
rect 8852 3606 8904 3612
rect 9048 3602 9076 4111
rect 9126 4040 9182 4049
rect 9126 3975 9182 3984
rect 9140 3942 9168 3975
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 9232 2990 9260 3674
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8404 2310 8432 2858
rect 9324 2854 9352 4422
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9416 3194 9444 3946
rect 9692 3738 9720 4762
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9784 4010 9812 4626
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9876 3942 9904 4490
rect 9968 4214 9996 6394
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 9956 4208 10008 4214
rect 9956 4150 10008 4156
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9876 3534 9904 3878
rect 9968 3738 9996 4014
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9968 3194 9996 3538
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 10060 2650 10088 4966
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 10244 4282 10272 4694
rect 10428 4554 10456 5714
rect 10520 5001 10548 7919
rect 10784 7890 10836 7896
rect 10796 7478 10824 7890
rect 10784 7472 10836 7478
rect 11164 7449 11192 11494
rect 11440 10198 11468 12038
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11532 10674 11560 11086
rect 11624 10810 11652 11222
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11624 10266 11652 10746
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11428 10192 11480 10198
rect 11428 10134 11480 10140
rect 11440 9722 11468 10134
rect 11624 9722 11652 10202
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11624 9178 11652 9658
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11256 8022 11284 8366
rect 11440 8362 11468 9114
rect 11716 9042 11744 10746
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11992 7936 12020 11698
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12084 9994 12112 11018
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 12176 8090 12204 15558
rect 12438 15520 12494 15558
rect 17144 15558 17554 15586
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10606 12480 10950
rect 13004 10742 13032 11154
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 12992 10736 13044 10742
rect 12992 10678 13044 10684
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12360 9654 12388 9998
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12268 9178 12296 9522
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12072 7948 12124 7954
rect 11992 7908 12072 7936
rect 12072 7890 12124 7896
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 10784 7414 10836 7420
rect 11150 7440 11206 7449
rect 11150 7375 11206 7384
rect 10966 7304 11022 7313
rect 12084 7290 12112 7890
rect 12176 7546 12204 7890
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 12348 7336 12400 7342
rect 12162 7304 12218 7313
rect 12084 7262 12162 7290
rect 10966 7239 11022 7248
rect 12348 7278 12400 7284
rect 12162 7239 12218 7248
rect 10980 7206 11008 7239
rect 12176 7206 12204 7239
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10888 6186 10916 6598
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10796 5642 10824 6122
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 11992 5574 12020 6734
rect 12176 6390 12204 6870
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 12084 5370 12112 5850
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 11428 5296 11480 5302
rect 11428 5238 11480 5244
rect 11440 5137 11468 5238
rect 11426 5128 11482 5137
rect 11426 5063 11482 5072
rect 10506 4992 10562 5001
rect 10506 4927 10562 4936
rect 12176 4826 12204 5646
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 11426 4584 11482 4593
rect 10416 4548 10468 4554
rect 11426 4519 11482 4528
rect 10416 4490 10468 4496
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10428 4078 10456 4490
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10244 3126 10272 3538
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10244 2514 10272 3062
rect 11440 2990 11468 4519
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 10060 2378 10088 2450
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 8298 82 8354 480
rect 8036 54 8354 82
rect 1674 0 1730 54
rect 4986 0 5042 54
rect 8298 0 8354 54
rect 11610 82 11666 480
rect 11716 82 11744 3878
rect 11900 2650 11928 4762
rect 12072 4684 12124 4690
rect 12268 4672 12296 6326
rect 12360 6225 12388 7278
rect 12452 7274 12480 10542
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12544 8634 12572 10406
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12820 8430 12848 8774
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 13004 8090 13032 10678
rect 13188 10674 13216 11018
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13176 9988 13228 9994
rect 13176 9930 13228 9936
rect 13188 8974 13216 9930
rect 13648 9586 13676 10202
rect 14200 10130 14228 10542
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13188 8090 13216 8910
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 12440 7268 12492 7274
rect 12440 7210 12492 7216
rect 12346 6216 12402 6225
rect 12402 6174 12572 6202
rect 12346 6151 12402 6160
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12360 4826 12388 5510
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12124 4644 12296 4672
rect 12440 4684 12492 4690
rect 12072 4626 12124 4632
rect 12440 4626 12492 4632
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11992 3602 12020 4218
rect 12084 4214 12112 4626
rect 12452 4593 12480 4626
rect 12438 4584 12494 4593
rect 12438 4519 12494 4528
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12072 4208 12124 4214
rect 12072 4150 12124 4156
rect 12360 4078 12388 4218
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12452 3738 12480 4519
rect 12544 4185 12572 6174
rect 12636 4282 12664 8026
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 5846 12940 7142
rect 13464 6390 13492 8774
rect 13556 7993 13584 9454
rect 13832 9194 13860 10066
rect 14200 9654 14228 10066
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13740 9166 13860 9194
rect 13740 8838 13768 9166
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13832 8634 13860 9046
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13542 7984 13598 7993
rect 13542 7919 13598 7928
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13648 7274 13676 7890
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13832 7410 13860 7686
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13636 7268 13688 7274
rect 13636 7210 13688 7216
rect 13452 6384 13504 6390
rect 13648 6361 13676 7210
rect 13452 6326 13504 6332
rect 13634 6352 13690 6361
rect 13634 6287 13690 6296
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12912 4758 12940 4966
rect 12900 4752 12952 4758
rect 12900 4694 12952 4700
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12530 4176 12586 4185
rect 13004 4146 13032 6190
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 13096 5914 13124 6122
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13452 5840 13504 5846
rect 13452 5782 13504 5788
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 13188 4826 13216 5034
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13188 4154 13216 4762
rect 13280 4758 13308 5034
rect 13464 4826 13492 5782
rect 13832 5642 13860 7346
rect 13924 5914 13952 9318
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14004 7268 14056 7274
rect 14004 7210 14056 7216
rect 14016 7002 14044 7210
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 14016 6458 14044 6938
rect 14108 6934 14136 7890
rect 14200 7546 14228 9590
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 14660 8022 14688 8366
rect 14648 8016 14700 8022
rect 14648 7958 14700 7964
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14568 7546 14596 7822
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14200 7002 14228 7482
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 14096 6928 14148 6934
rect 14096 6870 14148 6876
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 14752 6322 14780 6802
rect 14844 6798 14872 10406
rect 15120 10062 15148 10474
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15028 9178 15056 9522
rect 15212 9518 15240 10474
rect 15396 9994 15424 10610
rect 15488 10538 15516 11154
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 15396 9110 15424 9930
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15488 7546 15516 10474
rect 15580 10198 15608 11154
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 15304 6458 15332 7278
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14108 6089 14136 6190
rect 15304 6118 15332 6394
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 15292 6112 15344 6118
rect 14094 6080 14150 6089
rect 15292 6054 15344 6060
rect 14094 6015 14150 6024
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 14556 5840 14608 5846
rect 14556 5782 14608 5788
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13832 5166 13860 5578
rect 14568 5370 14596 5782
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 13820 5160 13872 5166
rect 14568 5137 14596 5306
rect 14752 5234 14780 5510
rect 14844 5234 14872 5646
rect 15396 5574 15424 6190
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14832 5228 14884 5234
rect 14884 5188 14964 5216
rect 14832 5170 14884 5176
rect 13820 5102 13872 5108
rect 14554 5128 14610 5137
rect 14554 5063 14610 5072
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13740 4282 13768 4694
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 12530 4111 12586 4120
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13096 4126 13216 4154
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12636 3738 12664 4014
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12452 3602 12480 3674
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 11992 2854 12020 3538
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12256 2916 12308 2922
rect 12256 2858 12308 2864
rect 11980 2848 12032 2854
rect 12268 2825 12296 2858
rect 11980 2790 12032 2796
rect 12254 2816 12310 2825
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11992 2281 12020 2790
rect 12254 2751 12310 2760
rect 12360 2553 12388 3470
rect 13096 3194 13124 4126
rect 13832 4078 13860 4966
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14289 4848 14585 4868
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14016 4146 14044 4558
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 13832 3058 13860 3538
rect 13910 3496 13966 3505
rect 13910 3431 13966 3440
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 13832 2582 13860 2994
rect 13924 2922 13952 3431
rect 14016 3194 14044 4082
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14384 3505 14412 3538
rect 14370 3496 14426 3505
rect 14370 3431 14426 3440
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14289 2672 14585 2692
rect 14752 2650 14780 5170
rect 14832 5092 14884 5098
rect 14832 5034 14884 5040
rect 14844 4826 14872 5034
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14936 4758 14964 5188
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 14832 3664 14884 3670
rect 14832 3606 14884 3612
rect 14844 2922 14872 3606
rect 15120 3126 15148 4014
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15212 3398 15240 3878
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 15108 3120 15160 3126
rect 15108 3062 15160 3068
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 14830 2680 14886 2689
rect 14740 2644 14792 2650
rect 14830 2615 14886 2624
rect 14740 2586 14792 2592
rect 13820 2576 13872 2582
rect 12346 2544 12402 2553
rect 13820 2518 13872 2524
rect 14844 2514 14872 2615
rect 12346 2479 12402 2488
rect 13360 2508 13412 2514
rect 12360 2310 12388 2479
rect 13360 2450 13412 2456
rect 14832 2508 14884 2514
rect 14832 2450 14884 2456
rect 13372 2310 13400 2450
rect 12348 2304 12400 2310
rect 11978 2272 12034 2281
rect 12348 2246 12400 2252
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 11978 2207 12034 2216
rect 13372 2009 13400 2246
rect 13358 2000 13414 2009
rect 13358 1935 13414 1944
rect 13372 1329 13400 1935
rect 13358 1320 13414 1329
rect 13358 1255 13414 1264
rect 11610 54 11744 82
rect 14936 82 14964 2926
rect 15120 2650 15148 3062
rect 15212 3058 15240 3334
rect 15672 3194 15700 11630
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15764 9042 15792 11290
rect 15948 10062 15976 11494
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16500 10810 16528 11154
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15948 9654 15976 9998
rect 16040 9722 16068 10134
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 15936 9648 15988 9654
rect 15936 9590 15988 9596
rect 15844 9444 15896 9450
rect 15844 9386 15896 9392
rect 15856 9110 15884 9386
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 15764 8634 15792 8978
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15752 8288 15804 8294
rect 15856 8276 15884 9046
rect 16132 8498 16160 9862
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 15804 8248 15884 8276
rect 15752 8230 15804 8236
rect 15764 8022 15792 8230
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15764 7342 15792 7958
rect 16120 7472 16172 7478
rect 16120 7414 16172 7420
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 16132 6798 16160 7414
rect 16212 7268 16264 7274
rect 16212 7210 16264 7216
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16040 6390 16068 6734
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 16132 5710 16160 6734
rect 16224 6118 16252 7210
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 16316 6458 16344 6870
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16224 5166 16252 6054
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15764 4146 15792 4966
rect 15936 4752 15988 4758
rect 15936 4694 15988 4700
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15948 3738 15976 4694
rect 16224 4554 16252 5102
rect 16316 5030 16344 5510
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16592 4622 16620 11494
rect 17144 10810 17172 15558
rect 17498 15520 17554 15558
rect 22112 15558 22522 15586
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16684 9178 16712 9658
rect 17500 9512 17552 9518
rect 17498 9480 17500 9489
rect 17552 9480 17554 9489
rect 17498 9415 17554 9424
rect 17512 9382 17540 9415
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 17328 8498 17356 9318
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16868 7750 16896 8366
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 17052 8090 17080 8298
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 17052 7410 17080 8026
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16684 6934 16712 7210
rect 16672 6928 16724 6934
rect 16672 6870 16724 6876
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16684 4690 16712 5510
rect 16764 4752 16816 4758
rect 16764 4694 16816 4700
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16580 4616 16632 4622
rect 16394 4584 16450 4593
rect 16212 4548 16264 4554
rect 16580 4558 16632 4564
rect 16488 4548 16540 4554
rect 16450 4528 16488 4536
rect 16394 4519 16488 4528
rect 16408 4508 16488 4519
rect 16212 4490 16264 4496
rect 16488 4490 16540 4496
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16316 4282 16344 4422
rect 16304 4276 16356 4282
rect 16304 4218 16356 4224
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 16224 3466 16252 4082
rect 16408 3602 16436 4218
rect 16684 4010 16712 4626
rect 16776 4146 16804 4694
rect 16868 4214 16896 6258
rect 16960 5846 16988 6598
rect 17144 6322 17172 8434
rect 17604 8022 17632 10950
rect 18156 10130 18184 12038
rect 19168 11558 19196 12242
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 22112 11898 22140 15558
rect 22466 15520 22522 15558
rect 27080 15558 27490 15586
rect 24124 12708 24176 12714
rect 24124 12650 24176 12656
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 19616 11824 19668 11830
rect 19616 11766 19668 11772
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19628 11218 19656 11766
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 18340 10810 18368 11154
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 19168 10742 19196 11154
rect 19156 10736 19208 10742
rect 19156 10678 19208 10684
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 19168 10266 19196 10474
rect 19536 10282 19564 10610
rect 19628 10452 19656 11154
rect 19720 10674 19748 11494
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 19708 10464 19760 10470
rect 19628 10424 19708 10452
rect 19708 10406 19760 10412
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 19248 10260 19300 10266
rect 19536 10254 19656 10282
rect 19248 10202 19300 10208
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 17696 9178 17724 10066
rect 18156 9722 18184 10066
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18786 10024 18842 10033
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17592 8016 17644 8022
rect 17592 7958 17644 7964
rect 17604 7002 17632 7958
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17604 6390 17632 6802
rect 17592 6384 17644 6390
rect 17592 6326 17644 6332
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17696 6254 17724 9114
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17972 8537 18000 8978
rect 17958 8528 18014 8537
rect 17958 8463 18014 8472
rect 17972 8430 18000 8463
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17868 8288 17920 8294
rect 17972 8265 18000 8366
rect 17868 8230 17920 8236
rect 17958 8256 18014 8265
rect 17880 8022 17908 8230
rect 17958 8191 18014 8200
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17880 7818 17908 7958
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 17880 7546 17908 7754
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 17788 6458 17816 6802
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16960 5234 16988 5782
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 17696 4690 17724 6190
rect 17788 5574 17816 6394
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17788 5370 17816 5510
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 18156 5166 18184 9658
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18248 8022 18276 8774
rect 18236 8016 18288 8022
rect 18236 7958 18288 7964
rect 18236 6384 18288 6390
rect 18236 6326 18288 6332
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 17774 4856 17830 4865
rect 17774 4791 17830 4800
rect 18144 4820 18196 4826
rect 17684 4684 17736 4690
rect 17604 4644 17684 4672
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 16960 4214 16988 4558
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 16856 4208 16908 4214
rect 16856 4150 16908 4156
rect 16948 4208 17000 4214
rect 16948 4150 17000 4156
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16776 3942 16804 4082
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 16224 3126 16252 3402
rect 16212 3120 16264 3126
rect 16212 3062 16264 3068
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 16408 2990 16436 3538
rect 16776 3058 16804 3878
rect 17144 3097 17172 4422
rect 17604 3738 17632 4644
rect 17684 4626 17736 4632
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17788 3670 17816 4791
rect 18144 4762 18196 4768
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 17788 3194 17816 3606
rect 17972 3534 18000 4014
rect 18064 3942 18092 4150
rect 18156 4078 18184 4762
rect 18248 4604 18276 6326
rect 18340 5778 18368 9998
rect 18786 9959 18842 9968
rect 18800 9722 18828 9959
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18800 9518 18828 9658
rect 19168 9586 19196 10202
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18616 9178 18644 9318
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18432 8362 18460 8774
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18420 8356 18472 8362
rect 18420 8298 18472 8304
rect 18524 8090 18552 8434
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18616 7886 18644 8434
rect 19076 8294 19104 9046
rect 19260 8634 19288 10202
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19536 9382 19564 10066
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 19076 8090 19104 8230
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 19260 8022 19288 8298
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 18604 7880 18656 7886
rect 18656 7840 18736 7868
rect 18604 7822 18656 7828
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18524 6322 18552 6938
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18616 6186 18644 7142
rect 18708 6866 18736 7840
rect 19260 7546 19288 7958
rect 19536 7886 19564 8842
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19536 7410 19564 7822
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19432 7268 19484 7274
rect 19432 7210 19484 7216
rect 19444 7002 19472 7210
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19340 6928 19392 6934
rect 19340 6870 19392 6876
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18708 6322 18736 6802
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18604 6180 18656 6186
rect 18604 6122 18656 6128
rect 18616 5914 18644 6122
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18696 5908 18748 5914
rect 18696 5850 18748 5856
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18340 4826 18368 5714
rect 18512 5092 18564 5098
rect 18512 5034 18564 5040
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18328 4616 18380 4622
rect 18248 4576 18328 4604
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17972 3126 18000 3470
rect 18052 3460 18104 3466
rect 18052 3402 18104 3408
rect 17960 3120 18012 3126
rect 17130 3088 17186 3097
rect 16764 3052 16816 3058
rect 17960 3062 18012 3068
rect 17130 3023 17186 3032
rect 16764 2994 16816 3000
rect 16396 2984 16448 2990
rect 16396 2926 16448 2932
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 16408 2650 16436 2926
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 16684 2514 16712 2926
rect 16776 2650 16804 2994
rect 18064 2650 18092 3402
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 15212 2310 15240 2450
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15014 82 15070 480
rect 15212 377 15240 2246
rect 15198 368 15254 377
rect 15198 303 15254 312
rect 14936 54 15070 82
rect 18156 82 18184 4014
rect 18248 3194 18276 4576
rect 18328 4558 18380 4564
rect 18420 4208 18472 4214
rect 18420 4150 18472 4156
rect 18432 4078 18460 4150
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18432 3534 18460 4014
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18328 3460 18380 3466
rect 18328 3402 18380 3408
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18340 2990 18368 3402
rect 18432 3058 18460 3470
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18524 2689 18552 5034
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 18510 2680 18566 2689
rect 18616 2650 18644 4626
rect 18708 3670 18736 5850
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18800 4690 18828 5170
rect 18892 4690 18920 6734
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18984 4758 19012 6598
rect 19352 6186 19380 6870
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 19352 5846 19380 6122
rect 19340 5840 19392 5846
rect 19340 5782 19392 5788
rect 19352 5370 19380 5782
rect 19628 5642 19656 10254
rect 19720 10130 19748 10406
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19720 9110 19748 10066
rect 19904 9586 19932 11086
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 20088 10266 20116 10610
rect 20180 10538 20208 10950
rect 20168 10532 20220 10538
rect 20168 10474 20220 10480
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20180 9722 20208 10474
rect 20640 10470 20668 11222
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 21272 10736 21324 10742
rect 21376 10713 21404 11630
rect 22008 11620 22060 11626
rect 22008 11562 22060 11568
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 21652 11150 21680 11494
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21640 11144 21692 11150
rect 21640 11086 21692 11092
rect 21468 10810 21496 11086
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21272 10678 21324 10684
rect 21362 10704 21418 10713
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19708 9104 19760 9110
rect 19708 9046 19760 9052
rect 20640 8634 20668 10406
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20732 9178 20760 9998
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 20810 9616 20866 9625
rect 20810 9551 20866 9560
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20824 9042 20852 9551
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 20548 7750 20576 8298
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 19616 5636 19668 5642
rect 19616 5578 19668 5584
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19628 5166 19656 5578
rect 20180 5574 20208 6190
rect 20168 5568 20220 5574
rect 20168 5510 20220 5516
rect 20180 5234 20208 5510
rect 20548 5370 20576 7686
rect 20732 7546 20760 8774
rect 20824 8634 20852 8978
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 21284 8634 21312 10678
rect 21652 10674 21680 11086
rect 21362 10639 21418 10648
rect 21640 10668 21692 10674
rect 21640 10610 21692 10616
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21364 9444 21416 9450
rect 21364 9386 21416 9392
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21284 8430 21312 8570
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 21376 8294 21404 9386
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20626 7440 20682 7449
rect 20626 7375 20682 7384
rect 20640 7342 20668 7375
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 21376 7274 21404 8230
rect 21364 7268 21416 7274
rect 21364 7210 21416 7216
rect 21272 6928 21324 6934
rect 21272 6870 21324 6876
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 21284 6458 21312 6870
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21376 6186 21404 7210
rect 21364 6180 21416 6186
rect 21364 6122 21416 6128
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20640 5846 20668 6054
rect 21468 5914 21496 10542
rect 21652 10130 21680 10610
rect 21732 10464 21784 10470
rect 21732 10406 21784 10412
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21744 9761 21772 10406
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 21730 9752 21786 9761
rect 21928 9722 21956 10134
rect 21730 9687 21786 9696
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 22020 9625 22048 11562
rect 23112 11212 23164 11218
rect 23112 11154 23164 11160
rect 23020 11008 23072 11014
rect 23020 10950 23072 10956
rect 22834 10704 22890 10713
rect 22834 10639 22890 10648
rect 22848 10606 22876 10639
rect 22836 10600 22888 10606
rect 22836 10542 22888 10548
rect 22006 9616 22062 9625
rect 21824 9580 21876 9586
rect 22006 9551 22062 9560
rect 21824 9522 21876 9528
rect 21732 9376 21784 9382
rect 21732 9318 21784 9324
rect 21548 8832 21600 8838
rect 21548 8774 21600 8780
rect 21560 8430 21588 8774
rect 21548 8424 21600 8430
rect 21548 8366 21600 8372
rect 21548 8288 21600 8294
rect 21548 8230 21600 8236
rect 21560 7410 21588 8230
rect 21640 8016 21692 8022
rect 21640 7958 21692 7964
rect 21652 7546 21680 7958
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 21560 7002 21588 7346
rect 21652 7002 21680 7482
rect 21548 6996 21600 7002
rect 21548 6938 21600 6944
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20168 5228 20220 5234
rect 20168 5170 20220 5176
rect 20548 5166 20576 5306
rect 19248 5160 19300 5166
rect 19248 5102 19300 5108
rect 19616 5160 19668 5166
rect 19616 5102 19668 5108
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18788 3936 18840 3942
rect 19156 3936 19208 3942
rect 18788 3878 18840 3884
rect 18970 3904 19026 3913
rect 18696 3664 18748 3670
rect 18696 3606 18748 3612
rect 18800 3097 18828 3878
rect 19156 3878 19208 3884
rect 18970 3839 19026 3848
rect 18880 3664 18932 3670
rect 18880 3606 18932 3612
rect 18786 3088 18842 3097
rect 18786 3023 18842 3032
rect 18510 2615 18566 2624
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 18892 2582 18920 3606
rect 18880 2576 18932 2582
rect 18880 2518 18932 2524
rect 18984 2446 19012 3839
rect 19168 2650 19196 3878
rect 19260 3602 19288 5102
rect 19708 5092 19760 5098
rect 19708 5034 19760 5040
rect 19432 4208 19484 4214
rect 19432 4150 19484 4156
rect 19444 4010 19472 4150
rect 19432 4004 19484 4010
rect 19432 3946 19484 3952
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19260 3505 19288 3538
rect 19246 3496 19302 3505
rect 19246 3431 19302 3440
rect 19260 2854 19288 3431
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19444 2922 19472 2994
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 19260 2310 19288 2790
rect 19720 2582 19748 5034
rect 20640 4826 20668 5782
rect 20812 5704 20864 5710
rect 20812 5646 20864 5652
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20732 5166 20760 5510
rect 20824 5370 20852 5646
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 20824 4826 20852 5306
rect 21456 5160 21508 5166
rect 21456 5102 21508 5108
rect 21638 5128 21694 5137
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 20812 4820 20864 4826
rect 20812 4762 20864 4768
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19904 4282 19932 4422
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 19892 4276 19944 4282
rect 19892 4218 19944 4224
rect 21180 4140 21232 4146
rect 21180 4082 21232 4088
rect 20628 4004 20680 4010
rect 20628 3946 20680 3952
rect 20640 3738 20668 3946
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20260 3664 20312 3670
rect 20260 3606 20312 3612
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19904 2961 19932 3470
rect 19890 2952 19946 2961
rect 20272 2922 20300 3606
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 19890 2887 19946 2896
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 20260 2916 20312 2922
rect 20260 2858 20312 2864
rect 19996 2582 20024 2858
rect 20640 2854 20668 3470
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 19708 2576 19760 2582
rect 19708 2518 19760 2524
rect 19984 2576 20036 2582
rect 19984 2518 20036 2524
rect 19248 2304 19300 2310
rect 20640 2281 20668 2790
rect 20824 2553 20852 3878
rect 21192 3602 21220 4082
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 20904 2916 20956 2922
rect 20904 2858 20956 2864
rect 20916 2825 20944 2858
rect 21468 2854 21496 5102
rect 21638 5063 21694 5072
rect 21652 4185 21680 5063
rect 21744 4758 21772 9318
rect 21836 9178 21864 9522
rect 21824 9172 21876 9178
rect 21824 9114 21876 9120
rect 22468 9036 22520 9042
rect 22468 8978 22520 8984
rect 22480 8294 22508 8978
rect 22468 8288 22520 8294
rect 22468 8230 22520 8236
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 21836 6866 21864 7822
rect 22480 7313 22508 8230
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 22466 7304 22522 7313
rect 22466 7239 22522 7248
rect 22664 7206 22692 7890
rect 22848 7342 22876 10542
rect 23032 10062 23060 10950
rect 23124 10470 23152 11154
rect 24136 10849 24164 12650
rect 24584 12640 24636 12646
rect 24584 12582 24636 12588
rect 24216 12300 24268 12306
rect 24216 12242 24268 12248
rect 24228 11801 24256 12242
rect 24400 12096 24452 12102
rect 24400 12038 24452 12044
rect 24214 11792 24270 11801
rect 24214 11727 24216 11736
rect 24268 11727 24270 11736
rect 24216 11698 24268 11704
rect 24228 11667 24256 11698
rect 24412 11286 24440 12038
rect 24400 11280 24452 11286
rect 24400 11222 24452 11228
rect 24492 11280 24544 11286
rect 24492 11222 24544 11228
rect 24122 10840 24178 10849
rect 23480 10804 23532 10810
rect 24412 10810 24440 11222
rect 24122 10775 24178 10784
rect 24400 10804 24452 10810
rect 23480 10746 23532 10752
rect 23296 10532 23348 10538
rect 23296 10474 23348 10480
rect 23112 10464 23164 10470
rect 23112 10406 23164 10412
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 23032 9722 23060 9998
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 23124 9602 23152 10406
rect 23204 10192 23256 10198
rect 23204 10134 23256 10140
rect 23216 9722 23244 10134
rect 23204 9716 23256 9722
rect 23204 9658 23256 9664
rect 23308 9654 23336 10474
rect 23492 10062 23520 10746
rect 23480 10056 23532 10062
rect 24136 10033 24164 10775
rect 24400 10746 24452 10752
rect 24400 10464 24452 10470
rect 24504 10452 24532 11222
rect 24596 10674 24624 12582
rect 25320 12300 25372 12306
rect 25320 12242 25372 12248
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24676 11552 24728 11558
rect 24676 11494 24728 11500
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24584 10532 24636 10538
rect 24584 10474 24636 10480
rect 24452 10424 24532 10452
rect 24400 10406 24452 10412
rect 23480 9998 23532 10004
rect 24122 10024 24178 10033
rect 24122 9959 24178 9968
rect 24412 9926 24440 10406
rect 24596 10198 24624 10474
rect 24584 10192 24636 10198
rect 24584 10134 24636 10140
rect 23664 9920 23716 9926
rect 23664 9862 23716 9868
rect 24400 9920 24452 9926
rect 24400 9862 24452 9868
rect 23296 9648 23348 9654
rect 23124 9574 23244 9602
rect 23296 9590 23348 9596
rect 23676 9586 23704 9862
rect 23020 9512 23072 9518
rect 23020 9454 23072 9460
rect 23032 9110 23060 9454
rect 23020 9104 23072 9110
rect 23020 9046 23072 9052
rect 22928 9036 22980 9042
rect 22928 8978 22980 8984
rect 22940 8294 22968 8978
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 22940 8090 22968 8230
rect 22928 8084 22980 8090
rect 22928 8026 22980 8032
rect 23112 7948 23164 7954
rect 23032 7908 23112 7936
rect 22836 7336 22888 7342
rect 22836 7278 22888 7284
rect 23032 7206 23060 7908
rect 23112 7890 23164 7896
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 22652 7200 22704 7206
rect 22652 7142 22704 7148
rect 23020 7200 23072 7206
rect 23020 7142 23072 7148
rect 21824 6860 21876 6866
rect 21824 6802 21876 6808
rect 21732 4752 21784 4758
rect 21732 4694 21784 4700
rect 21638 4176 21694 4185
rect 21638 4111 21694 4120
rect 21456 2848 21508 2854
rect 20902 2816 20958 2825
rect 21456 2790 21508 2796
rect 20902 2751 20958 2760
rect 20916 2650 20944 2751
rect 21652 2650 21680 4111
rect 21916 4072 21968 4078
rect 22020 4060 22048 7142
rect 22468 6860 22520 6866
rect 22468 6802 22520 6808
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22112 5574 22140 6190
rect 22284 6112 22336 6118
rect 22284 6054 22336 6060
rect 22296 5710 22324 6054
rect 22480 5914 22508 6802
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 22112 5098 22140 5510
rect 22296 5370 22324 5646
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22100 5092 22152 5098
rect 22100 5034 22152 5040
rect 23032 4865 23060 7142
rect 23112 6860 23164 6866
rect 23112 6802 23164 6808
rect 23124 6458 23152 6802
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23124 5642 23152 6394
rect 23112 5636 23164 5642
rect 23112 5578 23164 5584
rect 23018 4856 23074 4865
rect 23018 4791 23074 4800
rect 22192 4684 22244 4690
rect 22192 4626 22244 4632
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 22204 4146 22232 4626
rect 22376 4616 22428 4622
rect 22376 4558 22428 4564
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 22388 4078 22416 4558
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 21968 4032 22048 4060
rect 21916 4014 21968 4020
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 21836 3058 21864 3470
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 21916 2848 21968 2854
rect 22020 2836 22048 4032
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 22376 4072 22428 4078
rect 22376 4014 22428 4020
rect 22112 3670 22140 4014
rect 22664 3738 22692 4082
rect 22940 4010 22968 4626
rect 23216 4154 23244 9574
rect 23664 9580 23716 9586
rect 23664 9522 23716 9528
rect 23664 9444 23716 9450
rect 23664 9386 23716 9392
rect 23676 9110 23704 9386
rect 23664 9104 23716 9110
rect 23664 9046 23716 9052
rect 23676 8838 23704 9046
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23676 8294 23704 8774
rect 24412 8634 24440 9862
rect 24596 9722 24624 10134
rect 24584 9716 24636 9722
rect 24584 9658 24636 9664
rect 24688 9586 24716 11494
rect 24780 10198 24808 12038
rect 25332 11694 25360 12242
rect 25320 11688 25372 11694
rect 25320 11630 25372 11636
rect 25228 11144 25280 11150
rect 25228 11086 25280 11092
rect 25240 10538 25268 11086
rect 25228 10532 25280 10538
rect 25228 10474 25280 10480
rect 25240 10266 25268 10474
rect 25228 10260 25280 10266
rect 25228 10202 25280 10208
rect 24768 10192 24820 10198
rect 24768 10134 24820 10140
rect 24860 10192 24912 10198
rect 24860 10134 24912 10140
rect 24676 9580 24728 9586
rect 24676 9522 24728 9528
rect 24780 9178 24808 10134
rect 24872 9722 24900 10134
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24872 9382 24900 9658
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 24872 9042 24900 9318
rect 25136 9172 25188 9178
rect 25136 9114 25188 9120
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 25148 8974 25176 9114
rect 25136 8968 25188 8974
rect 25136 8910 25188 8916
rect 25148 8634 25176 8910
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 24216 8424 24268 8430
rect 24216 8366 24268 8372
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23664 8288 23716 8294
rect 23664 8230 23716 8236
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23492 6322 23520 7482
rect 23768 6390 23796 8298
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 24136 7342 24164 7890
rect 24228 7750 24256 8366
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 25136 8288 25188 8294
rect 25332 8265 25360 11630
rect 25412 11552 25464 11558
rect 25412 11494 25464 11500
rect 25424 8634 25452 11494
rect 27080 11354 27108 15558
rect 27434 15520 27490 15558
rect 31208 15564 31260 15570
rect 32494 15564 32550 16000
rect 37462 15586 37518 16000
rect 32494 15520 32496 15564
rect 31208 15506 31260 15512
rect 32548 15520 32550 15564
rect 37200 15558 37518 15586
rect 32496 15506 32548 15512
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 29552 12232 29604 12238
rect 29552 12174 29604 12180
rect 28448 11756 28500 11762
rect 28448 11698 28500 11704
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 27068 11348 27120 11354
rect 27068 11290 27120 11296
rect 27068 11212 27120 11218
rect 27068 11154 27120 11160
rect 27528 11212 27580 11218
rect 27528 11154 27580 11160
rect 28080 11212 28132 11218
rect 28080 11154 28132 11160
rect 27080 10810 27108 11154
rect 27068 10804 27120 10810
rect 26988 10764 27068 10792
rect 26240 10600 26292 10606
rect 26240 10542 26292 10548
rect 26148 10464 26200 10470
rect 26148 10406 26200 10412
rect 25964 10192 26016 10198
rect 25964 10134 26016 10140
rect 25780 9988 25832 9994
rect 25780 9930 25832 9936
rect 25792 9586 25820 9930
rect 25976 9926 26004 10134
rect 25964 9920 26016 9926
rect 25964 9862 26016 9868
rect 25976 9722 26004 9862
rect 25964 9716 26016 9722
rect 25964 9658 26016 9664
rect 25504 9580 25556 9586
rect 25504 9522 25556 9528
rect 25780 9580 25832 9586
rect 25780 9522 25832 9528
rect 25516 9110 25544 9522
rect 25504 9104 25556 9110
rect 25504 9046 25556 9052
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25872 8356 25924 8362
rect 25872 8298 25924 8304
rect 25136 8230 25188 8236
rect 25318 8256 25374 8265
rect 24688 8022 24716 8230
rect 24676 8016 24728 8022
rect 24676 7958 24728 7964
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 24216 7744 24268 7750
rect 24216 7686 24268 7692
rect 24228 7410 24256 7686
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24124 7336 24176 7342
rect 24124 7278 24176 7284
rect 24412 6866 24440 7822
rect 24688 7206 24716 7958
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 25056 7206 25084 7822
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 24400 6860 24452 6866
rect 24400 6802 24452 6808
rect 23756 6384 23808 6390
rect 23756 6326 23808 6332
rect 23480 6316 23532 6322
rect 23480 6258 23532 6264
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 23572 6112 23624 6118
rect 23572 6054 23624 6060
rect 23584 5914 23612 6054
rect 23676 5914 23704 6190
rect 23572 5908 23624 5914
rect 23572 5850 23624 5856
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 23584 5030 23612 5850
rect 23676 5030 23704 5850
rect 23768 5166 23796 6326
rect 24688 6186 24716 7142
rect 25056 6934 25084 7142
rect 25044 6928 25096 6934
rect 25044 6870 25096 6876
rect 24952 6724 25004 6730
rect 24952 6666 25004 6672
rect 24964 6458 24992 6666
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 25042 6352 25098 6361
rect 25148 6338 25176 8230
rect 25318 8191 25374 8200
rect 25884 8090 25912 8298
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 25688 7812 25740 7818
rect 25688 7754 25740 7760
rect 25320 6860 25372 6866
rect 25320 6802 25372 6808
rect 25332 6458 25360 6802
rect 25412 6656 25464 6662
rect 25412 6598 25464 6604
rect 25320 6452 25372 6458
rect 25320 6394 25372 6400
rect 25098 6310 25176 6338
rect 25042 6287 25098 6296
rect 24676 6180 24728 6186
rect 24676 6122 24728 6128
rect 24584 6112 24636 6118
rect 24584 6054 24636 6060
rect 24596 5846 24624 6054
rect 24584 5840 24636 5846
rect 24584 5782 24636 5788
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24124 5568 24176 5574
rect 24124 5510 24176 5516
rect 24136 5370 24164 5510
rect 24124 5364 24176 5370
rect 24124 5306 24176 5312
rect 23756 5160 23808 5166
rect 23756 5102 23808 5108
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 23664 5024 23716 5030
rect 23664 4966 23716 4972
rect 23478 4720 23534 4729
rect 23478 4655 23534 4664
rect 23388 4616 23440 4622
rect 23388 4558 23440 4564
rect 23216 4126 23336 4154
rect 23400 4146 23428 4558
rect 22928 4004 22980 4010
rect 22928 3946 22980 3952
rect 22744 3936 22796 3942
rect 22744 3878 22796 3884
rect 22652 3732 22704 3738
rect 22652 3674 22704 3680
rect 22100 3664 22152 3670
rect 22100 3606 22152 3612
rect 22112 3466 22140 3606
rect 22560 3596 22612 3602
rect 22560 3538 22612 3544
rect 22100 3460 22152 3466
rect 22100 3402 22152 3408
rect 22112 3058 22140 3402
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 22572 2854 22600 3538
rect 22756 2990 22784 3878
rect 23308 3369 23336 4126
rect 23388 4140 23440 4146
rect 23388 4082 23440 4088
rect 23294 3360 23350 3369
rect 23294 3295 23350 3304
rect 23492 3126 23520 4655
rect 23584 3992 23612 4966
rect 23768 4826 23796 5102
rect 24032 5092 24084 5098
rect 24032 5034 24084 5040
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 24044 4282 24072 5034
rect 24688 5030 24716 5714
rect 25056 5302 25084 6287
rect 25136 5772 25188 5778
rect 25136 5714 25188 5720
rect 25044 5296 25096 5302
rect 25044 5238 25096 5244
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24688 4865 24716 4966
rect 24674 4856 24730 4865
rect 24674 4791 24730 4800
rect 24952 4684 25004 4690
rect 24952 4626 25004 4632
rect 24492 4480 24544 4486
rect 24492 4422 24544 4428
rect 24032 4276 24084 4282
rect 24032 4218 24084 4224
rect 24124 4208 24176 4214
rect 24124 4150 24176 4156
rect 23756 4004 23808 4010
rect 23584 3964 23756 3992
rect 23756 3946 23808 3952
rect 23664 3596 23716 3602
rect 23664 3538 23716 3544
rect 23676 3194 23704 3538
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 23480 3120 23532 3126
rect 23480 3062 23532 3068
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 23768 2904 23796 3946
rect 24136 3913 24164 4150
rect 24504 4078 24532 4422
rect 24964 4154 24992 4626
rect 25148 4622 25176 5714
rect 25320 5092 25372 5098
rect 25320 5034 25372 5040
rect 25332 4690 25360 5034
rect 25320 4684 25372 4690
rect 25320 4626 25372 4632
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 24964 4146 25084 4154
rect 24964 4140 25096 4146
rect 24964 4126 25044 4140
rect 25044 4082 25096 4088
rect 24492 4072 24544 4078
rect 24492 4014 24544 4020
rect 24122 3904 24178 3913
rect 24122 3839 24178 3848
rect 24504 3738 24532 4014
rect 24952 4004 25004 4010
rect 24952 3946 25004 3952
rect 24492 3732 24544 3738
rect 24492 3674 24544 3680
rect 24964 3670 24992 3946
rect 24952 3664 25004 3670
rect 24952 3606 25004 3612
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24596 3058 24624 3334
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 23985 2916 24037 2922
rect 23768 2876 23985 2904
rect 22100 2848 22152 2854
rect 22020 2808 22100 2836
rect 21916 2790 21968 2796
rect 22100 2790 22152 2796
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 23572 2848 23624 2854
rect 23768 2825 23796 2876
rect 23985 2858 24037 2864
rect 24872 2854 24900 3538
rect 25228 3392 25280 3398
rect 25228 3334 25280 3340
rect 24860 2848 24912 2854
rect 23572 2790 23624 2796
rect 23754 2816 23810 2825
rect 21928 2650 21956 2790
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 21640 2644 21692 2650
rect 21640 2586 21692 2592
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 22112 2553 22140 2790
rect 23584 2582 23612 2790
rect 24860 2790 24912 2796
rect 23754 2751 23810 2760
rect 23768 2650 23796 2751
rect 24674 2680 24730 2689
rect 23756 2644 23808 2650
rect 25240 2650 25268 3334
rect 24674 2615 24730 2624
rect 25228 2644 25280 2650
rect 23756 2586 23808 2592
rect 23572 2576 23624 2582
rect 20810 2544 20866 2553
rect 20810 2479 20866 2488
rect 22098 2544 22154 2553
rect 23572 2518 23624 2524
rect 24492 2576 24544 2582
rect 24492 2518 24544 2524
rect 22098 2479 22154 2488
rect 24032 2508 24084 2514
rect 24032 2450 24084 2456
rect 24044 2417 24072 2450
rect 24030 2408 24086 2417
rect 24030 2343 24086 2352
rect 24504 2310 24532 2518
rect 21456 2304 21508 2310
rect 19248 2246 19300 2252
rect 20626 2272 20682 2281
rect 21456 2246 21508 2252
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 20626 2207 20682 2216
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 18326 82 18382 480
rect 18156 54 18382 82
rect 21468 82 21496 2246
rect 21638 82 21694 480
rect 21468 54 21694 82
rect 24688 82 24716 2615
rect 25228 2586 25280 2592
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 24872 2417 24900 2450
rect 24858 2408 24914 2417
rect 24858 2343 24914 2352
rect 24950 82 25006 480
rect 25424 134 25452 6598
rect 25504 5704 25556 5710
rect 25504 5646 25556 5652
rect 25516 3942 25544 5646
rect 25700 4146 25728 7754
rect 26160 7410 26188 10406
rect 26252 10130 26280 10542
rect 26240 10124 26292 10130
rect 26240 10066 26292 10072
rect 26148 7404 26200 7410
rect 26148 7346 26200 7352
rect 26160 7002 26188 7346
rect 26148 6996 26200 7002
rect 26148 6938 26200 6944
rect 26252 6730 26280 10066
rect 26332 10056 26384 10062
rect 26332 9998 26384 10004
rect 26344 9654 26372 9998
rect 26332 9648 26384 9654
rect 26332 9590 26384 9596
rect 26344 9110 26372 9590
rect 26332 9104 26384 9110
rect 26332 9046 26384 9052
rect 26516 9036 26568 9042
rect 26516 8978 26568 8984
rect 26528 8294 26556 8978
rect 26988 8498 27016 10764
rect 27068 10746 27120 10752
rect 27540 10470 27568 11154
rect 28092 11014 28120 11154
rect 28080 11008 28132 11014
rect 28080 10950 28132 10956
rect 28092 10606 28120 10950
rect 28080 10600 28132 10606
rect 28080 10542 28132 10548
rect 27528 10464 27580 10470
rect 27528 10406 27580 10412
rect 27068 9920 27120 9926
rect 27068 9862 27120 9868
rect 27080 9761 27108 9862
rect 27066 9752 27122 9761
rect 27066 9687 27122 9696
rect 27080 9654 27108 9687
rect 27068 9648 27120 9654
rect 27068 9590 27120 9596
rect 27068 9036 27120 9042
rect 27068 8978 27120 8984
rect 27080 8634 27108 8978
rect 27068 8628 27120 8634
rect 27068 8570 27120 8576
rect 26976 8492 27028 8498
rect 26976 8434 27028 8440
rect 26516 8288 26568 8294
rect 26516 8230 26568 8236
rect 26790 8256 26846 8265
rect 26790 8191 26846 8200
rect 26700 7880 26752 7886
rect 26700 7822 26752 7828
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 26240 6724 26292 6730
rect 26240 6666 26292 6672
rect 25872 6248 25924 6254
rect 25872 6190 25924 6196
rect 25884 5574 25912 6190
rect 25872 5568 25924 5574
rect 25872 5510 25924 5516
rect 25884 5234 25912 5510
rect 26252 5302 26280 6666
rect 26344 5914 26372 6734
rect 26712 6662 26740 7822
rect 26804 7449 26832 8191
rect 26988 7478 27016 8434
rect 27080 7954 27108 8570
rect 27540 8430 27568 10406
rect 27622 10364 27918 10384
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 28092 9926 28120 10542
rect 28356 10532 28408 10538
rect 28356 10474 28408 10480
rect 28080 9920 28132 9926
rect 28080 9862 28132 9868
rect 28092 9518 28120 9862
rect 28080 9512 28132 9518
rect 28080 9454 28132 9460
rect 28264 9444 28316 9450
rect 28264 9386 28316 9392
rect 27622 9276 27918 9296
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 27622 9200 27918 9220
rect 27712 8832 27764 8838
rect 27712 8774 27764 8780
rect 27724 8430 27752 8774
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27712 8424 27764 8430
rect 27712 8366 27764 8372
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27622 8112 27918 8132
rect 27344 8016 27396 8022
rect 27344 7958 27396 7964
rect 27068 7948 27120 7954
rect 27068 7890 27120 7896
rect 26976 7472 27028 7478
rect 26790 7440 26846 7449
rect 26976 7414 27028 7420
rect 26790 7375 26846 7384
rect 27356 7274 27384 7958
rect 27436 7744 27488 7750
rect 27436 7686 27488 7692
rect 27712 7744 27764 7750
rect 27712 7686 27764 7692
rect 27344 7268 27396 7274
rect 27344 7210 27396 7216
rect 27448 6934 27476 7686
rect 27528 7472 27580 7478
rect 27528 7414 27580 7420
rect 27436 6928 27488 6934
rect 27436 6870 27488 6876
rect 26700 6656 26752 6662
rect 26700 6598 26752 6604
rect 26332 5908 26384 5914
rect 26332 5850 26384 5856
rect 26240 5296 26292 5302
rect 26240 5238 26292 5244
rect 25872 5228 25924 5234
rect 25872 5170 25924 5176
rect 26712 4758 26740 6598
rect 27448 6458 27476 6870
rect 27540 6798 27568 7414
rect 27724 7410 27752 7686
rect 27712 7404 27764 7410
rect 27712 7346 27764 7352
rect 27988 7404 28040 7410
rect 27988 7346 28040 7352
rect 27622 7100 27918 7120
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 27528 6792 27580 6798
rect 27528 6734 27580 6740
rect 27436 6452 27488 6458
rect 27436 6394 27488 6400
rect 28000 6322 28028 7346
rect 28276 7002 28304 9386
rect 28368 9042 28396 10474
rect 28460 9058 28488 11698
rect 29564 11286 29592 12174
rect 29828 11824 29880 11830
rect 29828 11766 29880 11772
rect 29552 11280 29604 11286
rect 29552 11222 29604 11228
rect 29564 10810 29592 11222
rect 29644 11144 29696 11150
rect 29644 11086 29696 11092
rect 29552 10804 29604 10810
rect 29552 10746 29604 10752
rect 29460 10736 29512 10742
rect 29460 10678 29512 10684
rect 29472 10266 29500 10678
rect 29656 10266 29684 11086
rect 29460 10260 29512 10266
rect 29460 10202 29512 10208
rect 29644 10260 29696 10266
rect 29644 10202 29696 10208
rect 28632 10192 28684 10198
rect 28632 10134 28684 10140
rect 28540 10056 28592 10062
rect 28540 9998 28592 10004
rect 28552 9586 28580 9998
rect 28540 9580 28592 9586
rect 28540 9522 28592 9528
rect 28552 9178 28580 9522
rect 28644 9382 28672 10134
rect 29656 9586 29684 10202
rect 29840 9761 29868 11766
rect 30288 11552 30340 11558
rect 30288 11494 30340 11500
rect 29920 11280 29972 11286
rect 29920 11222 29972 11228
rect 29932 10742 29960 11222
rect 29920 10736 29972 10742
rect 29920 10678 29972 10684
rect 30012 10668 30064 10674
rect 30012 10610 30064 10616
rect 29826 9752 29882 9761
rect 29826 9687 29882 9696
rect 29644 9580 29696 9586
rect 29644 9522 29696 9528
rect 28632 9376 28684 9382
rect 28632 9318 28684 9324
rect 28816 9376 28868 9382
rect 28816 9318 28868 9324
rect 28540 9172 28592 9178
rect 28540 9114 28592 9120
rect 28828 9110 28856 9318
rect 28816 9104 28868 9110
rect 28356 9036 28408 9042
rect 28460 9030 28580 9058
rect 28816 9046 28868 9052
rect 28356 8978 28408 8984
rect 28368 8634 28396 8978
rect 28356 8628 28408 8634
rect 28356 8570 28408 8576
rect 28264 6996 28316 7002
rect 28264 6938 28316 6944
rect 28080 6384 28132 6390
rect 28080 6326 28132 6332
rect 27988 6316 28040 6322
rect 27988 6258 28040 6264
rect 27622 6012 27918 6032
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 28000 5846 28028 6258
rect 27528 5840 27580 5846
rect 27528 5782 27580 5788
rect 27988 5840 28040 5846
rect 27988 5782 28040 5788
rect 27068 5704 27120 5710
rect 27068 5646 27120 5652
rect 27080 5302 27108 5646
rect 27540 5370 27568 5782
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 27528 5364 27580 5370
rect 27528 5306 27580 5312
rect 27068 5296 27120 5302
rect 27068 5238 27120 5244
rect 27264 5098 27292 5306
rect 27252 5092 27304 5098
rect 27252 5034 27304 5040
rect 27540 4826 27568 5306
rect 28000 5234 28028 5782
rect 28092 5574 28120 6326
rect 28080 5568 28132 5574
rect 28080 5510 28132 5516
rect 27988 5228 28040 5234
rect 27988 5170 28040 5176
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 28092 4826 28120 5510
rect 28172 5024 28224 5030
rect 28172 4966 28224 4972
rect 27528 4820 27580 4826
rect 27528 4762 27580 4768
rect 28080 4820 28132 4826
rect 28080 4762 28132 4768
rect 26700 4752 26752 4758
rect 26700 4694 26752 4700
rect 27160 4684 27212 4690
rect 27160 4626 27212 4632
rect 26516 4616 26568 4622
rect 26516 4558 26568 4564
rect 26424 4276 26476 4282
rect 26424 4218 26476 4224
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 26436 4010 26464 4218
rect 26332 4004 26384 4010
rect 26252 3964 26332 3992
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 26160 3369 26188 3538
rect 26252 3398 26280 3964
rect 26332 3946 26384 3952
rect 26424 4004 26476 4010
rect 26424 3946 26476 3952
rect 26240 3392 26292 3398
rect 26146 3360 26202 3369
rect 26240 3334 26292 3340
rect 26332 3392 26384 3398
rect 26332 3334 26384 3340
rect 26146 3295 26202 3304
rect 26252 2650 26280 3334
rect 26344 3058 26372 3334
rect 26332 3052 26384 3058
rect 26332 2994 26384 3000
rect 26528 2922 26556 4558
rect 27172 4282 27200 4626
rect 27712 4616 27764 4622
rect 27712 4558 27764 4564
rect 27436 4548 27488 4554
rect 27488 4508 27568 4536
rect 27436 4490 27488 4496
rect 27160 4276 27212 4282
rect 27160 4218 27212 4224
rect 26976 4004 27028 4010
rect 26976 3946 27028 3952
rect 26988 3534 27016 3946
rect 27540 3602 27568 4508
rect 27724 4214 27752 4558
rect 27712 4208 27764 4214
rect 27712 4150 27764 4156
rect 28184 4146 28212 4966
rect 28276 4690 28304 6938
rect 28448 5840 28500 5846
rect 28448 5782 28500 5788
rect 28460 5370 28488 5782
rect 28448 5364 28500 5370
rect 28448 5306 28500 5312
rect 28264 4684 28316 4690
rect 28264 4626 28316 4632
rect 28276 4214 28304 4626
rect 28264 4208 28316 4214
rect 28264 4150 28316 4156
rect 28172 4140 28224 4146
rect 28172 4082 28224 4088
rect 28552 4078 28580 9030
rect 28828 8294 28856 9046
rect 29644 8356 29696 8362
rect 29644 8298 29696 8304
rect 28816 8288 28868 8294
rect 28816 8230 28868 8236
rect 28828 8022 28856 8230
rect 28816 8016 28868 8022
rect 28816 7958 28868 7964
rect 28828 7410 28856 7958
rect 29656 7886 29684 8298
rect 29460 7880 29512 7886
rect 29460 7822 29512 7828
rect 29644 7880 29696 7886
rect 29644 7822 29696 7828
rect 28908 7540 28960 7546
rect 28908 7482 28960 7488
rect 28816 7404 28868 7410
rect 28816 7346 28868 7352
rect 28816 6928 28868 6934
rect 28816 6870 28868 6876
rect 28724 6792 28776 6798
rect 28724 6734 28776 6740
rect 28632 5704 28684 5710
rect 28632 5646 28684 5652
rect 28644 5234 28672 5646
rect 28736 5370 28764 6734
rect 28828 6458 28856 6870
rect 28920 6458 28948 7482
rect 29472 7206 29500 7822
rect 29460 7200 29512 7206
rect 29460 7142 29512 7148
rect 28816 6452 28868 6458
rect 28816 6394 28868 6400
rect 28908 6452 28960 6458
rect 28908 6394 28960 6400
rect 28828 6186 28856 6394
rect 29184 6316 29236 6322
rect 29184 6258 29236 6264
rect 28816 6180 28868 6186
rect 28816 6122 28868 6128
rect 29000 6112 29052 6118
rect 29000 6054 29052 6060
rect 28724 5364 28776 5370
rect 28724 5306 28776 5312
rect 28632 5228 28684 5234
rect 28632 5170 28684 5176
rect 29012 5098 29040 6054
rect 29196 5914 29224 6258
rect 29368 6180 29420 6186
rect 29368 6122 29420 6128
rect 29184 5908 29236 5914
rect 29184 5850 29236 5856
rect 29196 5642 29224 5850
rect 29380 5710 29408 6122
rect 29368 5704 29420 5710
rect 29368 5646 29420 5652
rect 29184 5636 29236 5642
rect 29184 5578 29236 5584
rect 29000 5092 29052 5098
rect 29000 5034 29052 5040
rect 29472 4758 29500 7142
rect 29644 6792 29696 6798
rect 29644 6734 29696 6740
rect 29656 6322 29684 6734
rect 29644 6316 29696 6322
rect 29644 6258 29696 6264
rect 29840 5370 29868 9687
rect 30024 5760 30052 10610
rect 30104 10532 30156 10538
rect 30104 10474 30156 10480
rect 30116 9926 30144 10474
rect 30300 10198 30328 11494
rect 30564 11076 30616 11082
rect 30564 11018 30616 11024
rect 30576 10742 30604 11018
rect 30564 10736 30616 10742
rect 30564 10678 30616 10684
rect 30656 10532 30708 10538
rect 30656 10474 30708 10480
rect 30288 10192 30340 10198
rect 30288 10134 30340 10140
rect 30564 10192 30616 10198
rect 30564 10134 30616 10140
rect 30104 9920 30156 9926
rect 30104 9862 30156 9868
rect 30116 9178 30144 9862
rect 30300 9722 30328 10134
rect 30288 9716 30340 9722
rect 30288 9658 30340 9664
rect 30576 9654 30604 10134
rect 30564 9648 30616 9654
rect 30564 9590 30616 9596
rect 30104 9172 30156 9178
rect 30104 9114 30156 9120
rect 30564 9036 30616 9042
rect 30668 9024 30696 10474
rect 31116 10464 31168 10470
rect 31116 10406 31168 10412
rect 31128 10062 31156 10406
rect 31116 10056 31168 10062
rect 31116 9998 31168 10004
rect 30748 9444 30800 9450
rect 30748 9386 30800 9392
rect 30616 8996 30696 9024
rect 30564 8978 30616 8984
rect 30196 8832 30248 8838
rect 30196 8774 30248 8780
rect 30208 8362 30236 8774
rect 30288 8560 30340 8566
rect 30288 8502 30340 8508
rect 30104 8356 30156 8362
rect 30104 8298 30156 8304
rect 30196 8356 30248 8362
rect 30196 8298 30248 8304
rect 30116 8090 30144 8298
rect 30104 8084 30156 8090
rect 30104 8026 30156 8032
rect 30208 7954 30236 8298
rect 30196 7948 30248 7954
rect 30196 7890 30248 7896
rect 30104 7880 30156 7886
rect 30104 7822 30156 7828
rect 30116 7410 30144 7822
rect 30104 7404 30156 7410
rect 30104 7346 30156 7352
rect 30300 7002 30328 8502
rect 30472 8288 30524 8294
rect 30472 8230 30524 8236
rect 30288 6996 30340 7002
rect 30288 6938 30340 6944
rect 30484 6866 30512 8230
rect 30576 7818 30604 8978
rect 30760 8809 30788 9386
rect 30932 9036 30984 9042
rect 30932 8978 30984 8984
rect 30746 8800 30802 8809
rect 30746 8735 30802 8744
rect 30944 8566 30972 8978
rect 31220 8634 31248 15506
rect 32508 15475 32536 15506
rect 36634 15056 36690 15065
rect 36634 14991 36690 15000
rect 36266 14240 36322 14249
rect 36266 14175 36322 14184
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 35622 12336 35678 12345
rect 34612 12300 34664 12306
rect 34612 12242 34664 12248
rect 35440 12300 35492 12306
rect 35622 12271 35678 12280
rect 35440 12242 35492 12248
rect 34289 11996 34585 12016
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 33600 11892 33652 11898
rect 33600 11834 33652 11840
rect 32588 11688 32640 11694
rect 32588 11630 32640 11636
rect 31484 11552 31536 11558
rect 31484 11494 31536 11500
rect 31852 11552 31904 11558
rect 31852 11494 31904 11500
rect 31496 11354 31524 11494
rect 31484 11348 31536 11354
rect 31484 11290 31536 11296
rect 31392 11212 31444 11218
rect 31392 11154 31444 11160
rect 31404 10538 31432 11154
rect 31496 10742 31524 11290
rect 31760 10804 31812 10810
rect 31760 10746 31812 10752
rect 31484 10736 31536 10742
rect 31484 10678 31536 10684
rect 31392 10532 31444 10538
rect 31392 10474 31444 10480
rect 31668 10532 31720 10538
rect 31668 10474 31720 10480
rect 31680 10266 31708 10474
rect 31668 10260 31720 10266
rect 31668 10202 31720 10208
rect 31772 9518 31800 10746
rect 31760 9512 31812 9518
rect 31760 9454 31812 9460
rect 31758 9072 31814 9081
rect 31864 9058 31892 11494
rect 32496 11212 32548 11218
rect 32496 11154 32548 11160
rect 32508 10674 32536 11154
rect 32496 10668 32548 10674
rect 32496 10610 32548 10616
rect 32220 10532 32272 10538
rect 32220 10474 32272 10480
rect 32312 10532 32364 10538
rect 32312 10474 32364 10480
rect 32232 10198 32260 10474
rect 32220 10192 32272 10198
rect 32220 10134 32272 10140
rect 32324 9722 32352 10474
rect 32508 10470 32536 10610
rect 32496 10464 32548 10470
rect 32496 10406 32548 10412
rect 32508 9994 32536 10406
rect 32496 9988 32548 9994
rect 32496 9930 32548 9936
rect 32312 9716 32364 9722
rect 32312 9658 32364 9664
rect 32036 9376 32088 9382
rect 32036 9318 32088 9324
rect 31814 9030 31892 9058
rect 31758 9007 31814 9016
rect 31208 8628 31260 8634
rect 31208 8570 31260 8576
rect 30932 8560 30984 8566
rect 30932 8502 30984 8508
rect 30746 7984 30802 7993
rect 30746 7919 30802 7928
rect 30564 7812 30616 7818
rect 30564 7754 30616 7760
rect 30472 6860 30524 6866
rect 30472 6802 30524 6808
rect 30484 6390 30512 6802
rect 30472 6384 30524 6390
rect 30472 6326 30524 6332
rect 30104 5772 30156 5778
rect 30024 5732 30104 5760
rect 30104 5714 30156 5720
rect 30196 5772 30248 5778
rect 30196 5714 30248 5720
rect 30116 5370 30144 5714
rect 29828 5364 29880 5370
rect 29828 5306 29880 5312
rect 30104 5364 30156 5370
rect 30104 5306 30156 5312
rect 29840 5166 29868 5306
rect 29828 5160 29880 5166
rect 29828 5102 29880 5108
rect 30208 4826 30236 5714
rect 30760 5370 30788 7919
rect 31772 7342 31800 9007
rect 32048 8362 32076 9318
rect 32128 9036 32180 9042
rect 32128 8978 32180 8984
rect 32404 9036 32456 9042
rect 32404 8978 32456 8984
rect 32036 8356 32088 8362
rect 32036 8298 32088 8304
rect 31760 7336 31812 7342
rect 31760 7278 31812 7284
rect 32048 7274 32076 8298
rect 32140 8294 32168 8978
rect 32128 8288 32180 8294
rect 32128 8230 32180 8236
rect 32416 8090 32444 8978
rect 32404 8084 32456 8090
rect 32404 8026 32456 8032
rect 32600 7857 32628 11630
rect 33416 11620 33468 11626
rect 33416 11562 33468 11568
rect 32680 11144 32732 11150
rect 32680 11086 32732 11092
rect 32692 10266 32720 11086
rect 33324 10668 33376 10674
rect 33324 10610 33376 10616
rect 32956 10600 33008 10606
rect 32956 10542 33008 10548
rect 32680 10260 32732 10266
rect 32680 10202 32732 10208
rect 32692 9586 32720 10202
rect 32680 9580 32732 9586
rect 32680 9522 32732 9528
rect 32772 9104 32824 9110
rect 32772 9046 32824 9052
rect 32784 8430 32812 9046
rect 32772 8424 32824 8430
rect 32772 8366 32824 8372
rect 32678 7984 32734 7993
rect 32678 7919 32680 7928
rect 32732 7919 32734 7928
rect 32680 7890 32732 7896
rect 32586 7848 32642 7857
rect 32586 7783 32642 7792
rect 32036 7268 32088 7274
rect 32036 7210 32088 7216
rect 32048 6934 32076 7210
rect 32036 6928 32088 6934
rect 32036 6870 32088 6876
rect 31116 6860 31168 6866
rect 31116 6802 31168 6808
rect 31128 6236 31156 6802
rect 32048 6390 32076 6870
rect 32036 6384 32088 6390
rect 32036 6326 32088 6332
rect 32128 6316 32180 6322
rect 32128 6258 32180 6264
rect 31208 6248 31260 6254
rect 31128 6208 31208 6236
rect 31128 5914 31156 6208
rect 31208 6190 31260 6196
rect 31116 5908 31168 5914
rect 31116 5850 31168 5856
rect 32140 5778 32168 6258
rect 32128 5772 32180 5778
rect 32128 5714 32180 5720
rect 30748 5364 30800 5370
rect 30748 5306 30800 5312
rect 30760 5166 30788 5306
rect 31760 5228 31812 5234
rect 31760 5170 31812 5176
rect 30748 5160 30800 5166
rect 31772 5137 31800 5170
rect 30748 5102 30800 5108
rect 31758 5128 31814 5137
rect 31758 5063 31814 5072
rect 30196 4820 30248 4826
rect 30196 4762 30248 4768
rect 29460 4752 29512 4758
rect 29460 4694 29512 4700
rect 29644 4684 29696 4690
rect 29644 4626 29696 4632
rect 29656 4282 29684 4626
rect 30208 4622 30236 4762
rect 30196 4616 30248 4622
rect 30196 4558 30248 4564
rect 29644 4276 29696 4282
rect 29644 4218 29696 4224
rect 31772 4154 31800 5063
rect 32140 5030 32168 5714
rect 32128 5024 32180 5030
rect 32128 4966 32180 4972
rect 32140 4729 32168 4966
rect 32126 4720 32182 4729
rect 32126 4655 32182 4664
rect 32600 4154 32628 7783
rect 32692 7546 32720 7890
rect 32680 7540 32732 7546
rect 32680 7482 32732 7488
rect 32968 6458 32996 10542
rect 33140 10192 33192 10198
rect 33140 10134 33192 10140
rect 33152 9722 33180 10134
rect 33140 9716 33192 9722
rect 33140 9658 33192 9664
rect 33336 9042 33364 10610
rect 33324 9036 33376 9042
rect 33324 8978 33376 8984
rect 33428 8906 33456 11562
rect 33416 8900 33468 8906
rect 33416 8842 33468 8848
rect 33508 7880 33560 7886
rect 33508 7822 33560 7828
rect 33324 7812 33376 7818
rect 33324 7754 33376 7760
rect 33336 7274 33364 7754
rect 33416 7744 33468 7750
rect 33416 7686 33468 7692
rect 33428 7410 33456 7686
rect 33416 7404 33468 7410
rect 33416 7346 33468 7352
rect 33428 7274 33456 7346
rect 33324 7268 33376 7274
rect 33324 7210 33376 7216
rect 33416 7268 33468 7274
rect 33416 7210 33468 7216
rect 33336 7002 33364 7210
rect 33324 6996 33376 7002
rect 33324 6938 33376 6944
rect 33520 6662 33548 7822
rect 33048 6656 33100 6662
rect 33048 6598 33100 6604
rect 33324 6656 33376 6662
rect 33324 6598 33376 6604
rect 33508 6656 33560 6662
rect 33508 6598 33560 6604
rect 32956 6452 33008 6458
rect 32956 6394 33008 6400
rect 33060 6390 33088 6598
rect 33048 6384 33100 6390
rect 33048 6326 33100 6332
rect 32680 6248 32732 6254
rect 32680 6190 32732 6196
rect 32692 5914 32720 6190
rect 32680 5908 32732 5914
rect 32680 5850 32732 5856
rect 33336 5846 33364 6598
rect 33324 5840 33376 5846
rect 33324 5782 33376 5788
rect 33612 5778 33640 11834
rect 34428 11756 34480 11762
rect 34428 11698 34480 11704
rect 34152 11212 34204 11218
rect 34152 11154 34204 11160
rect 33692 11076 33744 11082
rect 33692 11018 33744 11024
rect 33704 10198 33732 11018
rect 34058 10840 34114 10849
rect 34164 10810 34192 11154
rect 34440 11082 34468 11698
rect 34624 11626 34652 12242
rect 34796 12096 34848 12102
rect 34796 12038 34848 12044
rect 34612 11620 34664 11626
rect 34612 11562 34664 11568
rect 34428 11076 34480 11082
rect 34428 11018 34480 11024
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 34058 10775 34114 10784
rect 34152 10804 34204 10810
rect 34072 10742 34100 10775
rect 34152 10746 34204 10752
rect 34060 10736 34112 10742
rect 34060 10678 34112 10684
rect 34152 10668 34204 10674
rect 34152 10610 34204 10616
rect 33784 10600 33836 10606
rect 33784 10542 33836 10548
rect 33692 10192 33744 10198
rect 33692 10134 33744 10140
rect 33796 8974 33824 10542
rect 34164 9761 34192 10610
rect 34612 10464 34664 10470
rect 34612 10406 34664 10412
rect 34624 10062 34652 10406
rect 34704 10192 34756 10198
rect 34704 10134 34756 10140
rect 34612 10056 34664 10062
rect 34612 9998 34664 10004
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34150 9752 34206 9761
rect 34289 9744 34585 9764
rect 34624 9722 34652 9998
rect 34150 9687 34206 9696
rect 34612 9716 34664 9722
rect 34612 9658 34664 9664
rect 34336 9376 34388 9382
rect 34336 9318 34388 9324
rect 34060 9172 34112 9178
rect 34060 9114 34112 9120
rect 33784 8968 33836 8974
rect 33784 8910 33836 8916
rect 34072 8634 34100 9114
rect 34348 9042 34376 9318
rect 34716 9042 34744 10134
rect 34808 9586 34836 12038
rect 35452 11898 35480 12242
rect 35636 11898 35664 12271
rect 35440 11892 35492 11898
rect 35440 11834 35492 11840
rect 35624 11892 35676 11898
rect 35624 11834 35676 11840
rect 35164 11688 35216 11694
rect 35164 11630 35216 11636
rect 34888 11552 34940 11558
rect 34888 11494 34940 11500
rect 34900 10198 34928 11494
rect 35072 11144 35124 11150
rect 35072 11086 35124 11092
rect 34980 11008 35032 11014
rect 34980 10950 35032 10956
rect 34992 10538 35020 10950
rect 35084 10538 35112 11086
rect 34980 10532 35032 10538
rect 34980 10474 35032 10480
rect 35072 10532 35124 10538
rect 35072 10474 35124 10480
rect 34888 10192 34940 10198
rect 34888 10134 34940 10140
rect 34796 9580 34848 9586
rect 34796 9522 34848 9528
rect 34808 9178 34836 9522
rect 35084 9450 35112 10474
rect 35072 9444 35124 9450
rect 35072 9386 35124 9392
rect 34796 9172 34848 9178
rect 34796 9114 34848 9120
rect 34336 9036 34388 9042
rect 34336 8978 34388 8984
rect 34704 9036 34756 9042
rect 34704 8978 34756 8984
rect 34980 8832 35032 8838
rect 34980 8774 35032 8780
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 34072 8362 34100 8570
rect 34992 8362 35020 8774
rect 34060 8356 34112 8362
rect 34060 8298 34112 8304
rect 34980 8356 35032 8362
rect 34980 8298 35032 8304
rect 34072 8022 34100 8298
rect 34060 8016 34112 8022
rect 34060 7958 34112 7964
rect 34072 7546 34100 7958
rect 34888 7744 34940 7750
rect 34888 7686 34940 7692
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34289 7568 34585 7588
rect 34060 7540 34112 7546
rect 34060 7482 34112 7488
rect 34900 7478 34928 7686
rect 34888 7472 34940 7478
rect 34888 7414 34940 7420
rect 34992 7206 35020 8298
rect 35176 7954 35204 11630
rect 35622 11520 35678 11529
rect 35622 11455 35678 11464
rect 35636 11354 35664 11455
rect 35624 11348 35676 11354
rect 35624 11290 35676 11296
rect 35440 11212 35492 11218
rect 35440 11154 35492 11160
rect 35452 10674 35480 11154
rect 35440 10668 35492 10674
rect 35440 10610 35492 10616
rect 35624 10532 35676 10538
rect 35624 10474 35676 10480
rect 35256 9988 35308 9994
rect 35256 9930 35308 9936
rect 35268 9586 35296 9930
rect 35636 9926 35664 10474
rect 36084 10464 36136 10470
rect 36084 10406 36136 10412
rect 36096 10130 36124 10406
rect 36280 10266 36308 14175
rect 36648 10810 36676 14991
rect 37200 11898 37228 15558
rect 37462 15520 37518 15558
rect 39578 13800 39634 13809
rect 39578 13735 39634 13744
rect 39592 12442 39620 13735
rect 39580 12436 39632 12442
rect 39580 12378 39632 12384
rect 37188 11892 37240 11898
rect 37188 11834 37240 11840
rect 37004 11212 37056 11218
rect 37004 11154 37056 11160
rect 36728 11008 36780 11014
rect 36728 10950 36780 10956
rect 36740 10849 36768 10950
rect 36726 10840 36782 10849
rect 36636 10804 36688 10810
rect 37016 10810 37044 11154
rect 39580 11076 39632 11082
rect 39580 11018 39632 11024
rect 36726 10775 36782 10784
rect 37004 10804 37056 10810
rect 36636 10746 36688 10752
rect 37004 10746 37056 10752
rect 37016 10713 37044 10746
rect 37002 10704 37058 10713
rect 37002 10639 37058 10648
rect 39592 10305 39620 11018
rect 39578 10296 39634 10305
rect 36268 10260 36320 10266
rect 39578 10231 39634 10240
rect 36268 10202 36320 10208
rect 36544 10192 36596 10198
rect 36544 10134 36596 10140
rect 36084 10124 36136 10130
rect 36084 10066 36136 10072
rect 35624 9920 35676 9926
rect 35624 9862 35676 9868
rect 35636 9586 35664 9862
rect 35256 9580 35308 9586
rect 35256 9522 35308 9528
rect 35624 9580 35676 9586
rect 35624 9522 35676 9528
rect 36096 9489 36124 10066
rect 36082 9480 36138 9489
rect 36556 9450 36584 10134
rect 36082 9415 36138 9424
rect 36360 9444 36412 9450
rect 36096 9382 36124 9415
rect 36360 9386 36412 9392
rect 36544 9444 36596 9450
rect 36544 9386 36596 9392
rect 36636 9444 36688 9450
rect 36636 9386 36688 9392
rect 36084 9376 36136 9382
rect 36084 9318 36136 9324
rect 36372 9178 36400 9386
rect 36648 9178 36676 9386
rect 35808 9172 35860 9178
rect 35808 9114 35860 9120
rect 36360 9172 36412 9178
rect 36360 9114 36412 9120
rect 36636 9172 36688 9178
rect 36636 9114 36688 9120
rect 35820 8634 35848 9114
rect 36268 8968 36320 8974
rect 36268 8910 36320 8916
rect 36280 8634 36308 8910
rect 39580 8900 39632 8906
rect 39580 8842 39632 8848
rect 36634 8800 36690 8809
rect 36634 8735 36690 8744
rect 36648 8634 36676 8735
rect 35808 8628 35860 8634
rect 35808 8570 35860 8576
rect 36268 8628 36320 8634
rect 36268 8570 36320 8576
rect 36636 8628 36688 8634
rect 36636 8570 36688 8576
rect 35624 8492 35676 8498
rect 35624 8434 35676 8440
rect 35440 8016 35492 8022
rect 35440 7958 35492 7964
rect 35164 7948 35216 7954
rect 35164 7890 35216 7896
rect 35348 7880 35400 7886
rect 35348 7822 35400 7828
rect 35360 7410 35388 7822
rect 35452 7546 35480 7958
rect 35636 7886 35664 8434
rect 36268 8424 36320 8430
rect 36268 8366 36320 8372
rect 35624 7880 35676 7886
rect 35624 7822 35676 7828
rect 35440 7540 35492 7546
rect 35440 7482 35492 7488
rect 35348 7404 35400 7410
rect 35348 7346 35400 7352
rect 35164 7268 35216 7274
rect 35164 7210 35216 7216
rect 34060 7200 34112 7206
rect 34060 7142 34112 7148
rect 34980 7200 35032 7206
rect 34980 7142 35032 7148
rect 33876 6792 33928 6798
rect 33876 6734 33928 6740
rect 33888 6458 33916 6734
rect 33876 6452 33928 6458
rect 33876 6394 33928 6400
rect 34072 6361 34100 7142
rect 34612 6928 34664 6934
rect 34612 6870 34664 6876
rect 34152 6792 34204 6798
rect 34152 6734 34204 6740
rect 34058 6352 34114 6361
rect 34058 6287 34114 6296
rect 34164 5914 34192 6734
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 34624 6390 34652 6870
rect 34612 6384 34664 6390
rect 34612 6326 34664 6332
rect 35176 6322 35204 7210
rect 35360 7002 35388 7346
rect 35348 6996 35400 7002
rect 35348 6938 35400 6944
rect 35360 6322 35388 6938
rect 36176 6928 36228 6934
rect 36176 6870 36228 6876
rect 36084 6792 36136 6798
rect 36084 6734 36136 6740
rect 36096 6458 36124 6734
rect 36084 6452 36136 6458
rect 36084 6394 36136 6400
rect 36188 6390 36216 6870
rect 36176 6384 36228 6390
rect 36176 6326 36228 6332
rect 35164 6316 35216 6322
rect 35164 6258 35216 6264
rect 35348 6316 35400 6322
rect 35348 6258 35400 6264
rect 34612 6248 34664 6254
rect 34612 6190 34664 6196
rect 34624 6118 34652 6190
rect 34980 6180 35032 6186
rect 34980 6122 35032 6128
rect 34612 6112 34664 6118
rect 34612 6054 34664 6060
rect 34152 5908 34204 5914
rect 34152 5850 34204 5856
rect 34624 5846 34652 6054
rect 34992 5914 35020 6122
rect 34980 5908 35032 5914
rect 34980 5850 35032 5856
rect 34612 5840 34664 5846
rect 34612 5782 34664 5788
rect 33600 5772 33652 5778
rect 33600 5714 33652 5720
rect 33612 5681 33640 5714
rect 34152 5704 34204 5710
rect 33598 5672 33654 5681
rect 34152 5646 34204 5652
rect 33598 5607 33654 5616
rect 33612 5370 33640 5607
rect 34164 5370 34192 5646
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 34289 5392 34585 5412
rect 34624 5370 34652 5782
rect 34992 5370 35020 5850
rect 36280 5778 36308 8366
rect 36634 7984 36690 7993
rect 36634 7919 36690 7928
rect 36648 7546 36676 7919
rect 36636 7540 36688 7546
rect 36636 7482 36688 7488
rect 36360 7200 36412 7206
rect 36360 7142 36412 7148
rect 36372 6798 36400 7142
rect 36360 6792 36412 6798
rect 36360 6734 36412 6740
rect 36372 5846 36400 6734
rect 39592 6633 39620 8842
rect 39578 6624 39634 6633
rect 39578 6559 39634 6568
rect 36452 6452 36504 6458
rect 36452 6394 36504 6400
rect 36464 5914 36492 6394
rect 36912 6112 36964 6118
rect 36912 6054 36964 6060
rect 36452 5908 36504 5914
rect 36452 5850 36504 5856
rect 36360 5840 36412 5846
rect 36360 5782 36412 5788
rect 36268 5772 36320 5778
rect 36268 5714 36320 5720
rect 36280 5370 36308 5714
rect 33600 5364 33652 5370
rect 33600 5306 33652 5312
rect 34152 5364 34204 5370
rect 34152 5306 34204 5312
rect 34612 5364 34664 5370
rect 34612 5306 34664 5312
rect 34980 5364 35032 5370
rect 34980 5306 35032 5312
rect 35992 5364 36044 5370
rect 35992 5306 36044 5312
rect 36268 5364 36320 5370
rect 36268 5306 36320 5312
rect 35440 5024 35492 5030
rect 35440 4966 35492 4972
rect 35452 4865 35480 4966
rect 35438 4856 35494 4865
rect 35438 4791 35494 4800
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 35452 4282 35480 4791
rect 35440 4276 35492 4282
rect 35440 4218 35492 4224
rect 29828 4140 29880 4146
rect 31772 4126 31892 4154
rect 29828 4082 29880 4088
rect 28540 4072 28592 4078
rect 29840 4049 29868 4082
rect 30288 4072 30340 4078
rect 28540 4014 28592 4020
rect 29826 4040 29882 4049
rect 30288 4014 30340 4020
rect 29826 3975 29882 3984
rect 27622 3836 27918 3856
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 29092 3732 29144 3738
rect 29092 3674 29144 3680
rect 28448 3664 28500 3670
rect 28448 3606 28500 3612
rect 27252 3596 27304 3602
rect 27252 3538 27304 3544
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 26976 3528 27028 3534
rect 26976 3470 27028 3476
rect 26988 2922 27016 3470
rect 27264 3194 27292 3538
rect 27540 3194 27568 3538
rect 27988 3460 28040 3466
rect 27988 3402 28040 3408
rect 28000 3194 28028 3402
rect 27252 3188 27304 3194
rect 27252 3130 27304 3136
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 27988 3188 28040 3194
rect 27988 3130 28040 3136
rect 26516 2916 26568 2922
rect 26516 2858 26568 2864
rect 26976 2916 27028 2922
rect 26976 2858 27028 2864
rect 26240 2644 26292 2650
rect 26240 2586 26292 2592
rect 27264 2009 27292 3130
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27724 2961 27752 2994
rect 27710 2952 27766 2961
rect 27710 2887 27766 2896
rect 28460 2854 28488 3606
rect 28448 2848 28500 2854
rect 28448 2790 28500 2796
rect 27622 2748 27918 2768
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 27622 2672 27918 2692
rect 27436 2508 27488 2514
rect 27436 2450 27488 2456
rect 27448 2417 27476 2450
rect 27434 2408 27490 2417
rect 27434 2343 27490 2352
rect 27448 2310 27476 2343
rect 27436 2304 27488 2310
rect 27436 2246 27488 2252
rect 28264 2304 28316 2310
rect 28264 2246 28316 2252
rect 27250 2000 27306 2009
rect 27250 1935 27306 1944
rect 27448 1329 27476 2246
rect 28276 1329 28304 2246
rect 27434 1320 27490 1329
rect 27434 1255 27490 1264
rect 28262 1320 28318 1329
rect 28262 1255 28318 1264
rect 24688 54 25006 82
rect 25412 128 25464 134
rect 25412 70 25464 76
rect 28354 82 28410 480
rect 28460 82 28488 2790
rect 29104 2650 29132 3674
rect 30104 3460 30156 3466
rect 30104 3402 30156 3408
rect 30116 3058 30144 3402
rect 30300 3097 30328 4014
rect 30472 3936 30524 3942
rect 30472 3878 30524 3884
rect 30286 3088 30342 3097
rect 29460 3052 29512 3058
rect 29460 2994 29512 3000
rect 30104 3052 30156 3058
rect 30286 3023 30342 3032
rect 30104 2994 30156 3000
rect 29472 2650 29500 2994
rect 29552 2916 29604 2922
rect 29552 2858 29604 2864
rect 29092 2644 29144 2650
rect 29092 2586 29144 2592
rect 29460 2644 29512 2650
rect 29460 2586 29512 2592
rect 29564 2582 29592 2858
rect 29828 2848 29880 2854
rect 29828 2790 29880 2796
rect 29552 2576 29604 2582
rect 29552 2518 29604 2524
rect 29840 2514 29868 2790
rect 30116 2514 30144 2994
rect 30484 2961 30512 3878
rect 30748 3528 30800 3534
rect 30748 3470 30800 3476
rect 30760 3194 30788 3470
rect 30748 3188 30800 3194
rect 30748 3130 30800 3136
rect 30470 2952 30526 2961
rect 30470 2887 30526 2896
rect 29828 2508 29880 2514
rect 29828 2450 29880 2456
rect 30104 2508 30156 2514
rect 30104 2450 30156 2456
rect 31864 1057 31892 4126
rect 32508 4126 32628 4154
rect 32508 2825 32536 4126
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 34289 3216 34585 3236
rect 32494 2816 32550 2825
rect 32494 2751 32550 2760
rect 36004 2417 36032 5306
rect 35990 2408 36046 2417
rect 35990 2343 36046 2352
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 36924 1873 36952 6054
rect 38384 2372 38436 2378
rect 38384 2314 38436 2320
rect 36910 1864 36966 1873
rect 36910 1799 36966 1808
rect 35070 1320 35126 1329
rect 35070 1255 35126 1264
rect 31850 1048 31906 1057
rect 31850 983 31906 992
rect 11610 0 11666 54
rect 15014 0 15070 54
rect 18326 0 18382 54
rect 21638 0 21694 54
rect 24950 0 25006 54
rect 28354 54 28488 82
rect 31666 128 31722 480
rect 31666 76 31668 128
rect 31720 76 31722 128
rect 28354 0 28410 54
rect 31666 0 31722 76
rect 34978 82 35034 480
rect 35084 82 35112 1255
rect 34978 54 35112 82
rect 38290 82 38346 480
rect 38396 82 38424 2314
rect 38290 54 38424 82
rect 34978 0 35034 54
rect 38290 0 38346 54
<< via2 >>
rect 2686 15000 2742 15056
rect 1582 14184 1638 14240
rect 110 13744 166 13800
rect 110 12008 166 12064
rect 1582 10784 1638 10840
rect 1398 10648 1454 10704
rect 110 10240 166 10296
rect 754 6704 810 6760
rect 1398 4528 1454 4584
rect 754 3576 810 3632
rect 1674 8472 1730 8528
rect 1582 7928 1638 7984
rect 2226 9968 2282 10024
rect 5814 12280 5870 12336
rect 2226 7792 2282 7848
rect 3054 9968 3110 10024
rect 2042 6160 2098 6216
rect 3146 8880 3202 8936
rect 3330 8472 3386 8528
rect 1674 4120 1730 4176
rect 2134 3984 2190 4040
rect 3606 6160 3662 6216
rect 3974 8744 4030 8800
rect 4618 4528 4674 4584
rect 4618 3984 4674 4040
rect 5078 5616 5134 5672
rect 4894 3848 4950 3904
rect 110 2216 166 2272
rect 4250 1944 4306 2000
rect 4342 992 4398 1048
rect 1950 312 2006 368
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 6642 11736 6698 11792
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 6090 4120 6146 4176
rect 6274 3032 6330 3088
rect 8022 8744 8078 8800
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 7470 6296 7526 6352
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 7286 3848 7342 3904
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 8390 9444 8446 9480
rect 8390 9424 8392 9444
rect 8392 9424 8444 9444
rect 8444 9424 8446 9444
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 9494 7792 9550 7848
rect 9678 9560 9734 9616
rect 10506 7928 10562 7984
rect 9954 7384 10010 7440
rect 9862 7248 9918 7304
rect 9954 6704 10010 6760
rect 8666 6024 8722 6080
rect 9034 4120 9090 4176
rect 9126 3984 9182 4040
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 11150 7384 11206 7440
rect 10966 7248 11022 7304
rect 12162 7248 12218 7304
rect 11426 5072 11482 5128
rect 10506 4936 10562 4992
rect 11426 4528 11482 4584
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 12346 6160 12402 6216
rect 12438 4528 12494 4584
rect 13542 7928 13598 7984
rect 13634 6296 13690 6352
rect 12530 4120 12586 4176
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 14094 6024 14150 6080
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 14554 5072 14610 5128
rect 12254 2760 12310 2816
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 13910 3440 13966 3496
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 14370 3440 14426 3496
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 14830 2624 14886 2680
rect 12346 2488 12402 2544
rect 11978 2216 12034 2272
rect 13358 1944 13414 2000
rect 13358 1264 13414 1320
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 17498 9460 17500 9480
rect 17500 9460 17552 9480
rect 17552 9460 17554 9480
rect 17498 9424 17554 9460
rect 16394 4528 16450 4584
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 17958 8472 18014 8528
rect 17958 8200 18014 8256
rect 17774 4800 17830 4856
rect 18786 9968 18842 10024
rect 17130 3032 17186 3088
rect 15198 312 15254 368
rect 18510 2624 18566 2680
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 20810 9560 20866 9616
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 21362 10648 21418 10704
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 20626 7384 20682 7440
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 21730 9696 21786 9752
rect 22834 10648 22890 10704
rect 22006 9560 22062 9616
rect 18970 3848 19026 3904
rect 18786 3032 18842 3088
rect 19246 3440 19302 3496
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 19890 2896 19946 2952
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 21638 5072 21694 5128
rect 22466 7248 22522 7304
rect 24214 11756 24270 11792
rect 24214 11736 24216 11756
rect 24216 11736 24268 11756
rect 24268 11736 24270 11756
rect 24122 10784 24178 10840
rect 24122 9968 24178 10024
rect 21638 4120 21694 4176
rect 20902 2760 20958 2816
rect 23018 4800 23074 4856
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 25042 6296 25098 6352
rect 25318 8200 25374 8256
rect 23478 4664 23534 4720
rect 23294 3304 23350 3360
rect 24674 4800 24730 4856
rect 24122 3848 24178 3904
rect 23754 2760 23810 2816
rect 24674 2624 24730 2680
rect 20810 2488 20866 2544
rect 22098 2488 22154 2544
rect 24030 2352 24086 2408
rect 20626 2216 20682 2272
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 24858 2352 24914 2408
rect 27066 9696 27122 9752
rect 26790 8200 26846 8256
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 26790 7384 26846 7440
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 29826 9696 29882 9752
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 26146 3304 26202 3360
rect 30746 8744 30802 8800
rect 36634 15000 36690 15056
rect 36266 14184 36322 14240
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 35622 12280 35678 12336
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 31758 9016 31814 9072
rect 30746 7928 30802 7984
rect 32678 7948 32734 7984
rect 32678 7928 32680 7948
rect 32680 7928 32732 7948
rect 32732 7928 32734 7948
rect 32586 7792 32642 7848
rect 31758 5072 31814 5128
rect 32126 4664 32182 4720
rect 34058 10784 34114 10840
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 34150 9696 34206 9752
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 35622 11464 35678 11520
rect 39578 13744 39634 13800
rect 36726 10784 36782 10840
rect 37002 10648 37058 10704
rect 39578 10240 39634 10296
rect 36082 9424 36138 9480
rect 36634 8744 36690 8800
rect 34058 6296 34114 6352
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 33598 5616 33654 5672
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 36634 7928 36690 7984
rect 39578 6568 39634 6624
rect 35438 4800 35494 4856
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 29826 3984 29882 4040
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 27710 2896 27766 2952
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 27434 2352 27490 2408
rect 27250 1944 27306 2000
rect 27434 1264 27490 1320
rect 28262 1264 28318 1320
rect 30286 3032 30342 3088
rect 30470 2896 30526 2952
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 32494 2760 32550 2816
rect 35990 2352 36046 2408
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 36910 1808 36966 1864
rect 35070 1264 35126 1320
rect 31850 992 31906 1048
<< metal3 >>
rect 0 15512 480 15632
rect 39520 15512 40000 15632
rect 62 15058 122 15512
rect 2681 15058 2747 15061
rect 62 15056 2747 15058
rect 62 15000 2686 15056
rect 2742 15000 2747 15056
rect 62 14998 2747 15000
rect 2681 14995 2747 14998
rect 36629 15058 36695 15061
rect 39622 15058 39682 15512
rect 36629 15056 39682 15058
rect 36629 15000 36634 15056
rect 36690 15000 39682 15056
rect 36629 14998 39682 15000
rect 36629 14995 36695 14998
rect 0 14560 480 14680
rect 39520 14560 40000 14680
rect 62 14242 122 14560
rect 1577 14242 1643 14245
rect 62 14240 1643 14242
rect 62 14184 1582 14240
rect 1638 14184 1643 14240
rect 62 14182 1643 14184
rect 1577 14179 1643 14182
rect 36261 14242 36327 14245
rect 39622 14242 39682 14560
rect 36261 14240 39682 14242
rect 36261 14184 36266 14240
rect 36322 14184 39682 14240
rect 36261 14182 39682 14184
rect 36261 14179 36327 14182
rect 0 13800 480 13864
rect 39520 13802 40000 13864
rect 0 13744 110 13800
rect 166 13744 480 13800
rect 39492 13800 40000 13802
rect 39492 13744 39578 13800
rect 39634 13744 40000 13800
rect 105 13742 252 13744
rect 39492 13742 39639 13744
rect 105 13739 171 13742
rect 39573 13739 39639 13742
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 7610 13088 7930 13089
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 13023 34597 13024
rect 0 12792 480 12912
rect 39520 12792 40000 12912
rect 62 12338 122 12792
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 12479 27930 12480
rect 5809 12338 5875 12341
rect 62 12336 5875 12338
rect 62 12280 5814 12336
rect 5870 12280 5875 12336
rect 62 12278 5875 12280
rect 5809 12275 5875 12278
rect 35617 12338 35683 12341
rect 39622 12338 39682 12792
rect 35617 12336 39682 12338
rect 35617 12280 35622 12336
rect 35678 12280 39682 12336
rect 35617 12278 39682 12280
rect 35617 12275 35683 12278
rect 0 12064 480 12096
rect 0 12008 110 12064
rect 166 12008 480 12064
rect 0 11976 480 12008
rect 7610 12000 7930 12001
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 39520 11976 40000 12096
rect 34277 11935 34597 11936
rect 6637 11794 6703 11797
rect 24209 11794 24275 11797
rect 6637 11792 24275 11794
rect 6637 11736 6642 11792
rect 6698 11736 24214 11792
rect 24270 11736 24275 11792
rect 6637 11734 24275 11736
rect 6637 11731 6703 11734
rect 24209 11731 24275 11734
rect 35617 11522 35683 11525
rect 39622 11522 39682 11976
rect 35617 11520 39682 11522
rect 35617 11464 35622 11520
rect 35678 11464 39682 11520
rect 35617 11462 39682 11464
rect 35617 11459 35683 11462
rect 14277 11456 14597 11457
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 11391 27930 11392
rect 0 11116 480 11144
rect 0 11052 60 11116
rect 124 11052 480 11116
rect 39520 11116 40000 11144
rect 39520 11114 39620 11116
rect 39492 11054 39620 11114
rect 0 11024 480 11052
rect 39520 11052 39620 11054
rect 39684 11052 40000 11116
rect 39520 11024 40000 11052
rect 7610 10912 7930 10913
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 10847 34597 10848
rect 54 10780 60 10844
rect 124 10842 130 10844
rect 1577 10842 1643 10845
rect 124 10840 1643 10842
rect 124 10784 1582 10840
rect 1638 10784 1643 10840
rect 124 10782 1643 10784
rect 124 10780 130 10782
rect 1577 10779 1643 10782
rect 24117 10842 24183 10845
rect 34053 10842 34119 10845
rect 24117 10840 34119 10842
rect 24117 10784 24122 10840
rect 24178 10784 34058 10840
rect 34114 10784 34119 10840
rect 24117 10782 34119 10784
rect 24117 10779 24183 10782
rect 34053 10779 34119 10782
rect 36721 10842 36787 10845
rect 39614 10842 39620 10844
rect 36721 10840 39620 10842
rect 36721 10784 36726 10840
rect 36782 10784 39620 10840
rect 36721 10782 39620 10784
rect 36721 10779 36787 10782
rect 39614 10780 39620 10782
rect 39684 10780 39690 10844
rect 1393 10706 1459 10709
rect 21357 10706 21423 10709
rect 1393 10704 21423 10706
rect 1393 10648 1398 10704
rect 1454 10648 21362 10704
rect 21418 10648 21423 10704
rect 1393 10646 21423 10648
rect 1393 10643 1459 10646
rect 21357 10643 21423 10646
rect 22829 10706 22895 10709
rect 36997 10706 37063 10709
rect 22829 10704 37063 10706
rect 22829 10648 22834 10704
rect 22890 10648 37002 10704
rect 37058 10648 37063 10704
rect 22829 10646 37063 10648
rect 22829 10643 22895 10646
rect 36997 10643 37063 10646
rect 14277 10368 14597 10369
rect 0 10296 480 10328
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 10303 27930 10304
rect 39520 10298 40000 10328
rect 0 10240 110 10296
rect 166 10240 480 10296
rect 0 10208 480 10240
rect 39492 10296 40000 10298
rect 39492 10240 39578 10296
rect 39634 10240 40000 10296
rect 39492 10238 40000 10240
rect 39520 10208 40000 10238
rect 2221 10026 2287 10029
rect 3049 10026 3115 10029
rect 18781 10026 18847 10029
rect 24117 10026 24183 10029
rect 2221 10024 24183 10026
rect 2221 9968 2226 10024
rect 2282 9968 3054 10024
rect 3110 9968 18786 10024
rect 18842 9968 24122 10024
rect 24178 9968 24183 10024
rect 2221 9966 24183 9968
rect 2221 9963 2287 9966
rect 3049 9963 3115 9966
rect 18781 9963 18847 9966
rect 24117 9963 24183 9966
rect 7610 9824 7930 9825
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 9759 34597 9760
rect 21725 9754 21791 9757
rect 27061 9754 27127 9757
rect 21725 9752 27127 9754
rect 21725 9696 21730 9752
rect 21786 9696 27066 9752
rect 27122 9696 27127 9752
rect 21725 9694 27127 9696
rect 21725 9691 21791 9694
rect 27061 9691 27127 9694
rect 29821 9754 29887 9757
rect 34145 9754 34211 9757
rect 29821 9752 34211 9754
rect 29821 9696 29826 9752
rect 29882 9696 34150 9752
rect 34206 9696 34211 9752
rect 29821 9694 34211 9696
rect 29821 9691 29887 9694
rect 34145 9691 34211 9694
rect 9673 9618 9739 9621
rect 20805 9618 20871 9621
rect 22001 9618 22067 9621
rect 9673 9616 22067 9618
rect 9673 9560 9678 9616
rect 9734 9560 20810 9616
rect 20866 9560 22006 9616
rect 22062 9560 22067 9616
rect 9673 9558 22067 9560
rect 9673 9555 9739 9558
rect 20805 9555 20871 9558
rect 22001 9555 22067 9558
rect 8385 9482 8451 9485
rect 17493 9482 17559 9485
rect 36077 9482 36143 9485
rect 8385 9480 36143 9482
rect 8385 9424 8390 9480
rect 8446 9424 17498 9480
rect 17554 9424 36082 9480
rect 36138 9424 36143 9480
rect 8385 9422 36143 9424
rect 8385 9419 8451 9422
rect 17493 9419 17559 9422
rect 36077 9419 36143 9422
rect 0 9256 480 9376
rect 14277 9280 14597 9281
rect 62 8802 122 9256
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 39520 9256 40000 9376
rect 27610 9215 27930 9216
rect 31753 9074 31819 9077
rect 13770 9072 31819 9074
rect 13770 9016 31758 9072
rect 31814 9016 31819 9072
rect 13770 9014 31819 9016
rect 3141 8938 3207 8941
rect 13770 8938 13830 9014
rect 31753 9011 31819 9014
rect 3141 8936 13830 8938
rect 3141 8880 3146 8936
rect 3202 8880 13830 8936
rect 3141 8878 13830 8880
rect 18646 8878 21466 8938
rect 3141 8875 3207 8878
rect 3969 8802 4035 8805
rect 62 8800 4035 8802
rect 62 8744 3974 8800
rect 4030 8744 4035 8800
rect 62 8742 4035 8744
rect 3969 8739 4035 8742
rect 8017 8802 8083 8805
rect 18646 8802 18706 8878
rect 8017 8800 18706 8802
rect 8017 8744 8022 8800
rect 8078 8744 18706 8800
rect 8017 8742 18706 8744
rect 21406 8802 21466 8878
rect 30741 8802 30807 8805
rect 21406 8800 30807 8802
rect 21406 8744 30746 8800
rect 30802 8744 30807 8800
rect 21406 8742 30807 8744
rect 8017 8739 8083 8742
rect 30741 8739 30807 8742
rect 36629 8802 36695 8805
rect 39622 8802 39682 9256
rect 36629 8800 39682 8802
rect 36629 8744 36634 8800
rect 36690 8744 39682 8800
rect 36629 8742 39682 8744
rect 36629 8739 36695 8742
rect 7610 8736 7930 8737
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 8671 34597 8672
rect 0 8440 480 8560
rect 1669 8530 1735 8533
rect 3325 8530 3391 8533
rect 17953 8530 18019 8533
rect 1669 8528 18019 8530
rect 1669 8472 1674 8528
rect 1730 8472 3330 8528
rect 3386 8472 17958 8528
rect 18014 8472 18019 8528
rect 1669 8470 18019 8472
rect 1669 8467 1735 8470
rect 3325 8467 3391 8470
rect 17953 8467 18019 8470
rect 39520 8440 40000 8560
rect 62 7986 122 8440
rect 17953 8258 18019 8261
rect 25313 8258 25379 8261
rect 26785 8258 26851 8261
rect 17953 8256 26851 8258
rect 17953 8200 17958 8256
rect 18014 8200 25318 8256
rect 25374 8200 26790 8256
rect 26846 8200 26851 8256
rect 17953 8198 26851 8200
rect 17953 8195 18019 8198
rect 25313 8195 25379 8198
rect 26785 8195 26851 8198
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 8127 27930 8128
rect 1577 7986 1643 7989
rect 62 7984 1643 7986
rect 62 7928 1582 7984
rect 1638 7928 1643 7984
rect 62 7926 1643 7928
rect 1577 7923 1643 7926
rect 10501 7986 10567 7989
rect 13537 7986 13603 7989
rect 30741 7986 30807 7989
rect 32673 7986 32739 7989
rect 10501 7984 32739 7986
rect 10501 7928 10506 7984
rect 10562 7928 13542 7984
rect 13598 7928 30746 7984
rect 30802 7928 32678 7984
rect 32734 7928 32739 7984
rect 10501 7926 32739 7928
rect 10501 7923 10567 7926
rect 13537 7923 13603 7926
rect 30741 7923 30807 7926
rect 32673 7923 32739 7926
rect 36629 7986 36695 7989
rect 39622 7986 39682 8440
rect 36629 7984 39682 7986
rect 36629 7928 36634 7984
rect 36690 7928 39682 7984
rect 36629 7926 39682 7928
rect 36629 7923 36695 7926
rect 2221 7850 2287 7853
rect 62 7848 2287 7850
rect 62 7792 2226 7848
rect 2282 7792 2287 7848
rect 62 7790 2287 7792
rect 62 7608 122 7790
rect 2221 7787 2287 7790
rect 9489 7850 9555 7853
rect 32581 7850 32647 7853
rect 9489 7848 32647 7850
rect 9489 7792 9494 7848
rect 9550 7792 32586 7848
rect 32642 7792 32647 7848
rect 9489 7790 32647 7792
rect 9489 7787 9555 7790
rect 32581 7787 32647 7790
rect 7610 7648 7930 7649
rect 0 7488 480 7608
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 7583 34597 7584
rect 39520 7580 40000 7608
rect 39520 7578 39620 7580
rect 39492 7518 39620 7578
rect 39520 7516 39620 7518
rect 39684 7516 40000 7580
rect 39520 7488 40000 7516
rect 9949 7442 10015 7445
rect 11145 7442 11211 7445
rect 20621 7442 20687 7445
rect 9949 7440 20687 7442
rect 9949 7384 9954 7440
rect 10010 7384 11150 7440
rect 11206 7384 20626 7440
rect 20682 7384 20687 7440
rect 9949 7382 20687 7384
rect 9949 7379 10015 7382
rect 11145 7379 11211 7382
rect 20621 7379 20687 7382
rect 26785 7442 26851 7445
rect 26785 7440 29010 7442
rect 26785 7384 26790 7440
rect 26846 7384 29010 7440
rect 26785 7382 29010 7384
rect 26785 7379 26851 7382
rect 9857 7306 9923 7309
rect 10961 7306 11027 7309
rect 9857 7304 11027 7306
rect 9857 7248 9862 7304
rect 9918 7248 10966 7304
rect 11022 7248 11027 7304
rect 9857 7246 11027 7248
rect 9857 7243 9923 7246
rect 10961 7243 11027 7246
rect 12157 7306 12223 7309
rect 22461 7306 22527 7309
rect 12157 7304 22527 7306
rect 12157 7248 12162 7304
rect 12218 7248 22466 7304
rect 22522 7248 22527 7304
rect 12157 7246 22527 7248
rect 28950 7306 29010 7382
rect 39614 7306 39620 7308
rect 28950 7246 39620 7306
rect 12157 7243 12223 7246
rect 22461 7243 22527 7246
rect 39614 7244 39620 7246
rect 39684 7244 39690 7308
rect 14277 7104 14597 7105
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 7039 27930 7040
rect 749 6762 815 6765
rect 9949 6762 10015 6765
rect 749 6760 10015 6762
rect 749 6704 754 6760
rect 810 6704 9954 6760
rect 10010 6704 10015 6760
rect 749 6702 10015 6704
rect 749 6699 815 6702
rect 9949 6699 10015 6702
rect 0 6536 480 6656
rect 39520 6626 40000 6656
rect 39492 6624 40000 6626
rect 39492 6568 39578 6624
rect 39634 6568 40000 6624
rect 39492 6566 40000 6568
rect 7610 6560 7930 6561
rect 62 6354 122 6536
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 39520 6536 40000 6566
rect 34277 6495 34597 6496
rect 7465 6354 7531 6357
rect 62 6352 7531 6354
rect 62 6296 7470 6352
rect 7526 6296 7531 6352
rect 62 6294 7531 6296
rect 7465 6291 7531 6294
rect 13629 6354 13695 6357
rect 25037 6354 25103 6357
rect 13629 6352 25103 6354
rect 13629 6296 13634 6352
rect 13690 6296 25042 6352
rect 25098 6296 25103 6352
rect 13629 6294 25103 6296
rect 13629 6291 13695 6294
rect 25037 6291 25103 6294
rect 34053 6354 34119 6357
rect 34053 6352 39682 6354
rect 34053 6296 34058 6352
rect 34114 6296 39682 6352
rect 34053 6294 39682 6296
rect 34053 6291 34119 6294
rect 2037 6218 2103 6221
rect 3601 6218 3667 6221
rect 12341 6218 12407 6221
rect 2037 6216 12407 6218
rect 2037 6160 2042 6216
rect 2098 6160 3606 6216
rect 3662 6160 12346 6216
rect 12402 6160 12407 6216
rect 2037 6158 12407 6160
rect 2037 6155 2103 6158
rect 3601 6155 3667 6158
rect 12341 6155 12407 6158
rect 8661 6082 8727 6085
rect 14089 6082 14155 6085
rect 8661 6080 14155 6082
rect 8661 6024 8666 6080
rect 8722 6024 14094 6080
rect 14150 6024 14155 6080
rect 8661 6022 14155 6024
rect 8661 6019 8727 6022
rect 14089 6019 14155 6022
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 5951 27930 5952
rect 39622 5840 39682 6294
rect 0 5720 480 5840
rect 39520 5720 40000 5840
rect 62 5266 122 5720
rect 5073 5674 5139 5677
rect 33593 5674 33659 5677
rect 4110 5672 33659 5674
rect 4110 5616 5078 5672
rect 5134 5616 33598 5672
rect 33654 5616 33659 5672
rect 4110 5614 33659 5616
rect 4110 5266 4170 5614
rect 5073 5611 5139 5614
rect 33593 5611 33659 5614
rect 7610 5472 7930 5473
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 62 5206 4170 5266
rect 54 5068 60 5132
rect 124 5130 130 5132
rect 11421 5130 11487 5133
rect 14549 5130 14615 5133
rect 124 5070 9690 5130
rect 124 5068 130 5070
rect 9630 4994 9690 5070
rect 11421 5128 14615 5130
rect 11421 5072 11426 5128
rect 11482 5072 14554 5128
rect 14610 5072 14615 5128
rect 11421 5070 14615 5072
rect 11421 5067 11487 5070
rect 14549 5067 14615 5070
rect 21633 5130 21699 5133
rect 31753 5130 31819 5133
rect 21633 5128 31819 5130
rect 21633 5072 21638 5128
rect 21694 5072 31758 5128
rect 31814 5072 31819 5128
rect 21633 5070 31819 5072
rect 21633 5067 21699 5070
rect 31753 5067 31819 5070
rect 10501 4994 10567 4997
rect 9630 4992 10567 4994
rect 9630 4936 10506 4992
rect 10562 4936 10567 4992
rect 9630 4934 10567 4936
rect 10501 4931 10567 4934
rect 14277 4928 14597 4929
rect 0 4860 480 4888
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 4863 27930 4864
rect 0 4796 60 4860
rect 124 4796 480 4860
rect 0 4768 480 4796
rect 17769 4858 17835 4861
rect 23013 4858 23079 4861
rect 24669 4858 24735 4861
rect 17769 4856 24735 4858
rect 17769 4800 17774 4856
rect 17830 4800 23018 4856
rect 23074 4800 24674 4856
rect 24730 4800 24735 4856
rect 17769 4798 24735 4800
rect 17769 4795 17835 4798
rect 23013 4795 23079 4798
rect 24669 4795 24735 4798
rect 35433 4858 35499 4861
rect 39520 4858 40000 4888
rect 35433 4856 40000 4858
rect 35433 4800 35438 4856
rect 35494 4800 40000 4856
rect 35433 4798 40000 4800
rect 35433 4795 35499 4798
rect 39520 4768 40000 4798
rect 23473 4722 23539 4725
rect 32121 4722 32187 4725
rect 23473 4720 32187 4722
rect 23473 4664 23478 4720
rect 23534 4664 32126 4720
rect 32182 4664 32187 4720
rect 23473 4662 32187 4664
rect 23473 4659 23539 4662
rect 32121 4659 32187 4662
rect 54 4524 60 4588
rect 124 4586 130 4588
rect 1393 4586 1459 4589
rect 4613 4586 4679 4589
rect 11421 4586 11487 4589
rect 124 4584 1459 4586
rect 124 4528 1398 4584
rect 1454 4528 1459 4584
rect 124 4526 1459 4528
rect 124 4524 130 4526
rect 1393 4523 1459 4526
rect 4110 4584 11487 4586
rect 4110 4528 4618 4584
rect 4674 4528 11426 4584
rect 11482 4528 11487 4584
rect 4110 4526 11487 4528
rect 1669 4178 1735 4181
rect 4110 4178 4170 4526
rect 4613 4523 4679 4526
rect 11421 4523 11487 4526
rect 12433 4586 12499 4589
rect 16389 4586 16455 4589
rect 12433 4584 16455 4586
rect 12433 4528 12438 4584
rect 12494 4528 16394 4584
rect 16450 4528 16455 4584
rect 12433 4526 16455 4528
rect 12433 4523 12499 4526
rect 16389 4523 16455 4526
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 4319 34597 4320
rect 1669 4176 4170 4178
rect 1669 4120 1674 4176
rect 1730 4120 4170 4176
rect 1669 4118 4170 4120
rect 6085 4178 6151 4181
rect 9029 4178 9095 4181
rect 6085 4176 9095 4178
rect 6085 4120 6090 4176
rect 6146 4120 9034 4176
rect 9090 4120 9095 4176
rect 6085 4118 9095 4120
rect 1669 4115 1735 4118
rect 6085 4115 6151 4118
rect 9029 4115 9095 4118
rect 12525 4178 12591 4181
rect 21633 4178 21699 4181
rect 12525 4176 21699 4178
rect 12525 4120 12530 4176
rect 12586 4120 21638 4176
rect 21694 4120 21699 4176
rect 12525 4118 21699 4120
rect 12525 4115 12591 4118
rect 21633 4115 21699 4118
rect 0 4044 480 4072
rect 0 3980 60 4044
rect 124 3980 480 4044
rect 0 3952 480 3980
rect 2129 4042 2195 4045
rect 4613 4042 4679 4045
rect 9121 4042 9187 4045
rect 2129 4040 9187 4042
rect 2129 3984 2134 4040
rect 2190 3984 4618 4040
rect 4674 3984 9126 4040
rect 9182 3984 9187 4040
rect 2129 3982 9187 3984
rect 2129 3979 2195 3982
rect 4613 3979 4679 3982
rect 9121 3979 9187 3982
rect 29821 4042 29887 4045
rect 39520 4042 40000 4072
rect 29821 4040 40000 4042
rect 29821 3984 29826 4040
rect 29882 3984 40000 4040
rect 29821 3982 40000 3984
rect 29821 3979 29887 3982
rect 39520 3952 40000 3982
rect 4889 3906 4955 3909
rect 7281 3906 7347 3909
rect 4889 3904 7347 3906
rect 4889 3848 4894 3904
rect 4950 3848 7286 3904
rect 7342 3848 7347 3904
rect 4889 3846 7347 3848
rect 4889 3843 4955 3846
rect 7281 3843 7347 3846
rect 18965 3906 19031 3909
rect 24117 3906 24183 3909
rect 18965 3904 24183 3906
rect 18965 3848 18970 3904
rect 19026 3848 24122 3904
rect 24178 3848 24183 3904
rect 18965 3846 24183 3848
rect 18965 3843 19031 3846
rect 24117 3843 24183 3846
rect 14277 3840 14597 3841
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 3775 27930 3776
rect 749 3634 815 3637
rect 62 3632 815 3634
rect 62 3576 754 3632
rect 810 3576 815 3632
rect 62 3574 815 3576
rect 62 3120 122 3574
rect 749 3571 815 3574
rect 13905 3498 13971 3501
rect 14365 3498 14431 3501
rect 19241 3498 19307 3501
rect 13905 3496 19307 3498
rect 13905 3440 13910 3496
rect 13966 3440 14370 3496
rect 14426 3440 19246 3496
rect 19302 3440 19307 3496
rect 13905 3438 19307 3440
rect 13905 3435 13971 3438
rect 14365 3435 14431 3438
rect 19241 3435 19307 3438
rect 23430 3438 39682 3498
rect 23289 3362 23355 3365
rect 23430 3362 23490 3438
rect 23289 3360 23490 3362
rect 23289 3304 23294 3360
rect 23350 3304 23490 3360
rect 23289 3302 23490 3304
rect 23289 3299 23355 3302
rect 25998 3300 26004 3364
rect 26068 3362 26074 3364
rect 26141 3362 26207 3365
rect 26068 3360 26207 3362
rect 26068 3304 26146 3360
rect 26202 3304 26207 3360
rect 26068 3302 26207 3304
rect 26068 3300 26074 3302
rect 26141 3299 26207 3302
rect 7610 3296 7930 3297
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 39622 3120 39682 3438
rect 0 3000 480 3120
rect 6269 3090 6335 3093
rect 17125 3090 17191 3093
rect 6269 3088 17191 3090
rect 6269 3032 6274 3088
rect 6330 3032 17130 3088
rect 17186 3032 17191 3088
rect 6269 3030 17191 3032
rect 6269 3027 6335 3030
rect 17125 3027 17191 3030
rect 18781 3090 18847 3093
rect 30281 3090 30347 3093
rect 18781 3088 30347 3090
rect 18781 3032 18786 3088
rect 18842 3032 30286 3088
rect 30342 3032 30347 3088
rect 18781 3030 30347 3032
rect 18781 3027 18847 3030
rect 30281 3027 30347 3030
rect 39520 3000 40000 3120
rect 19885 2954 19951 2957
rect 27705 2954 27771 2957
rect 30465 2954 30531 2957
rect 19885 2952 27771 2954
rect 19885 2896 19890 2952
rect 19946 2896 27710 2952
rect 27766 2896 27771 2952
rect 19885 2894 27771 2896
rect 19885 2891 19951 2894
rect 27705 2891 27771 2894
rect 28950 2952 30531 2954
rect 28950 2896 30470 2952
rect 30526 2896 30531 2952
rect 28950 2894 30531 2896
rect 12249 2818 12315 2821
rect 12382 2818 12388 2820
rect 12249 2816 12388 2818
rect 12249 2760 12254 2816
rect 12310 2760 12388 2816
rect 12249 2758 12388 2760
rect 12249 2755 12315 2758
rect 12382 2756 12388 2758
rect 12452 2756 12458 2820
rect 20897 2818 20963 2821
rect 23749 2818 23815 2821
rect 20897 2816 23815 2818
rect 20897 2760 20902 2816
rect 20958 2760 23754 2816
rect 23810 2760 23815 2816
rect 20897 2758 23815 2760
rect 20897 2755 20963 2758
rect 23749 2755 23815 2758
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2687 27930 2688
rect 14825 2682 14891 2685
rect 18505 2682 18571 2685
rect 24669 2682 24735 2685
rect 14825 2680 24735 2682
rect 14825 2624 14830 2680
rect 14886 2624 18510 2680
rect 18566 2624 24674 2680
rect 24730 2624 24735 2680
rect 14825 2622 24735 2624
rect 14825 2619 14891 2622
rect 18505 2619 18571 2622
rect 24669 2619 24735 2622
rect 12341 2546 12407 2549
rect 20805 2546 20871 2549
rect 12341 2544 20871 2546
rect 12341 2488 12346 2544
rect 12402 2488 20810 2544
rect 20866 2488 20871 2544
rect 12341 2486 20871 2488
rect 12341 2483 12407 2486
rect 20805 2483 20871 2486
rect 22093 2546 22159 2549
rect 28950 2546 29010 2894
rect 30465 2891 30531 2894
rect 32489 2818 32555 2821
rect 32489 2816 39682 2818
rect 32489 2760 32494 2816
rect 32550 2760 39682 2816
rect 32489 2758 39682 2760
rect 32489 2755 32555 2758
rect 22093 2544 29010 2546
rect 22093 2488 22098 2544
rect 22154 2488 29010 2544
rect 22093 2486 29010 2488
rect 22093 2483 22159 2486
rect 24025 2410 24091 2413
rect 24853 2410 24919 2413
rect 24025 2408 24919 2410
rect 24025 2352 24030 2408
rect 24086 2352 24858 2408
rect 24914 2352 24919 2408
rect 24025 2350 24919 2352
rect 24025 2347 24091 2350
rect 24853 2347 24919 2350
rect 27429 2410 27495 2413
rect 35985 2410 36051 2413
rect 27429 2408 36051 2410
rect 27429 2352 27434 2408
rect 27490 2352 35990 2408
rect 36046 2352 36051 2408
rect 27429 2350 36051 2352
rect 27429 2347 27495 2350
rect 35985 2347 36051 2350
rect 39622 2304 39682 2758
rect 0 2272 480 2304
rect 0 2216 110 2272
rect 166 2216 480 2272
rect 0 2184 480 2216
rect 11973 2274 12039 2277
rect 20621 2274 20687 2277
rect 11973 2272 20687 2274
rect 11973 2216 11978 2272
rect 12034 2216 20626 2272
rect 20682 2216 20687 2272
rect 11973 2214 20687 2216
rect 11973 2211 12039 2214
rect 20621 2211 20687 2214
rect 7610 2208 7930 2209
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 39520 2184 40000 2304
rect 34277 2143 34597 2144
rect 4245 2002 4311 2005
rect 13353 2002 13419 2005
rect 62 2000 13419 2002
rect 62 1944 4250 2000
rect 4306 1944 13358 2000
rect 13414 1944 13419 2000
rect 62 1942 13419 1944
rect 62 1352 122 1942
rect 4245 1939 4311 1942
rect 13353 1939 13419 1942
rect 27245 2002 27311 2005
rect 27245 2000 33150 2002
rect 27245 1944 27250 2000
rect 27306 1944 33150 2000
rect 27245 1942 33150 1944
rect 27245 1939 27311 1942
rect 33090 1866 33150 1942
rect 36905 1866 36971 1869
rect 33090 1864 39682 1866
rect 33090 1808 36910 1864
rect 36966 1808 39682 1864
rect 33090 1806 39682 1808
rect 36905 1803 36971 1806
rect 39622 1352 39682 1806
rect 0 1232 480 1352
rect 13353 1322 13419 1325
rect 27429 1322 27495 1325
rect 13353 1320 27495 1322
rect 13353 1264 13358 1320
rect 13414 1264 27434 1320
rect 27490 1264 27495 1320
rect 13353 1262 27495 1264
rect 13353 1259 13419 1262
rect 27429 1259 27495 1262
rect 28257 1322 28323 1325
rect 35065 1322 35131 1325
rect 28257 1320 35131 1322
rect 28257 1264 28262 1320
rect 28318 1264 35070 1320
rect 35126 1264 35131 1320
rect 28257 1262 35131 1264
rect 28257 1259 28323 1262
rect 35065 1259 35131 1262
rect 39520 1232 40000 1352
rect 4337 1050 4403 1053
rect 62 1048 4403 1050
rect 62 992 4342 1048
rect 4398 992 4403 1048
rect 62 990 4403 992
rect 62 536 122 990
rect 4337 987 4403 990
rect 31845 1050 31911 1053
rect 31845 1048 39682 1050
rect 31845 992 31850 1048
rect 31906 992 39682 1048
rect 31845 990 39682 992
rect 31845 987 31911 990
rect 39622 536 39682 990
rect 0 416 480 536
rect 39520 416 40000 536
rect 1945 370 2011 373
rect 15193 370 15259 373
rect 1945 368 15259 370
rect 1945 312 1950 368
rect 2006 312 15198 368
rect 15254 312 15259 368
rect 1945 310 15259 312
rect 1945 307 2011 310
rect 15193 307 15259 310
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 60 11052 124 11116
rect 39620 11052 39684 11116
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 60 10780 124 10844
rect 39620 10780 39684 10844
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 39620 7516 39684 7580
rect 39620 7244 39684 7308
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 60 5068 124 5132
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 60 4796 124 4860
rect 60 4524 124 4588
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 60 3980 124 4044
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 26004 3300 26068 3364
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 12388 2756 12452 2820
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 59 11116 125 11117
rect 59 11052 60 11116
rect 124 11052 125 11116
rect 59 11051 125 11052
rect 62 10845 122 11051
rect 7610 10912 7931 11936
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 59 10844 125 10845
rect 59 10780 60 10844
rect 124 10780 125 10844
rect 59 10779 125 10780
rect 7610 9824 7931 10848
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 7610 8736 7931 9760
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 7610 6560 7931 7584
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 59 5132 125 5133
rect 59 5068 60 5132
rect 124 5068 125 5132
rect 59 5067 125 5068
rect 62 4861 122 5067
rect 59 4860 125 4861
rect 59 4796 60 4860
rect 124 4796 125 4860
rect 59 4795 125 4796
rect 59 4588 125 4589
rect 59 4524 60 4588
rect 124 4524 125 4588
rect 59 4523 125 4524
rect 62 4045 122 4523
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 59 4044 125 4045
rect 59 3980 60 4044
rect 124 3980 125 4044
rect 59 3979 125 3980
rect 7610 3296 7931 4320
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 7610 2208 7931 3232
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 12390 2821 12450 2942
rect 12387 2820 12453 2821
rect 12387 2756 12388 2820
rect 12452 2756 12453 2820
rect 12387 2755 12453 2756
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 14277 2752 14597 3776
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 10368 27930 11392
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 8192 27930 9216
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 7104 27930 8128
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 26003 3364 26069 3365
rect 26003 3300 26004 3364
rect 26068 3300 26069 3364
rect 26003 3299 26069 3300
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 26006 3178 26066 3299
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 27610 2752 27930 3776
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2128 27930 2688
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 10912 34597 11936
rect 39619 11116 39685 11117
rect 39619 11052 39620 11116
rect 39684 11052 39685 11116
rect 39619 11051 39685 11052
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 9824 34597 10848
rect 39622 10845 39682 11051
rect 39619 10844 39685 10845
rect 39619 10780 39620 10844
rect 39684 10780 39685 10844
rect 39619 10779 39685 10780
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 7648 34597 8672
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 39619 7580 39685 7581
rect 39619 7516 39620 7580
rect 39684 7516 39685 7580
rect 39619 7515 39685 7516
rect 39622 7309 39682 7515
rect 39619 7308 39685 7309
rect 39619 7244 39620 7308
rect 39684 7244 39685 7308
rect 39619 7243 39685 7244
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 5472 34597 6496
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 3296 34597 4320
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 2208 34597 3232
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
<< via4 >>
rect 12302 2942 12538 3178
rect 25918 2942 26154 3178
<< metal5 >>
rect 12260 3178 26196 3220
rect 12260 2942 12302 3178
rect 12538 2942 25918 3178
rect 26154 2942 26196 3178
rect 12260 2900 26196 2942
use scs8hd_decap_3  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__085__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_8 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_11
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _082_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 3312 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_19 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_18
timestamp 1586364061
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_22
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_26
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_31
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_35
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_39 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 406 592
use scs8hd_buf_1  _164_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5060 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_45
timestamp 1586364061
transform 1 0 5244 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_56
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_66
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 7360 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _067_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7084 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _069_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 866 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__C
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_74
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_78
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_70
timestamp 1586364061
transform 1 0 7544 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_80
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _177_
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _178_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_97
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_105
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_129
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_130
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 314 592
use scs8hd_inv_8  _108_
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use scs8hd_or4_4  _110_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_139
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 406 592
use scs8hd_inv_8  _073_
timestamp 1586364061
transform 1 0 15548 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _075_
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_166
timestamp 1586364061
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_158
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_164
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _093_
timestamp 1586364061
transform 1 0 17112 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__075__C
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__D
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_170
timestamp 1586364061
transform 1 0 16744 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_177
timestamp 1586364061
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_181
timestamp 1586364061
transform 1 0 17756 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 17940 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_buf_1  _076_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_187
timestamp 1586364061
transform 1 0 18308 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_185
timestamp 1586364061
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 18492 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _148_
timestamp 1586364061
transform 1 0 18492 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_191
timestamp 1586364061
transform 1 0 18676 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_192
timestamp 1586364061
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 18952 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_206
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20792 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__C
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_221
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_225
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_225
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_229
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_229
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__C
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23644 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_256
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_260
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_268
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_264
timestamp 1586364061
transform 1 0 25392 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 -1 2720
box -38 -48 222 592
use scs8hd_conb_1  _190_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25668 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_270
timestamp 1586364061
transform 1 0 25944 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26496 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26128 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26036 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26220 0 1 2720
box -38 -48 866 592
use scs8hd_fill_1  FILLER_0_278
timestamp 1586364061
transform 1 0 26680 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_286
timestamp 1586364061
transform 1 0 27416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_282
timestamp 1586364061
transform 1 0 27048 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_283
timestamp 1586364061
transform 1 0 27140 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27232 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27324 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_287
timestamp 1586364061
transform 1 0 27508 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27600 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _146_
timestamp 1586364061
transform 1 0 27784 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_293
timestamp 1586364061
transform 1 0 28060 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_294
timestamp 1586364061
transform 1 0 28152 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 28244 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27876 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_297
timestamp 1586364061
transform 1 0 28428 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_298
timestamp 1586364061
transform 1 0 28520 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28336 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 28612 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_301
timestamp 1586364061
transform 1 0 28796 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_302
timestamp 1586364061
transform 1 0 28888 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 28980 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_309
timestamp 1586364061
transform 1 0 29532 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_305
timestamp 1586364061
transform 1 0 29164 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29348 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_316
timestamp 1586364061
transform 1 0 30176 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29348 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _161_
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 866 592
use scs8hd_conb_1  _191_
timestamp 1586364061
transform 1 0 30912 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31280 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30728 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_320 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 30544 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_331
timestamp 1586364061
transform 1 0 31556 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_320
timestamp 1586364061
transform 1 0 30544 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_327
timestamp 1586364061
transform 1 0 31188 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31740 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_339
timestamp 1586364061
transform 1 0 32292 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_354
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_351
timestamp 1586364061
transform 1 0 33396 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_363
timestamp 1586364061
transform 1 0 34500 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2668 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_35
timestamp 1586364061
transform 1 0 4324 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_46
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_2_52
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_1  _084_
timestamp 1586364061
transform 1 0 6348 0 -1 3808
box -38 -48 314 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__C
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_77
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_81
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 590 592
use scs8hd_nor2_4  _176_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_87
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_90
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 590 592
use scs8hd_inv_8  _068_
timestamp 1586364061
transform 1 0 11500 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_112
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_122
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 222 592
use scs8hd_nand2_4  _109_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_126
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_130
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_151
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _094_
timestamp 1586364061
transform 1 0 16008 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_158
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__C
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_171
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_175
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 406 592
use scs8hd_or4_4  _137_
timestamp 1586364061
transform 1 0 17756 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__C
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use scs8hd_or2_4  _145_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19320 0 -1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 19136 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_194
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_nor3_4  _156_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 22264 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 22632 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_232
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 222 592
use scs8hd_nor3_4  _158_
timestamp 1586364061
transform 1 0 22816 0 -1 3808
box -38 -48 1234 592
use scs8hd_fill_2  FILLER_2_249
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _159_
timestamp 1586364061
transform 1 0 24748 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_253
timestamp 1586364061
transform 1 0 24380 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_266
timestamp 1586364061
transform 1 0 25576 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_272
timestamp 1586364061
transform 1 0 26128 0 -1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 27692 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26956 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_279
timestamp 1586364061
transform 1 0 26772 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_283
timestamp 1586364061
transform 1 0 27140 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_8  FILLER_2_300
timestamp 1586364061
transform 1 0 28704 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29440 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_12  FILLER_2_317
timestamp 1586364061
transform 1 0 30268 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_2_329
timestamp 1586364061
transform 1 0 31372 0 -1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_335
timestamp 1586364061
transform 1 0 31924 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_337
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_349
timestamp 1586364061
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_361
timestamp 1586364061
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_373
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_385
timestamp 1586364061
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_17
timestamp 1586364061
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_21
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _081_
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__C
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_42
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_46
timestamp 1586364061
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_75
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _179_
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__C
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_88
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_92
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_109
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _174_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_113
timestamp 1586364061
transform 1 0 11500 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _074_
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_146
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 130 592
use scs8hd_or4_4  _095_
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_158
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_162
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _119_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_or4_4  _147_
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__C
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__D
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_210
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_214
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_219
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use scs8hd_nor3_4  _155_
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 23920 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_236
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 24288 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_250
timestamp 1586364061
transform 1 0 24104 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26220 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 25668 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26036 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_265
timestamp 1586364061
transform 1 0 25484 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _130_
timestamp 1586364061
transform 1 0 27784 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 27600 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 27232 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_282
timestamp 1586364061
transform 1 0 27048 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_286
timestamp 1586364061
transform 1 0 27416 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 28244 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 28612 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_293
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_297
timestamp 1586364061
transform 1 0 28428 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_301
timestamp 1586364061
transform 1 0 28796 0 1 3808
box -38 -48 406 592
use scs8hd_buf_1  _120_
timestamp 1586364061
transform 1 0 30268 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30084 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_309
timestamp 1586364061
transform 1 0 29532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_313
timestamp 1586364061
transform 1 0 29900 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 30728 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_320
timestamp 1586364061
transform 1 0 30544 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_324
timestamp 1586364061
transform 1 0 30912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_336
timestamp 1586364061
transform 1 0 32016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_348
timestamp 1586364061
transform 1 0 33120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_360
timestamp 1586364061
transform 1 0 34224 0 1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_379
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_391
timestamp 1586364061
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_4  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 590 592
use scs8hd_or3_4  _098_
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use scs8hd_or3_4  _090_
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_58
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_75
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_81
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_or3_4  _080_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_85
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_89
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 774 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_114
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_128
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_132
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_or2_4  _171_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_161
timestamp 1586364061
transform 1 0 15916 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_165
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 130 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_1  FILLER_4_168
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_182
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_1  _078_
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_195
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_199
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_218
timestamp 1586364061
transform 1 0 21160 0 -1 4896
box -38 -48 406 592
use scs8hd_nor3_4  _157_
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 21620 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_222
timestamp 1586364061
transform 1 0 21528 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_225
timestamp 1586364061
transform 1 0 21804 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_241
timestamp 1586364061
transform 1 0 23276 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_6  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 590 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 24748 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24472 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_253
timestamp 1586364061
transform 1 0 24380 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_256
timestamp 1586364061
transform 1 0 24656 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_8  _162_
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 25760 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_266
timestamp 1586364061
transform 1 0 25576 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_270
timestamp 1586364061
transform 1 0 25944 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27508 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_285
timestamp 1586364061
transform 1 0 27324 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_289
timestamp 1586364061
transform 1 0 27692 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 28060 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_302
timestamp 1586364061
transform 1 0 28888 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29624 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 30084 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_313
timestamp 1586364061
transform 1 0 29900 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_317
timestamp 1586364061
transform 1 0 30268 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_4_329
timestamp 1586364061
transform 1 0 31372 0 -1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_335
timestamp 1586364061
transform 1 0 31924 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_373
timestamp 1586364061
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_385
timestamp 1586364061
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_16
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_20
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_24
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3680 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _070_
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_43
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_47
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _099_
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_68
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_72
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_139
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _173_
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_160
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_177
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use scs8hd_or2_4  _072_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_191
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _160_
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_212
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_217
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_228
timestamp 1586364061
transform 1 0 22080 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_234
timestamp 1586364061
transform 1 0 22632 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_238
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_242
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 26220 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_271
timestamp 1586364061
transform 1 0 26036 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_275
timestamp 1586364061
transform 1 0 26404 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27048 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26864 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_279
timestamp 1586364061
transform 1 0 26772 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28520 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28888 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28060 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_291
timestamp 1586364061
transform 1 0 27876 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_295
timestamp 1586364061
transform 1 0 28244 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_300
timestamp 1586364061
transform 1 0 28704 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_304
timestamp 1586364061
transform 1 0 29072 0 1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30268 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 30084 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_309
timestamp 1586364061
transform 1 0 29532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_313
timestamp 1586364061
transform 1 0 29900 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31280 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30728 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_320
timestamp 1586364061
transform 1 0 30544 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_324
timestamp 1586364061
transform 1 0 30912 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_331
timestamp 1586364061
transform 1 0 31556 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32108 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31740 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_335
timestamp 1586364061
transform 1 0 31924 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_339
timestamp 1586364061
transform 1 0 32292 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33396 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34040 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_353
timestamp 1586364061
transform 1 0 33580 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_357
timestamp 1586364061
transform 1 0 33948 0 1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35328 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34408 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_360
timestamp 1586364061
transform 1 0 34224 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_364
timestamp 1586364061
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_370
timestamp 1586364061
transform 1 0 35144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_374
timestamp 1586364061
transform 1 0 35512 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_378
timestamp 1586364061
transform 1 0 35880 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_381
timestamp 1586364061
transform 1 0 36156 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_393
timestamp 1586364061
transform 1 0 37260 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_405
timestamp 1586364061
transform 1 0 38364 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _200_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_17
timestamp 1586364061
transform 1 0 2668 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_21
timestamp 1586364061
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_25
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_26
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_29
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_30
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_43
timestamp 1586364061
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_47
timestamp 1586364061
transform 1 0 5428 0 1 5984
box -38 -48 774 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_58
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_62
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _167_
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_75
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_81
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_85
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_88
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_92
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_104
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_108
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_116
timestamp 1586364061
transform 1 0 11776 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_113
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_117
timestamp 1586364061
transform 1 0 11868 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_120
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_128
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_132
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _071_
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_145
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_149
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__D
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_166
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_168
timestamp 1586364061
transform 1 0 16560 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_170
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_178
timestamp 1586364061
transform 1 0 17480 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_181
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_184
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_180
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 18216 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_201
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_201
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_209
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_216
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_229
timestamp 1586364061
transform 1 0 22172 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_6_234
timestamp 1586364061
transform 1 0 22632 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_224
timestamp 1586364061
transform 1 0 21712 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 23184 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_or2_4  _129_
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24380 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_255
timestamp 1586364061
transform 1 0 24564 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_256
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_260
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_265
timestamp 1586364061
transform 1 0 25484 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_266
timestamp 1586364061
transform 1 0 25576 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25852 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 25668 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_271
timestamp 1586364061
transform 1 0 26036 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26956 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27416 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27048 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26772 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_290
timestamp 1586364061
transform 1 0 27784 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_280
timestamp 1586364061
transform 1 0 26864 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_284
timestamp 1586364061
transform 1 0 27232 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28520 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27968 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_294
timestamp 1586364061
transform 1 0 28152 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_297
timestamp 1586364061
transform 1 0 28428 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_301
timestamp 1586364061
transform 1 0 28796 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 30084 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29532 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_307
timestamp 1586364061
transform 1 0 29348 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_311
timestamp 1586364061
transform 1 0 29716 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_315
timestamp 1586364061
transform 1 0 30084 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 31096 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 30452 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 30912 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 31096 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_324
timestamp 1586364061
transform 1 0 30912 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_328
timestamp 1586364061
transform 1 0 31280 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_321
timestamp 1586364061
transform 1 0 30636 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_339
timestamp 1586364061
transform 1 0 32292 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_335
timestamp 1586364061
transform 1 0 31924 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 32108 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_6_345
timestamp 1586364061
transform 1 0 32844 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_3  FILLER_6_340
timestamp 1586364061
transform 1 0 32384 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32660 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 32476 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 32660 0 1 5984
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33396 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33856 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_354
timestamp 1586364061
transform 1 0 33672 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_354
timestamp 1586364061
transform 1 0 33672 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_358
timestamp 1586364061
transform 1 0 34040 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34408 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34224 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_371
timestamp 1586364061
transform 1 0 35236 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_362
timestamp 1586364061
transform 1 0 34408 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_376
timestamp 1586364061
transform 1 0 35696 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_375
timestamp 1586364061
transform 1 0 35604 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35972 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35972 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_387
timestamp 1586364061
transform 1 0 36708 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_381
timestamp 1586364061
transform 1 0 36156 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_382
timestamp 1586364061
transform 1 0 36248 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36432 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36432 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_386
timestamp 1586364061
transform 1 0 36616 0 -1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36892 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_394
timestamp 1586364061
transform 1 0 37352 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_391
timestamp 1586364061
transform 1 0 37076 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_403
timestamp 1586364061
transform 1 0 38180 0 1 5984
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_9
timestamp 1586364061
transform 1 0 1932 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 314 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_70
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_8_75
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_104
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_8_116
timestamp 1586364061
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_135
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 130 592
use scs8hd_or2_4  _077_
timestamp 1586364061
transform 1 0 17572 0 -1 7072
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_170
timestamp 1586364061
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_174
timestamp 1586364061
transform 1 0 17112 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18768 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_8_205
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_211
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_228
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_235
timestamp 1586364061
transform 1 0 22724 0 -1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 23736 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  FILLER_8_243
timestamp 1586364061
transform 1 0 23460 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_255
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25852 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_266
timestamp 1586364061
transform 1 0 25576 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_271
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27048 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26680 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_280
timestamp 1586364061
transform 1 0 26864 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28612 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28428 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_291
timestamp 1586364061
transform 1 0 27876 0 -1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 30268 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_308
timestamp 1586364061
transform 1 0 29440 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_316
timestamp 1586364061
transform 1 0 30176 0 -1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 30452 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_328
timestamp 1586364061
transform 1 0 31280 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33488 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33856 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_348
timestamp 1586364061
transform 1 0 33120 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_354
timestamp 1586364061
transform 1 0 33672 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_358
timestamp 1586364061
transform 1 0 34040 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34408 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_371
timestamp 1586364061
transform 1 0 35236 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35972 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_4  FILLER_8_375
timestamp 1586364061
transform 1 0 35604 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_388
timestamp 1586364061
transform 1 0 36800 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_396
timestamp 1586364061
transform 1 0 37536 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_9_9
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 5612 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_44
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_48
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 406 592
use scs8hd_buf_1  _091_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_65
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_69
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_84
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_90
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_107
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_111
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_117
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_121
timestamp 1586364061
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_131
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_144
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_148
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_155
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_199
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_210
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_214
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_218
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 22632 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_262
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 25668 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_266
timestamp 1586364061
transform 1 0 25576 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 27048 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27416 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_280
timestamp 1586364061
transform 1 0 26864 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_284
timestamp 1586364061
transform 1 0 27232 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 28888 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_297
timestamp 1586364061
transform 1 0 28428 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_301
timestamp 1586364061
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_304
timestamp 1586364061
transform 1 0 29072 0 1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 30084 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 29900 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29440 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_306
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_310
timestamp 1586364061
transform 1 0 29624 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_326
timestamp 1586364061
transform 1 0 31096 0 1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32200 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32660 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_341
timestamp 1586364061
transform 1 0 32476 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_345
timestamp 1586364061
transform 1 0 32844 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_358
timestamp 1586364061
transform 1 0 34040 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 34224 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_362
timestamp 1586364061
transform 1 0 34408 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 36432 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_376
timestamp 1586364061
transform 1 0 35696 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_380
timestamp 1586364061
transform 1 0 36064 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 36984 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_388
timestamp 1586364061
transform 1 0 36800 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_392
timestamp 1586364061
transform 1 0 37168 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_404
timestamp 1586364061
transform 1 0 38272 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_18
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_22
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_53
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_57
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_60
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_73
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_4  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_99
timestamp 1586364061
transform 1 0 10212 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_111
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_128
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_132
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_165
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_169
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_173
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_177
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_187
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_191
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_204
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_208
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_4  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_230
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 774 592
use scs8hd_or2_4  _121_
timestamp 1586364061
transform 1 0 23000 0 -1 8160
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_245
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_249
timestamp 1586364061
transform 1 0 24012 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 24472 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_253
timestamp 1586364061
transform 1 0 24380 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_265
timestamp 1586364061
transform 1 0 25484 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_269
timestamp 1586364061
transform 1 0 25852 0 -1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27692 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_287
timestamp 1586364061
transform 1 0 27508 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 28888 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_10_291
timestamp 1586364061
transform 1 0 27876 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_299
timestamp 1586364061
transform 1 0 28612 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30084 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_313
timestamp 1586364061
transform 1 0 29900 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_317
timestamp 1586364061
transform 1 0 30268 0 -1 8160
box -38 -48 222 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 30636 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 30452 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_324
timestamp 1586364061
transform 1 0 30912 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32476 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 32292 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_344
timestamp 1586364061
transform 1 0 32752 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 33488 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33212 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_348
timestamp 1586364061
transform 1 0 33120 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_351
timestamp 1586364061
transform 1 0 33396 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35236 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_363
timestamp 1586364061
transform 1 0 34500 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_369
timestamp 1586364061
transform 1 0 35052 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_380
timestamp 1586364061
transform 1 0 36064 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_392
timestamp 1586364061
transform 1 0 37168 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_396
timestamp 1586364061
transform 1 0 37536 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_21
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_25
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_37
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_41
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6900 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_78
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_82
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_89
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_108
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_116
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_157
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_161
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 19688 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_194
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_198
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_213
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_230
timestamp 1586364061
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_234
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_238
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_256
timestamp 1586364061
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_260
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_264
timestamp 1586364061
transform 1 0 25392 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_276
timestamp 1586364061
transform 1 0 26496 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 27600 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 27416 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 26680 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 27048 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_280
timestamp 1586364061
transform 1 0 26864 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_284
timestamp 1586364061
transform 1 0 27232 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_297
timestamp 1586364061
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_301
timestamp 1586364061
transform 1 0 28796 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29992 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29808 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31556 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 31004 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31372 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_323
timestamp 1586364061
transform 1 0 30820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_327
timestamp 1586364061
transform 1 0 31188 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 32752 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 32568 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 32108 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_334
timestamp 1586364061
transform 1 0 31832 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_339
timestamp 1586364061
transform 1 0 32292 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 33948 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_355
timestamp 1586364061
transform 1 0 33764 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_359
timestamp 1586364061
transform 1 0 34132 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_363
timestamp 1586364061
transform 1 0 34500 0 1 8160
box -38 -48 130 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 36432 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 35880 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_376
timestamp 1586364061
transform 1 0 35696 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_380
timestamp 1586364061
transform 1 0 36064 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 36984 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_388
timestamp 1586364061
transform 1 0 36800 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_392
timestamp 1586364061
transform 1 0 37168 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_404
timestamp 1586364061
transform 1 0 38272 0 1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_38
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_50
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_67
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_12_71
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_96
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_100
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_104
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_119
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_133
timestamp 1586364061
transform 1 0 13340 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15732 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_158
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_170
timestamp 1586364061
transform 1 0 16744 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_181
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_185
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_189
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 19872 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 590 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_218
timestamp 1586364061
transform 1 0 21160 0 -1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 22264 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21804 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_223
timestamp 1586364061
transform 1 0 21620 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_258
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_262
timestamp 1586364061
transform 1 0 25208 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25392 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_266
timestamp 1586364061
transform 1 0 25576 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_272
timestamp 1586364061
transform 1 0 26128 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 27600 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_285
timestamp 1586364061
transform 1 0 27324 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_12_290
timestamp 1586364061
transform 1 0 27784 0 -1 9248
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 28612 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28428 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_296
timestamp 1586364061
transform 1 0 28336 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29992 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_310
timestamp 1586364061
transform 1 0 29624 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_12_316
timestamp 1586364061
transform 1 0 30176 0 -1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 30452 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_328
timestamp 1586364061
transform 1 0 31280 0 -1 9248
box -38 -48 774 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 33672 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33120 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33488 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_346
timestamp 1586364061
transform 1 0 32936 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_350
timestamp 1586364061
transform 1 0 33304 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 35420 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35236 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_365
timestamp 1586364061
transform 1 0 34684 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_369
timestamp 1586364061
transform 1 0 35052 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36616 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_384
timestamp 1586364061
transform 1 0 36432 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_388
timestamp 1586364061
transform 1 0 36800 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_396
timestamp 1586364061
transform 1 0 37536 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_21
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_25
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_18
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 1142 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_29
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_30
timestamp 1586364061
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_42
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_46
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_43
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_55
timestamp 1586364061
transform 1 0 6164 0 -1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _180_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_62
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_73
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_90
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_94
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_109
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_110
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_127
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_135
timestamp 1586364061
transform 1 0 13524 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_162
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_166
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_158
timestamp 1586364061
transform 1 0 15640 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _175_
timestamp 1586364061
transform 1 0 17572 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_169
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_177
timestamp 1586364061
transform 1 0 17388 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_188
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_189
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_192
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_212
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_209
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_227
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_231
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_236
timestamp 1586364061
transform 1 0 22816 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_248
timestamp 1586364061
transform 1 0 23920 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24656 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24472 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_256
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_260
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_252
timestamp 1586364061
transform 1 0 24288 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25392 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 26036 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_273
timestamp 1586364061
transform 1 0 26220 0 1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_265
timestamp 1586364061
transform 1 0 25484 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_273
timestamp 1586364061
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 27600 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 27416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 27784 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 27048 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_278
timestamp 1586364061
transform 1 0 26680 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_284
timestamp 1586364061
transform 1 0 27232 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_285
timestamp 1586364061
transform 1 0 27324 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_289
timestamp 1586364061
transform 1 0 27692 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 28520 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_297
timestamp 1586364061
transform 1 0 28428 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_301
timestamp 1586364061
transform 1 0 28796 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_292
timestamp 1586364061
transform 1 0 27968 0 -1 10336
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30360 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29716 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30084 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_317
timestamp 1586364061
transform 1 0 30268 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_309
timestamp 1586364061
transform 1 0 29532 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_313
timestamp 1586364061
transform 1 0 29900 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_317
timestamp 1586364061
transform 1 0 30268 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31280 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30452 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31464 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30820 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_321
timestamp 1586364061
transform 1 0 30636 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_325
timestamp 1586364061
transform 1 0 31004 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_331
timestamp 1586364061
transform 1 0 31556 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_327
timestamp 1586364061
transform 1 0 31188 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_332
timestamp 1586364061
transform 1 0 31648 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_335
timestamp 1586364061
transform 1 0 31924 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 32292 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 32108 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31740 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_345
timestamp 1586364061
transform 1 0 32844 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_341
timestamp 1586364061
transform 1 0 32476 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32660 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 32292 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32936 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33488 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33856 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33948 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_350
timestamp 1586364061
transform 1 0 33304 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_354
timestamp 1586364061
transform 1 0 33672 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_358
timestamp 1586364061
transform 1 0 34040 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_355
timestamp 1586364061
transform 1 0 33764 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_359
timestamp 1586364061
transform 1 0 34132 0 -1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34500 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_362
timestamp 1586364061
transform 1 0 34408 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_372
timestamp 1586364061
transform 1 0 35328 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 36064 0 -1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 36064 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36616 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_376
timestamp 1586364061
transform 1 0 35696 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_382
timestamp 1586364061
transform 1 0 36248 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_384
timestamp 1586364061
transform 1 0 36432 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_393
timestamp 1586364061
transform 1 0 37260 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_388
timestamp 1586364061
transform 1 0 36800 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_396
timestamp 1586364061
transform 1 0 37536 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_405
timestamp 1586364061
transform 1 0 38364 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_18
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_22
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_26
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_33
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_37
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_41
timestamp 1586364061
transform 1 0 4876 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 774 592
use scs8hd_conb_1  _181_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_65
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 774 592
use scs8hd_buf_1  _104_
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_73
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_79
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_83
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_90
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_94
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_15_107
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 406 592
use scs8hd_conb_1  _182_
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 590 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_201
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_214
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_218
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _138_
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_225
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_250
timestamp 1586364061
transform 1 0 24104 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 26036 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_267
timestamp 1586364061
transform 1 0 25668 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 27600 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 27416 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27048 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_280
timestamp 1586364061
transform 1 0 26864 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_284
timestamp 1586364061
transform 1 0 27232 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 28612 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_297
timestamp 1586364061
transform 1 0 28428 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_301
timestamp 1586364061
transform 1 0 28796 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29900 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29716 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_310
timestamp 1586364061
transform 1 0 29624 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31464 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 31280 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30912 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_322
timestamp 1586364061
transform 1 0 30728 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_326
timestamp 1586364061
transform 1 0 31096 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 32844 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 32476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_339
timestamp 1586364061
transform 1 0 32292 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_343
timestamp 1586364061
transform 1 0 32660 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 33028 0 1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_15_356
timestamp 1586364061
transform 1 0 33856 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 34316 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_360
timestamp 1586364061
transform 1 0 34224 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_363
timestamp 1586364061
transform 1 0 34500 0 1 10336
box -38 -48 314 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 36432 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 35880 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 36248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_376
timestamp 1586364061
transform 1 0 35696 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_380
timestamp 1586364061
transform 1 0 36064 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37536 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 36984 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37996 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_388
timestamp 1586364061
transform 1 0 36800 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_392
timestamp 1586364061
transform 1 0 37168 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_399
timestamp 1586364061
transform 1 0 37812 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_403
timestamp 1586364061
transform 1 0 38180 0 1 10336
box -38 -48 406 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 774 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_35
timestamp 1586364061
transform 1 0 4324 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_47
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_59
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_71
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_79
timestamp 1586364061
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_104
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_108
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_121
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _113_
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_132
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_165
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_177
timestamp 1586364061
transform 1 0 17388 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_188
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 19136 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_205
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_209
timestamp 1586364061
transform 1 0 20332 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_236
timestamp 1586364061
transform 1 0 22816 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_240
timestamp 1586364061
transform 1 0 23184 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_244
timestamp 1586364061
transform 1 0 23552 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24288 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_12  FILLER_16_261
timestamp 1586364061
transform 1 0 25116 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_273
timestamp 1586364061
transform 1 0 26220 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 27784 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 27600 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_279
timestamp 1586364061
transform 1 0 26772 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_287
timestamp 1586364061
transform 1 0 27508 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_299
timestamp 1586364061
transform 1 0 28612 0 -1 11424
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29716 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31464 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_320
timestamp 1586364061
transform 1 0 30544 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_328
timestamp 1586364061
transform 1 0 31280 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_332
timestamp 1586364061
transform 1 0 31648 0 -1 11424
box -38 -48 406 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_346
timestamp 1586364061
transform 1 0 32936 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_16_358
timestamp 1586364061
transform 1 0 34040 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 406 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 34316 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34868 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35236 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_365
timestamp 1586364061
transform 1 0 34684 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_369
timestamp 1586364061
transform 1 0 35052 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 36524 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_377
timestamp 1586364061
transform 1 0 35788 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_389
timestamp 1586364061
transform 1 0 36892 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_18
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_22
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_26
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_38
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_50
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_58
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_17_94
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 774 592
use scs8hd_conb_1  _184_
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_155
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_161
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_173
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 774 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 18584 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _185_
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_205
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_216
timestamp 1586364061
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24012 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24380 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_251
timestamp 1586364061
transform 1 0 24196 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_256
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_260
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _186_
timestamp 1586364061
transform 1 0 25392 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_267
timestamp 1586364061
transform 1 0 25668 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_279
timestamp 1586364061
transform 1 0 26772 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_291
timestamp 1586364061
transform 1 0 27876 0 1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_17_303
timestamp 1586364061
transform 1 0 28980 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29992 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_317
timestamp 1586364061
transform 1 0 30268 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31188 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31648 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30452 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_321
timestamp 1586364061
transform 1 0 30636 0 1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_17_330
timestamp 1586364061
transform 1 0 31464 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_334
timestamp 1586364061
transform 1 0 31832 0 1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_346
timestamp 1586364061
transform 1 0 32936 0 1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_17_354
timestamp 1586364061
transform 1 0 33672 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_358
timestamp 1586364061
transform 1 0 34040 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 35420 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 35236 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_362
timestamp 1586364061
transform 1 0 34408 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36524 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_377
timestamp 1586364061
transform 1 0 35788 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_381
timestamp 1586364061
transform 1 0 36156 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36984 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_388
timestamp 1586364061
transform 1 0 36800 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_392
timestamp 1586364061
transform 1 0 37168 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_404
timestamp 1586364061
transform 1 0 38272 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_9
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2668 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_20
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_28
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_99
timestamp 1586364061
transform 1 0 10212 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_110
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_122
timestamp 1586364061
transform 1 0 12328 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_134
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_18_146
timestamp 1586364061
transform 1 0 14536 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 590 592
use scs8hd_buf_1  _172_
timestamp 1586364061
transform 1 0 19136 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_199
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_211
timestamp 1586364061
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_247
timestamp 1586364061
transform 1 0 23828 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_252
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_288
timestamp 1586364061
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_300
timestamp 1586364061
transform 1 0 28704 0 -1 12512
box -38 -48 774 592
use scs8hd_conb_1  _188_
timestamp 1586364061
transform 1 0 29532 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_308
timestamp 1586364061
transform 1 0 29440 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_312
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_324
timestamp 1586364061
transform 1 0 30912 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_349
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34316 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_364
timestamp 1586364061
transform 1 0 34592 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_372
timestamp 1586364061
transform 1 0 35328 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_377
timestamp 1586364061
transform 1 0 35788 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_389
timestamp 1586364061
transform 1 0 36892 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 590 592
use scs8hd_decap_6  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24196 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_254
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_258
timestamp 1586364061
transform 1 0 24840 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_261
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_270
timestamp 1586364061
transform 1 0 25944 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_282
timestamp 1586364061
transform 1 0 27048 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_280
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_294
timestamp 1586364061
transform 1 0 28152 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_302
timestamp 1586364061
transform 1 0 28888 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_292
timestamp 1586364061
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_304
timestamp 1586364061
transform 1 0 29072 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_330
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_323
timestamp 1586364061
transform 1 0 30820 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_342
timestamp 1586364061
transform 1 0 32568 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_354
timestamp 1586364061
transform 1 0 33672 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_354
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_366
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_379
timestamp 1586364061
transform 1 0 35972 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_385
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_391
timestamp 1586364061
transform 1 0 37076 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_397
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_403
timestamp 1586364061
transform 1 0 38180 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal2 s 4986 0 5042 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 8298 0 8354 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 11610 0 11666 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 15014 0 15070 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 18326 0 18382 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 21638 0 21694 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 24950 0 25006 480 6 address[6]
port 6 nsew default input
rlabel metal2 s 31666 0 31722 480 6 bottom_grid_pin_0_
port 7 nsew default tristate
rlabel metal2 s 34978 0 35034 480 6 bottom_grid_pin_4_
port 8 nsew default tristate
rlabel metal2 s 38290 0 38346 480 6 bottom_grid_pin_8_
port 9 nsew default tristate
rlabel metal3 s 0 416 480 536 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal3 s 0 1232 480 1352 6 chanx_left_in[1]
port 11 nsew default input
rlabel metal3 s 0 2184 480 2304 6 chanx_left_in[2]
port 12 nsew default input
rlabel metal3 s 0 3000 480 3120 6 chanx_left_in[3]
port 13 nsew default input
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[4]
port 14 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[5]
port 15 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[6]
port 16 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[7]
port 17 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[8]
port 18 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_out[0]
port 19 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[1]
port 20 nsew default tristate
rlabel metal3 s 0 10208 480 10328 6 chanx_left_out[2]
port 21 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[3]
port 22 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 chanx_left_out[4]
port 23 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 chanx_left_out[5]
port 24 nsew default tristate
rlabel metal3 s 0 13744 480 13864 6 chanx_left_out[6]
port 25 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[7]
port 26 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[8]
port 27 nsew default tristate
rlabel metal3 s 39520 416 40000 536 6 chanx_right_in[0]
port 28 nsew default input
rlabel metal3 s 39520 1232 40000 1352 6 chanx_right_in[1]
port 29 nsew default input
rlabel metal3 s 39520 2184 40000 2304 6 chanx_right_in[2]
port 30 nsew default input
rlabel metal3 s 39520 3000 40000 3120 6 chanx_right_in[3]
port 31 nsew default input
rlabel metal3 s 39520 3952 40000 4072 6 chanx_right_in[4]
port 32 nsew default input
rlabel metal3 s 39520 4768 40000 4888 6 chanx_right_in[5]
port 33 nsew default input
rlabel metal3 s 39520 5720 40000 5840 6 chanx_right_in[6]
port 34 nsew default input
rlabel metal3 s 39520 6536 40000 6656 6 chanx_right_in[7]
port 35 nsew default input
rlabel metal3 s 39520 7488 40000 7608 6 chanx_right_in[8]
port 36 nsew default input
rlabel metal3 s 39520 8440 40000 8560 6 chanx_right_out[0]
port 37 nsew default tristate
rlabel metal3 s 39520 9256 40000 9376 6 chanx_right_out[1]
port 38 nsew default tristate
rlabel metal3 s 39520 10208 40000 10328 6 chanx_right_out[2]
port 39 nsew default tristate
rlabel metal3 s 39520 11024 40000 11144 6 chanx_right_out[3]
port 40 nsew default tristate
rlabel metal3 s 39520 11976 40000 12096 6 chanx_right_out[4]
port 41 nsew default tristate
rlabel metal3 s 39520 12792 40000 12912 6 chanx_right_out[5]
port 42 nsew default tristate
rlabel metal3 s 39520 13744 40000 13864 6 chanx_right_out[6]
port 43 nsew default tristate
rlabel metal3 s 39520 14560 40000 14680 6 chanx_right_out[7]
port 44 nsew default tristate
rlabel metal3 s 39520 15512 40000 15632 6 chanx_right_out[8]
port 45 nsew default tristate
rlabel metal2 s 28354 0 28410 480 6 data_in
port 46 nsew default input
rlabel metal2 s 1674 0 1730 480 6 enable
port 47 nsew default input
rlabel metal2 s 2502 15520 2558 16000 6 top_grid_pin_0_
port 48 nsew default tristate
rlabel metal2 s 27434 15520 27490 16000 6 top_grid_pin_10_
port 49 nsew default tristate
rlabel metal2 s 32494 15520 32550 16000 6 top_grid_pin_12_
port 50 nsew default tristate
rlabel metal2 s 37462 15520 37518 16000 6 top_grid_pin_14_
port 51 nsew default tristate
rlabel metal2 s 7470 15520 7526 16000 6 top_grid_pin_2_
port 52 nsew default tristate
rlabel metal2 s 12438 15520 12494 16000 6 top_grid_pin_4_
port 53 nsew default tristate
rlabel metal2 s 17498 15520 17554 16000 6 top_grid_pin_6_
port 54 nsew default tristate
rlabel metal2 s 22466 15520 22522 16000 6 top_grid_pin_8_
port 55 nsew default tristate
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 56 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 57 nsew default input
<< end >>
