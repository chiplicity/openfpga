magic
tech EFS8A
magscale 1 2
timestamp 1604399383
<< locali >>
rect 2697 26095 2731 26537
rect 11471 26061 11839 26095
rect 16715 26061 16807 26095
rect 11805 25891 11839 26061
rect 15393 25687 15427 25789
rect 16773 25687 16807 26061
rect 16865 25959 16899 26129
rect 19349 25959 19383 26333
rect 14565 25279 14599 25449
rect 17601 25143 17635 25313
rect 21557 25143 21591 25245
rect 19349 21947 19383 22185
rect 20453 21879 20487 22117
rect 20913 21879 20947 22185
rect 12081 20315 12115 20485
rect 19441 19771 19475 19873
rect 24685 19703 24719 19873
rect 3249 16439 3283 16745
rect 8861 15351 8895 15453
rect 18889 14875 18923 15045
rect 2421 13719 2455 14025
rect 19073 13787 19107 14025
rect 19165 13855 19199 13957
rect 23213 12631 23247 12869
rect 6285 12155 6319 12257
rect 22477 10455 22511 10761
rect 22385 9367 22419 9537
rect 22201 8823 22235 8925
rect 22143 8789 22235 8823
rect 18613 7735 18647 7973
rect 19901 6647 19935 6885
rect 3249 5559 3283 5661
rect 24869 4063 24903 4233
rect 3249 2839 3283 2941
<< viali >>
rect 2697 26537 2731 26571
rect 19349 26333 19383 26367
rect 16865 26129 16899 26163
rect 2697 26061 2731 26095
rect 11437 26061 11471 26095
rect 16681 26061 16715 26095
rect 11805 25857 11839 25891
rect 15393 25789 15427 25823
rect 15393 25653 15427 25687
rect 16865 25925 16899 25959
rect 19349 25925 19383 25959
rect 16773 25653 16807 25687
rect 9965 25449 9999 25483
rect 14381 25449 14415 25483
rect 14565 25449 14599 25483
rect 15761 25449 15795 25483
rect 19717 25449 19751 25483
rect 20085 25449 20119 25483
rect 21373 25449 21407 25483
rect 5181 25381 5215 25415
rect 10517 25381 10551 25415
rect 1409 25313 1443 25347
rect 2513 25313 2547 25347
rect 4077 25313 4111 25347
rect 7941 25313 7975 25347
rect 9781 25313 9815 25347
rect 11345 25313 11379 25347
rect 13001 25313 13035 25347
rect 14197 25313 14231 25347
rect 15577 25313 15611 25347
rect 17049 25313 17083 25347
rect 17141 25313 17175 25347
rect 17601 25313 17635 25347
rect 17785 25313 17819 25347
rect 18705 25313 18739 25347
rect 19901 25313 19935 25347
rect 21189 25313 21223 25347
rect 22293 25313 22327 25347
rect 24041 25313 24075 25347
rect 3801 25245 3835 25279
rect 8033 25245 8067 25279
rect 8125 25245 8159 25279
rect 11437 25245 11471 25279
rect 11529 25245 11563 25279
rect 13093 25245 13127 25279
rect 13277 25245 13311 25279
rect 14105 25245 14139 25279
rect 14565 25245 14599 25279
rect 16497 25245 16531 25279
rect 17325 25245 17359 25279
rect 10793 25177 10827 25211
rect 10977 25177 11011 25211
rect 18797 25245 18831 25279
rect 18981 25245 19015 25279
rect 21557 25245 21591 25279
rect 20453 25177 20487 25211
rect 22477 25177 22511 25211
rect 1593 25109 1627 25143
rect 2053 25109 2087 25143
rect 2329 25109 2363 25143
rect 2697 25109 2731 25143
rect 3157 25109 3191 25143
rect 3433 25109 3467 25143
rect 4261 25109 4295 25143
rect 4721 25109 4755 25143
rect 4997 25109 5031 25143
rect 7389 25109 7423 25143
rect 7573 25109 7607 25143
rect 8677 25109 8711 25143
rect 9597 25109 9631 25143
rect 11989 25109 12023 25143
rect 12449 25109 12483 25143
rect 12633 25109 12667 25143
rect 13645 25109 13679 25143
rect 14841 25109 14875 25143
rect 15209 25109 15243 25143
rect 16681 25109 16715 25143
rect 17601 25109 17635 25143
rect 18153 25109 18187 25143
rect 18337 25109 18371 25143
rect 21557 25109 21591 25143
rect 21741 25109 21775 25143
rect 24225 25109 24259 25143
rect 13461 24905 13495 24939
rect 4537 24837 4571 24871
rect 11069 24837 11103 24871
rect 5089 24769 5123 24803
rect 8677 24769 8711 24803
rect 10241 24769 10275 24803
rect 13093 24769 13127 24803
rect 14197 24769 14231 24803
rect 14841 24769 14875 24803
rect 14933 24769 14967 24803
rect 17049 24769 17083 24803
rect 18613 24769 18647 24803
rect 19533 24769 19567 24803
rect 20085 24769 20119 24803
rect 20269 24769 20303 24803
rect 20729 24769 20763 24803
rect 24961 24769 24995 24803
rect 1409 24701 1443 24735
rect 2329 24701 2363 24735
rect 2513 24701 2547 24735
rect 3065 24701 3099 24735
rect 4905 24701 4939 24735
rect 10149 24701 10183 24735
rect 11253 24701 11287 24735
rect 12817 24701 12851 24735
rect 18429 24701 18463 24735
rect 19993 24701 20027 24735
rect 21649 24701 21683 24735
rect 23857 24701 23891 24735
rect 7113 24633 7147 24667
rect 9137 24633 9171 24667
rect 10057 24633 10091 24667
rect 11897 24633 11931 24667
rect 12909 24633 12943 24667
rect 14749 24633 14783 24667
rect 16313 24633 16347 24667
rect 16865 24633 16899 24667
rect 17877 24633 17911 24667
rect 18521 24633 18555 24667
rect 19073 24633 19107 24667
rect 1593 24565 1627 24599
rect 2053 24565 2087 24599
rect 2697 24565 2731 24599
rect 3709 24565 3743 24599
rect 4077 24565 4111 24599
rect 4997 24565 5031 24599
rect 6561 24565 6595 24599
rect 7665 24565 7699 24599
rect 7941 24565 7975 24599
rect 8125 24565 8159 24599
rect 8493 24565 8527 24599
rect 8585 24565 8619 24599
rect 9505 24565 9539 24599
rect 9689 24565 9723 24599
rect 11437 24565 11471 24599
rect 12265 24565 12299 24599
rect 12449 24565 12483 24599
rect 13829 24565 13863 24599
rect 14381 24565 14415 24599
rect 15669 24565 15703 24599
rect 16405 24565 16439 24599
rect 16773 24565 16807 24599
rect 17509 24565 17543 24599
rect 18061 24565 18095 24599
rect 19625 24565 19659 24599
rect 21281 24565 21315 24599
rect 21833 24565 21867 24599
rect 22385 24565 22419 24599
rect 23489 24565 23523 24599
rect 24041 24565 24075 24599
rect 24409 24565 24443 24599
rect 4813 24361 4847 24395
rect 5181 24361 5215 24395
rect 15301 24361 15335 24395
rect 15669 24361 15703 24395
rect 16497 24361 16531 24395
rect 19165 24361 19199 24395
rect 20637 24361 20671 24395
rect 22661 24361 22695 24395
rect 24685 24361 24719 24395
rect 6193 24293 6227 24327
rect 15025 24293 15059 24327
rect 2053 24225 2087 24259
rect 5273 24225 5307 24259
rect 6920 24225 6954 24259
rect 10681 24225 10715 24259
rect 13277 24225 13311 24259
rect 17509 24225 17543 24259
rect 19073 24225 19107 24259
rect 21281 24225 21315 24259
rect 22477 24225 22511 24259
rect 24501 24225 24535 24259
rect 2145 24157 2179 24191
rect 2329 24157 2363 24191
rect 4721 24157 4755 24191
rect 5457 24157 5491 24191
rect 6653 24157 6687 24191
rect 10425 24157 10459 24191
rect 13369 24157 13403 24191
rect 13461 24157 13495 24191
rect 15761 24157 15795 24191
rect 15853 24157 15887 24191
rect 16865 24157 16899 24191
rect 17601 24157 17635 24191
rect 17785 24157 17819 24191
rect 18245 24157 18279 24191
rect 18613 24157 18647 24191
rect 19257 24157 19291 24191
rect 21373 24157 21407 24191
rect 21465 24157 21499 24191
rect 3341 24089 3375 24123
rect 8953 24089 8987 24123
rect 1685 24021 1719 24055
rect 2789 24021 2823 24055
rect 3709 24021 3743 24055
rect 4353 24021 4387 24055
rect 5917 24021 5951 24055
rect 8033 24021 8067 24055
rect 8677 24021 8711 24055
rect 9965 24021 9999 24055
rect 10333 24021 10367 24055
rect 11805 24021 11839 24055
rect 12633 24021 12667 24055
rect 12909 24021 12943 24055
rect 13921 24021 13955 24055
rect 14473 24021 14507 24055
rect 17141 24021 17175 24055
rect 18705 24021 18739 24055
rect 19809 24021 19843 24055
rect 20269 24021 20303 24055
rect 20913 24021 20947 24055
rect 21925 24021 21959 24055
rect 3617 23817 3651 23851
rect 6193 23817 6227 23851
rect 7481 23817 7515 23851
rect 12173 23817 12207 23851
rect 14749 23817 14783 23851
rect 16589 23817 16623 23851
rect 17233 23817 17267 23851
rect 20361 23817 20395 23851
rect 22293 23817 22327 23851
rect 24777 23817 24811 23851
rect 5181 23749 5215 23783
rect 15025 23749 15059 23783
rect 2145 23681 2179 23715
rect 2237 23681 2271 23715
rect 4077 23681 4111 23715
rect 4261 23681 4295 23715
rect 5641 23681 5675 23715
rect 5825 23681 5859 23715
rect 11253 23681 11287 23715
rect 11437 23681 11471 23715
rect 21189 23681 21223 23715
rect 25145 23681 25179 23715
rect 3985 23613 4019 23647
rect 4629 23613 4663 23647
rect 5549 23613 5583 23647
rect 6837 23613 6871 23647
rect 8033 23613 8067 23647
rect 8125 23613 8159 23647
rect 8392 23613 8426 23647
rect 12449 23613 12483 23647
rect 15209 23613 15243 23647
rect 17877 23613 17911 23647
rect 18061 23613 18095 23647
rect 20913 23613 20947 23647
rect 21925 23613 21959 23647
rect 22109 23613 22143 23647
rect 24593 23613 24627 23647
rect 2053 23545 2087 23579
rect 2789 23545 2823 23579
rect 3065 23545 3099 23579
rect 3525 23545 3559 23579
rect 5089 23545 5123 23579
rect 6653 23545 6687 23579
rect 10517 23545 10551 23579
rect 11897 23545 11931 23579
rect 12694 23545 12728 23579
rect 15454 23545 15488 23579
rect 18306 23545 18340 23579
rect 20085 23545 20119 23579
rect 21649 23545 21683 23579
rect 1685 23477 1719 23511
rect 7021 23477 7055 23511
rect 9505 23477 9539 23511
rect 10149 23477 10183 23511
rect 10793 23477 10827 23511
rect 11161 23477 11195 23511
rect 13829 23477 13863 23511
rect 19441 23477 19475 23511
rect 20545 23477 20579 23511
rect 21005 23477 21039 23511
rect 22661 23477 22695 23511
rect 24409 23477 24443 23511
rect 1593 23273 1627 23307
rect 2421 23273 2455 23307
rect 4813 23273 4847 23307
rect 7205 23273 7239 23307
rect 7849 23273 7883 23307
rect 9137 23273 9171 23307
rect 10057 23273 10091 23307
rect 10885 23273 10919 23307
rect 12357 23273 12391 23307
rect 13185 23273 13219 23307
rect 13277 23273 13311 23307
rect 13921 23273 13955 23307
rect 15025 23273 15059 23307
rect 15485 23273 15519 23307
rect 19441 23273 19475 23307
rect 21925 23273 21959 23307
rect 22937 23273 22971 23307
rect 24777 23273 24811 23307
rect 4445 23205 4479 23239
rect 5150 23205 5184 23239
rect 16764 23205 16798 23239
rect 22293 23205 22327 23239
rect 1409 23137 1443 23171
rect 2789 23137 2823 23171
rect 2881 23137 2915 23171
rect 4905 23137 4939 23171
rect 8401 23137 8435 23171
rect 10149 23137 10183 23171
rect 11621 23137 11655 23171
rect 11713 23137 11747 23171
rect 14565 23137 14599 23171
rect 15301 23137 15335 23171
rect 19349 23137 19383 23171
rect 21281 23137 21315 23171
rect 22845 23137 22879 23171
rect 24593 23137 24627 23171
rect 2329 23069 2363 23103
rect 3065 23069 3099 23103
rect 8493 23069 8527 23103
rect 8585 23069 8619 23103
rect 10333 23069 10367 23103
rect 11805 23069 11839 23103
rect 13369 23069 13403 23103
rect 14197 23069 14231 23103
rect 15945 23069 15979 23103
rect 16497 23069 16531 23103
rect 19533 23069 19567 23103
rect 21373 23069 21407 23103
rect 21557 23069 21591 23103
rect 23121 23069 23155 23103
rect 3525 23001 3559 23035
rect 8033 23001 8067 23035
rect 9689 23001 9723 23035
rect 11253 23001 11287 23035
rect 12725 23001 12759 23035
rect 17877 23001 17911 23035
rect 1869 22933 1903 22967
rect 3893 22933 3927 22967
rect 6285 22933 6319 22967
rect 6929 22933 6963 22967
rect 9505 22933 9539 22967
rect 12817 22933 12851 22967
rect 16405 22933 16439 22967
rect 18705 22933 18739 22967
rect 18981 22933 19015 22967
rect 20269 22933 20303 22967
rect 20545 22933 20579 22967
rect 20913 22933 20947 22967
rect 22477 22933 22511 22967
rect 23489 22933 23523 22967
rect 2053 22729 2087 22763
rect 6837 22729 6871 22763
rect 11069 22729 11103 22763
rect 11437 22729 11471 22763
rect 12449 22729 12483 22763
rect 15669 22729 15703 22763
rect 16221 22729 16255 22763
rect 19533 22729 19567 22763
rect 21005 22729 21039 22763
rect 22845 22729 22879 22763
rect 23857 22729 23891 22763
rect 1593 22661 1627 22695
rect 10793 22661 10827 22695
rect 12265 22661 12299 22695
rect 17049 22661 17083 22695
rect 17877 22661 17911 22695
rect 19625 22661 19659 22695
rect 20729 22661 20763 22695
rect 22569 22661 22603 22695
rect 3157 22593 3191 22627
rect 3341 22593 3375 22627
rect 6193 22593 6227 22627
rect 7481 22593 7515 22627
rect 8585 22593 8619 22627
rect 8677 22593 8711 22627
rect 12909 22593 12943 22627
rect 13001 22593 13035 22627
rect 18521 22593 18555 22627
rect 18705 22593 18739 22627
rect 20269 22593 20303 22627
rect 21741 22593 21775 22627
rect 1409 22525 1443 22559
rect 2605 22525 2639 22559
rect 3065 22525 3099 22559
rect 4169 22525 4203 22559
rect 4261 22525 4295 22559
rect 4528 22525 4562 22559
rect 7205 22525 7239 22559
rect 11253 22525 11287 22559
rect 12817 22525 12851 22559
rect 14289 22525 14323 22559
rect 16865 22525 16899 22559
rect 17417 22525 17451 22559
rect 18429 22525 18463 22559
rect 20085 22525 20119 22559
rect 21557 22525 21591 22559
rect 21649 22525 21683 22559
rect 23673 22525 23707 22559
rect 24225 22525 24259 22559
rect 3709 22457 3743 22491
rect 6653 22457 6687 22491
rect 7297 22457 7331 22491
rect 8217 22457 8251 22491
rect 8944 22457 8978 22491
rect 14556 22457 14590 22491
rect 16681 22457 16715 22491
rect 19165 22457 19199 22491
rect 19993 22457 20027 22491
rect 24685 22457 24719 22491
rect 2697 22389 2731 22423
rect 5641 22389 5675 22423
rect 10057 22389 10091 22423
rect 11897 22389 11931 22423
rect 13461 22389 13495 22423
rect 14197 22389 14231 22423
rect 18061 22389 18095 22423
rect 21189 22389 21223 22423
rect 23213 22389 23247 22423
rect 24777 22389 24811 22423
rect 4813 22185 4847 22219
rect 5457 22185 5491 22219
rect 6837 22185 6871 22219
rect 8033 22185 8067 22219
rect 9873 22185 9907 22219
rect 10333 22185 10367 22219
rect 13553 22185 13587 22219
rect 18521 22185 18555 22219
rect 19349 22185 19383 22219
rect 20269 22185 20303 22219
rect 20913 22185 20947 22219
rect 22477 22185 22511 22219
rect 22661 22185 22695 22219
rect 23029 22185 23063 22219
rect 1777 22117 1811 22151
rect 2237 22117 2271 22151
rect 8401 22117 8435 22151
rect 13921 22117 13955 22151
rect 18061 22117 18095 22151
rect 4353 22049 4387 22083
rect 6377 22049 6411 22083
rect 9413 22049 9447 22083
rect 9689 22049 9723 22083
rect 11336 22049 11370 22083
rect 14933 22049 14967 22083
rect 15301 22049 15335 22083
rect 15568 22049 15602 22083
rect 17233 22049 17267 22083
rect 17693 22049 17727 22083
rect 2329 21981 2363 22015
rect 2421 21981 2455 22015
rect 4905 21981 4939 22015
rect 4997 21981 5031 22015
rect 6929 21981 6963 22015
rect 7113 21981 7147 22015
rect 8493 21981 8527 22015
rect 8585 21981 8619 22015
rect 9137 21981 9171 22015
rect 11069 21981 11103 22015
rect 14013 21981 14047 22015
rect 14105 21981 14139 22015
rect 18613 21981 18647 22015
rect 18705 21981 18739 22015
rect 20453 22117 20487 22151
rect 19717 22049 19751 22083
rect 1869 21913 1903 21947
rect 6469 21913 6503 21947
rect 12449 21913 12483 21947
rect 18153 21913 18187 21947
rect 19349 21913 19383 21947
rect 19625 21913 19659 21947
rect 21465 22117 21499 22151
rect 22109 22117 22143 22151
rect 24593 22117 24627 22151
rect 21557 21981 21591 22015
rect 21741 21981 21775 22015
rect 23121 21981 23155 22015
rect 23305 21981 23339 22015
rect 24685 21981 24719 22015
rect 24777 21981 24811 22015
rect 2973 21845 3007 21879
rect 3525 21845 3559 21879
rect 3801 21845 3835 21879
rect 4445 21845 4479 21879
rect 6009 21845 6043 21879
rect 7665 21845 7699 21879
rect 10609 21845 10643 21879
rect 13369 21845 13403 21879
rect 14657 21845 14691 21879
rect 16681 21845 16715 21879
rect 19257 21845 19291 21879
rect 19901 21845 19935 21879
rect 20453 21845 20487 21879
rect 20729 21845 20763 21879
rect 20913 21845 20947 21879
rect 21097 21845 21131 21879
rect 23765 21845 23799 21879
rect 24041 21845 24075 21879
rect 24225 21845 24259 21879
rect 1685 21641 1719 21675
rect 1869 21641 1903 21675
rect 4997 21641 5031 21675
rect 9045 21641 9079 21675
rect 10149 21641 10183 21675
rect 11529 21641 11563 21675
rect 12817 21641 12851 21675
rect 13185 21641 13219 21675
rect 15301 21641 15335 21675
rect 17509 21641 17543 21675
rect 20545 21641 20579 21675
rect 21097 21641 21131 21675
rect 23029 21641 23063 21675
rect 25053 21641 25087 21675
rect 25421 21641 25455 21675
rect 3249 21573 3283 21607
rect 3433 21573 3467 21607
rect 9781 21573 9815 21607
rect 23397 21573 23431 21607
rect 2329 21505 2363 21539
rect 2513 21505 2547 21539
rect 3985 21505 4019 21539
rect 4537 21505 4571 21539
rect 5549 21505 5583 21539
rect 10701 21505 10735 21539
rect 11897 21505 11931 21539
rect 13277 21505 13311 21539
rect 16313 21505 16347 21539
rect 17049 21505 17083 21539
rect 18613 21505 18647 21539
rect 21741 21505 21775 21539
rect 24133 21505 24167 21539
rect 24317 21505 24351 21539
rect 2237 21437 2271 21471
rect 2881 21437 2915 21471
rect 3893 21437 3927 21471
rect 6101 21437 6135 21471
rect 7665 21437 7699 21471
rect 11253 21437 11287 21471
rect 16773 21437 16807 21471
rect 17877 21437 17911 21471
rect 21465 21437 21499 21471
rect 25237 21437 25271 21471
rect 4813 21369 4847 21403
rect 5365 21369 5399 21403
rect 7021 21369 7055 21403
rect 7910 21369 7944 21403
rect 10609 21369 10643 21403
rect 13544 21369 13578 21403
rect 18858 21369 18892 21403
rect 24041 21369 24075 21403
rect 3801 21301 3835 21335
rect 5457 21301 5491 21335
rect 6561 21301 6595 21335
rect 7573 21301 7607 21335
rect 10517 21301 10551 21335
rect 14657 21301 14691 21335
rect 15669 21301 15703 21335
rect 16405 21301 16439 21335
rect 16865 21301 16899 21335
rect 18429 21301 18463 21335
rect 19993 21301 20027 21335
rect 20913 21301 20947 21335
rect 21557 21301 21591 21335
rect 22109 21301 22143 21335
rect 22753 21301 22787 21335
rect 23673 21301 23707 21335
rect 24685 21301 24719 21335
rect 25789 21301 25823 21335
rect 1777 21097 1811 21131
rect 1961 21097 1995 21131
rect 2421 21097 2455 21131
rect 4077 21097 4111 21131
rect 5457 21097 5491 21131
rect 5641 21097 5675 21131
rect 7113 21097 7147 21131
rect 8309 21097 8343 21131
rect 9045 21097 9079 21131
rect 11805 21097 11839 21131
rect 12265 21097 12299 21131
rect 13645 21097 13679 21131
rect 14289 21097 14323 21131
rect 15761 21097 15795 21131
rect 16865 21097 16899 21131
rect 17601 21097 17635 21131
rect 18061 21097 18095 21131
rect 19257 21097 19291 21131
rect 20361 21097 20395 21131
rect 20729 21097 20763 21131
rect 21189 21097 21223 21131
rect 24593 21097 24627 21131
rect 4537 21029 4571 21063
rect 7665 21029 7699 21063
rect 15117 21029 15151 21063
rect 16497 21029 16531 21063
rect 18153 21029 18187 21063
rect 19073 21029 19107 21063
rect 21557 21029 21591 21063
rect 24685 21029 24719 21063
rect 2329 20961 2363 20995
rect 2973 20961 3007 20995
rect 4445 20961 4479 20995
rect 6009 20961 6043 20995
rect 7573 20961 7607 20995
rect 9781 20961 9815 20995
rect 10037 20961 10071 20995
rect 12173 20961 12207 20995
rect 12633 20961 12667 20995
rect 12725 20961 12759 20995
rect 14105 20961 14139 20995
rect 15669 20961 15703 20995
rect 18797 20961 18831 20995
rect 19625 20961 19659 20995
rect 21997 20961 22031 20995
rect 25237 20961 25271 20995
rect 2605 20893 2639 20927
rect 3893 20893 3927 20927
rect 4721 20893 4755 20927
rect 6101 20893 6135 20927
rect 6285 20893 6319 20927
rect 7757 20893 7791 20927
rect 12909 20893 12943 20927
rect 15853 20893 15887 20927
rect 18337 20893 18371 20927
rect 19717 20893 19751 20927
rect 19809 20893 19843 20927
rect 21741 20893 21775 20927
rect 24777 20893 24811 20927
rect 8677 20825 8711 20859
rect 11161 20825 11195 20859
rect 14749 20825 14783 20859
rect 15301 20825 15335 20859
rect 17233 20825 17267 20859
rect 17693 20825 17727 20859
rect 3525 20757 3559 20791
rect 5089 20757 5123 20791
rect 6745 20757 6779 20791
rect 7205 20757 7239 20791
rect 9413 20757 9447 20791
rect 14013 20757 14047 20791
rect 23121 20757 23155 20791
rect 23673 20757 23707 20791
rect 24041 20757 24075 20791
rect 24225 20757 24259 20791
rect 1777 20553 1811 20587
rect 1961 20553 1995 20587
rect 3065 20553 3099 20587
rect 6193 20553 6227 20587
rect 6561 20553 6595 20587
rect 10241 20553 10275 20587
rect 12449 20553 12483 20587
rect 13461 20553 13495 20587
rect 14013 20553 14047 20587
rect 15761 20553 15795 20587
rect 17785 20553 17819 20587
rect 18521 20553 18555 20587
rect 21097 20553 21131 20587
rect 3341 20485 3375 20519
rect 12081 20485 12115 20519
rect 12173 20485 12207 20519
rect 13921 20485 13955 20519
rect 16405 20485 16439 20519
rect 2421 20417 2455 20451
rect 2605 20417 2639 20451
rect 10793 20417 10827 20451
rect 11253 20417 11287 20451
rect 11805 20417 11839 20451
rect 3709 20349 3743 20383
rect 3893 20349 3927 20383
rect 5825 20349 5859 20383
rect 7757 20349 7791 20383
rect 8013 20349 8047 20383
rect 9689 20349 9723 20383
rect 10701 20349 10735 20383
rect 13001 20417 13035 20451
rect 14473 20417 14507 20451
rect 14657 20417 14691 20451
rect 16957 20417 16991 20451
rect 18981 20417 19015 20451
rect 19073 20417 19107 20451
rect 22017 20417 22051 20451
rect 22201 20417 22235 20451
rect 22937 20417 22971 20451
rect 19340 20349 19374 20383
rect 22661 20349 22695 20383
rect 23489 20349 23523 20383
rect 23673 20349 23707 20383
rect 25973 20349 26007 20383
rect 4138 20281 4172 20315
rect 7665 20281 7699 20315
rect 10609 20281 10643 20315
rect 12081 20281 12115 20315
rect 12817 20281 12851 20315
rect 15301 20281 15335 20315
rect 16773 20281 16807 20315
rect 18061 20281 18095 20315
rect 21465 20281 21499 20315
rect 21925 20281 21959 20315
rect 23918 20281 23952 20315
rect 25605 20281 25639 20315
rect 2329 20213 2363 20247
rect 5273 20213 5307 20247
rect 7205 20213 7239 20247
rect 9137 20213 9171 20247
rect 10057 20213 10091 20247
rect 12909 20213 12943 20247
rect 14381 20213 14415 20247
rect 16221 20213 16255 20247
rect 16865 20213 16899 20247
rect 20453 20213 20487 20247
rect 21557 20213 21591 20247
rect 25053 20213 25087 20247
rect 2053 20009 2087 20043
rect 6837 20009 6871 20043
rect 7849 20009 7883 20043
rect 8309 20009 8343 20043
rect 9689 20009 9723 20043
rect 10333 20009 10367 20043
rect 11161 20009 11195 20043
rect 12541 20009 12575 20043
rect 15117 20009 15151 20043
rect 15761 20009 15795 20043
rect 16497 20009 16531 20043
rect 17417 20009 17451 20043
rect 18153 20009 18187 20043
rect 19625 20009 19659 20043
rect 23213 20009 23247 20043
rect 23857 20009 23891 20043
rect 24501 20009 24535 20043
rect 24869 20009 24903 20043
rect 25145 20009 25179 20043
rect 2881 19941 2915 19975
rect 3525 19941 3559 19975
rect 3893 19941 3927 19975
rect 12081 19941 12115 19975
rect 17509 19941 17543 19975
rect 19073 19941 19107 19975
rect 21180 19941 21214 19975
rect 2789 19873 2823 19907
rect 4077 19873 4111 19907
rect 4721 19873 4755 19907
rect 5457 19873 5491 19907
rect 5724 19873 5758 19907
rect 7481 19873 7515 19907
rect 8401 19873 8435 19907
rect 11069 19873 11103 19907
rect 12981 19873 13015 19907
rect 15669 19873 15703 19907
rect 18981 19873 19015 19907
rect 19441 19873 19475 19907
rect 23765 19873 23799 19907
rect 24685 19873 24719 19907
rect 24949 19873 24983 19907
rect 1409 19805 1443 19839
rect 3065 19805 3099 19839
rect 8585 19805 8619 19839
rect 11253 19805 11287 19839
rect 11713 19805 11747 19839
rect 12725 19805 12759 19839
rect 15853 19805 15887 19839
rect 17601 19805 17635 19839
rect 18429 19805 18463 19839
rect 19257 19805 19291 19839
rect 20913 19805 20947 19839
rect 22845 19805 22879 19839
rect 24041 19805 24075 19839
rect 5089 19737 5123 19771
rect 7941 19737 7975 19771
rect 9137 19737 9171 19771
rect 10701 19737 10735 19771
rect 14657 19737 14691 19771
rect 17049 19737 17083 19771
rect 19441 19737 19475 19771
rect 20729 19737 20763 19771
rect 2421 19669 2455 19703
rect 4261 19669 4295 19703
rect 9505 19669 9539 19703
rect 14105 19669 14139 19703
rect 15301 19669 15335 19703
rect 16957 19669 16991 19703
rect 18613 19669 18647 19703
rect 20361 19669 20395 19703
rect 22293 19669 22327 19703
rect 23397 19669 23431 19703
rect 24685 19669 24719 19703
rect 7849 19465 7883 19499
rect 9413 19465 9447 19499
rect 12725 19465 12759 19499
rect 16865 19465 16899 19499
rect 17417 19465 17451 19499
rect 24961 19465 24995 19499
rect 12173 19397 12207 19431
rect 15117 19397 15151 19431
rect 23489 19397 23523 19431
rect 3801 19329 3835 19363
rect 8033 19329 8067 19363
rect 11345 19329 11379 19363
rect 11897 19329 11931 19363
rect 13737 19329 13771 19363
rect 15669 19329 15703 19363
rect 19257 19329 19291 19363
rect 20913 19329 20947 19363
rect 22477 19329 22511 19363
rect 22661 19329 22695 19363
rect 24225 19329 24259 19363
rect 1777 19261 1811 19295
rect 4077 19261 4111 19295
rect 4261 19261 4295 19295
rect 4528 19261 4562 19295
rect 6837 19261 6871 19295
rect 14289 19261 14323 19295
rect 15577 19261 15611 19295
rect 16957 19261 16991 19295
rect 19073 19261 19107 19295
rect 20085 19261 20119 19295
rect 20729 19261 20763 19295
rect 23121 19261 23155 19295
rect 24041 19261 24075 19295
rect 25237 19261 25271 19295
rect 25789 19261 25823 19295
rect 2044 19193 2078 19227
rect 8278 19193 8312 19227
rect 10701 19193 10735 19227
rect 11161 19193 11195 19227
rect 15485 19193 15519 19227
rect 19165 19193 19199 19227
rect 19717 19193 19751 19227
rect 21649 19193 21683 19227
rect 22385 19193 22419 19227
rect 1685 19125 1719 19159
rect 3157 19125 3191 19159
rect 5641 19125 5675 19159
rect 6285 19125 6319 19159
rect 6653 19125 6687 19159
rect 7021 19125 7055 19159
rect 7481 19125 7515 19159
rect 10241 19125 10275 19159
rect 10793 19125 10827 19159
rect 11253 19125 11287 19159
rect 13185 19125 13219 19159
rect 13553 19125 13587 19159
rect 13645 19125 13679 19159
rect 14565 19125 14599 19159
rect 14933 19125 14967 19159
rect 16221 19125 16255 19159
rect 17141 19125 17175 19159
rect 17785 19125 17819 19159
rect 18521 19125 18555 19159
rect 18705 19125 18739 19159
rect 20269 19125 20303 19159
rect 20637 19125 20671 19159
rect 21373 19125 21407 19159
rect 22017 19125 22051 19159
rect 23673 19125 23707 19159
rect 24133 19125 24167 19159
rect 25421 19125 25455 19159
rect 1593 18921 1627 18955
rect 2789 18921 2823 18955
rect 4629 18921 4663 18955
rect 6745 18921 6779 18955
rect 8033 18921 8067 18955
rect 12173 18921 12207 18955
rect 12817 18921 12851 18955
rect 13277 18921 13311 18955
rect 14841 18921 14875 18955
rect 15485 18921 15519 18955
rect 16129 18921 16163 18955
rect 17785 18921 17819 18955
rect 19993 18921 20027 18955
rect 20913 18921 20947 18955
rect 22109 18921 22143 18955
rect 23857 18921 23891 18955
rect 24777 18921 24811 18955
rect 25145 18921 25179 18955
rect 2881 18853 2915 18887
rect 5632 18853 5666 18887
rect 9413 18853 9447 18887
rect 13829 18853 13863 18887
rect 15853 18853 15887 18887
rect 20729 18853 20763 18887
rect 21373 18853 21407 18887
rect 22744 18853 22778 18887
rect 1409 18785 1443 18819
rect 4077 18785 4111 18819
rect 5365 18785 5399 18819
rect 8401 18785 8435 18819
rect 8493 18785 8527 18819
rect 9689 18785 9723 18819
rect 10793 18785 10827 18819
rect 11060 18785 11094 18819
rect 13737 18785 13771 18819
rect 15301 18785 15335 18819
rect 16672 18785 16706 18819
rect 19257 18785 19291 18819
rect 19349 18785 19383 18819
rect 21281 18785 21315 18819
rect 22477 18785 22511 18819
rect 24961 18785 24995 18819
rect 3065 18717 3099 18751
rect 8585 18717 8619 18751
rect 10241 18717 10275 18751
rect 10609 18717 10643 18751
rect 13921 18717 13955 18751
rect 16405 18717 16439 18751
rect 18429 18717 18463 18751
rect 19441 18717 19475 18751
rect 21465 18717 21499 18751
rect 9873 18649 9907 18683
rect 1961 18581 1995 18615
rect 2421 18581 2455 18615
rect 3433 18581 3467 18615
rect 3801 18581 3835 18615
rect 4261 18581 4295 18615
rect 5273 18581 5307 18615
rect 7573 18581 7607 18615
rect 7941 18581 7975 18615
rect 9045 18581 9079 18615
rect 13369 18581 13403 18615
rect 14381 18581 14415 18615
rect 18705 18581 18739 18615
rect 18889 18581 18923 18615
rect 20361 18581 20395 18615
rect 24409 18581 24443 18615
rect 1869 18377 1903 18411
rect 4169 18377 4203 18411
rect 5089 18377 5123 18411
rect 6285 18377 6319 18411
rect 7113 18377 7147 18411
rect 9229 18377 9263 18411
rect 10241 18377 10275 18411
rect 13461 18377 13495 18411
rect 13829 18377 13863 18411
rect 14933 18377 14967 18411
rect 17049 18377 17083 18411
rect 17417 18377 17451 18411
rect 18705 18377 18739 18411
rect 20545 18377 20579 18411
rect 21649 18377 21683 18411
rect 22753 18377 22787 18411
rect 23029 18377 23063 18411
rect 23673 18377 23707 18411
rect 25421 18377 25455 18411
rect 4445 18309 4479 18343
rect 9137 18309 9171 18343
rect 10609 18309 10643 18343
rect 18337 18309 18371 18343
rect 25053 18309 25087 18343
rect 5825 18241 5859 18275
rect 6653 18241 6687 18275
rect 8125 18241 8159 18275
rect 8217 18241 8251 18275
rect 9689 18241 9723 18275
rect 9781 18241 9815 18275
rect 11345 18241 11379 18275
rect 12265 18241 12299 18275
rect 13001 18241 13035 18275
rect 14013 18241 14047 18275
rect 15117 18241 15151 18275
rect 18981 18241 19015 18275
rect 19165 18241 19199 18275
rect 22201 18241 22235 18275
rect 24225 18241 24259 18275
rect 24685 18241 24719 18275
rect 1961 18173 1995 18207
rect 8033 18173 8067 18207
rect 11161 18173 11195 18207
rect 12817 18173 12851 18207
rect 15384 18173 15418 18207
rect 17877 18173 17911 18207
rect 18153 18173 18187 18207
rect 19432 18173 19466 18207
rect 24133 18173 24167 18207
rect 25237 18173 25271 18207
rect 25789 18173 25823 18207
rect 2228 18105 2262 18139
rect 5549 18105 5583 18139
rect 9597 18105 9631 18139
rect 14657 18105 14691 18139
rect 21097 18105 21131 18139
rect 21557 18105 21591 18139
rect 22109 18105 22143 18139
rect 23489 18105 23523 18139
rect 24041 18105 24075 18139
rect 3341 18037 3375 18071
rect 5181 18037 5215 18071
rect 5641 18037 5675 18071
rect 7481 18037 7515 18071
rect 7665 18037 7699 18071
rect 8769 18037 8803 18071
rect 10793 18037 10827 18071
rect 11253 18037 11287 18071
rect 11805 18037 11839 18071
rect 12449 18037 12483 18071
rect 12909 18037 12943 18071
rect 16497 18037 16531 18071
rect 22017 18037 22051 18071
rect 1593 17833 1627 17867
rect 2329 17833 2363 17867
rect 4905 17833 4939 17867
rect 7757 17833 7791 17867
rect 10057 17833 10091 17867
rect 10885 17833 10919 17867
rect 11161 17833 11195 17867
rect 11529 17833 11563 17867
rect 12081 17833 12115 17867
rect 12633 17833 12667 17867
rect 13461 17833 13495 17867
rect 14565 17833 14599 17867
rect 15117 17833 15151 17867
rect 18245 17833 18279 17867
rect 18797 17833 18831 17867
rect 19257 17833 19291 17867
rect 20269 17833 20303 17867
rect 20729 17833 20763 17867
rect 22569 17833 22603 17867
rect 24133 17833 24167 17867
rect 25421 17833 25455 17867
rect 2789 17765 2823 17799
rect 3525 17765 3559 17799
rect 3893 17765 3927 17799
rect 6837 17765 6871 17799
rect 14197 17765 14231 17799
rect 15568 17765 15602 17799
rect 22017 17765 22051 17799
rect 22998 17765 23032 17799
rect 1409 17697 1443 17731
rect 4813 17697 4847 17731
rect 5273 17697 5307 17731
rect 6285 17697 6319 17731
rect 8401 17697 8435 17731
rect 12541 17697 12575 17731
rect 13737 17697 13771 17731
rect 18153 17697 18187 17731
rect 19809 17697 19843 17731
rect 21281 17697 21315 17731
rect 21373 17697 21407 17731
rect 22753 17697 22787 17731
rect 25237 17697 25271 17731
rect 2881 17629 2915 17663
rect 2973 17629 3007 17663
rect 5365 17629 5399 17663
rect 5457 17629 5491 17663
rect 6929 17629 6963 17663
rect 7021 17629 7055 17663
rect 8493 17629 8527 17663
rect 8585 17629 8619 17663
rect 10149 17629 10183 17663
rect 10333 17629 10367 17663
rect 12817 17629 12851 17663
rect 15301 17629 15335 17663
rect 18429 17629 18463 17663
rect 21465 17629 21499 17663
rect 1961 17561 1995 17595
rect 4445 17561 4479 17595
rect 5917 17561 5951 17595
rect 9137 17561 9171 17595
rect 9689 17561 9723 17595
rect 13921 17561 13955 17595
rect 17325 17561 17359 17595
rect 17785 17561 17819 17595
rect 20913 17561 20947 17595
rect 2421 17493 2455 17527
rect 6469 17493 6503 17527
rect 8033 17493 8067 17527
rect 9413 17493 9447 17527
rect 12173 17493 12207 17527
rect 16681 17493 16715 17527
rect 17601 17493 17635 17527
rect 19717 17493 19751 17527
rect 19993 17493 20027 17527
rect 24685 17493 24719 17527
rect 25053 17493 25087 17527
rect 1961 17289 1995 17323
rect 4261 17289 4295 17323
rect 5181 17289 5215 17323
rect 6561 17289 6595 17323
rect 8125 17289 8159 17323
rect 9413 17289 9447 17323
rect 11897 17289 11931 17323
rect 15301 17289 15335 17323
rect 15853 17289 15887 17323
rect 17509 17289 17543 17323
rect 17877 17289 17911 17323
rect 19165 17289 19199 17323
rect 21649 17289 21683 17323
rect 22385 17289 22419 17323
rect 23029 17289 23063 17323
rect 23489 17289 23523 17323
rect 23673 17289 23707 17323
rect 25421 17289 25455 17323
rect 25881 17289 25915 17323
rect 4629 17221 4663 17255
rect 9689 17221 9723 17255
rect 11253 17221 11287 17255
rect 5733 17153 5767 17187
rect 8769 17153 8803 17187
rect 8953 17153 8987 17187
rect 12173 17153 12207 17187
rect 12449 17153 12483 17187
rect 15393 17153 15427 17187
rect 16957 17153 16991 17187
rect 18613 17153 18647 17187
rect 24225 17153 24259 17187
rect 2053 17085 2087 17119
rect 6837 17085 6871 17119
rect 7389 17085 7423 17119
rect 8677 17085 8711 17119
rect 9873 17085 9907 17119
rect 14381 17085 14415 17119
rect 16773 17085 16807 17119
rect 18521 17085 18555 17119
rect 19533 17085 19567 17119
rect 19625 17085 19659 17119
rect 22477 17085 22511 17119
rect 24041 17085 24075 17119
rect 25237 17085 25271 17119
rect 2320 17017 2354 17051
rect 5549 17017 5583 17051
rect 10140 17017 10174 17051
rect 12694 17017 12728 17051
rect 16313 17017 16347 17051
rect 18429 17017 18463 17051
rect 19870 17017 19904 17051
rect 24133 17017 24167 17051
rect 24777 17017 24811 17051
rect 3433 16949 3467 16983
rect 4997 16949 5031 16983
rect 5641 16949 5675 16983
rect 7021 16949 7055 16983
rect 8309 16949 8343 16983
rect 13829 16949 13863 16983
rect 14933 16949 14967 16983
rect 16405 16949 16439 16983
rect 16865 16949 16899 16983
rect 18061 16949 18095 16983
rect 21005 16949 21039 16983
rect 22661 16949 22695 16983
rect 25053 16949 25087 16983
rect 2789 16745 2823 16779
rect 3249 16745 3283 16779
rect 3801 16745 3835 16779
rect 6377 16745 6411 16779
rect 8861 16745 8895 16779
rect 9505 16745 9539 16779
rect 9965 16745 9999 16779
rect 14565 16745 14599 16779
rect 15577 16745 15611 16779
rect 16129 16745 16163 16779
rect 18337 16745 18371 16779
rect 19257 16745 19291 16779
rect 19717 16745 19751 16779
rect 20269 16745 20303 16779
rect 20637 16745 20671 16779
rect 20913 16745 20947 16779
rect 21281 16745 21315 16779
rect 21925 16745 21959 16779
rect 22477 16745 22511 16779
rect 24133 16745 24167 16779
rect 25053 16745 25087 16779
rect 25421 16745 25455 16779
rect 2145 16677 2179 16711
rect 1409 16609 1443 16643
rect 2881 16609 2915 16643
rect 2973 16541 3007 16575
rect 1593 16473 1627 16507
rect 4322 16677 4356 16711
rect 6101 16677 6135 16711
rect 6806 16677 6840 16711
rect 8585 16677 8619 16711
rect 10600 16677 10634 16711
rect 13921 16677 13955 16711
rect 18613 16677 18647 16711
rect 21373 16677 21407 16711
rect 23020 16677 23054 16711
rect 4077 16609 4111 16643
rect 10333 16609 10367 16643
rect 12541 16609 12575 16643
rect 13185 16609 13219 16643
rect 14197 16609 14231 16643
rect 15117 16609 15151 16643
rect 16037 16609 16071 16643
rect 17049 16609 17083 16643
rect 17601 16609 17635 16643
rect 19165 16609 19199 16643
rect 19625 16609 19659 16643
rect 22753 16609 22787 16643
rect 25237 16609 25271 16643
rect 6561 16541 6595 16575
rect 13277 16541 13311 16575
rect 13461 16541 13495 16575
rect 16221 16541 16255 16575
rect 17693 16541 17727 16575
rect 17785 16541 17819 16575
rect 19809 16541 19843 16575
rect 21557 16541 21591 16575
rect 24685 16473 24719 16507
rect 2421 16405 2455 16439
rect 3249 16405 3283 16439
rect 3433 16405 3467 16439
rect 5457 16405 5491 16439
rect 7941 16405 7975 16439
rect 11713 16405 11747 16439
rect 12817 16405 12851 16439
rect 15669 16405 15703 16439
rect 16773 16405 16807 16439
rect 17233 16405 17267 16439
rect 25789 16405 25823 16439
rect 2053 16201 2087 16235
rect 3433 16201 3467 16235
rect 5089 16201 5123 16235
rect 8217 16201 8251 16235
rect 9505 16201 9539 16235
rect 9689 16201 9723 16235
rect 10701 16201 10735 16235
rect 11161 16201 11195 16235
rect 11897 16201 11931 16235
rect 12449 16201 12483 16235
rect 13461 16201 13495 16235
rect 14013 16201 14047 16235
rect 16405 16201 16439 16235
rect 18613 16201 18647 16235
rect 20453 16201 20487 16235
rect 21097 16201 21131 16235
rect 22753 16201 22787 16235
rect 23213 16201 23247 16235
rect 23673 16201 23707 16235
rect 25421 16201 25455 16235
rect 3617 16133 3651 16167
rect 16313 16133 16347 16167
rect 17877 16133 17911 16167
rect 18889 16133 18923 16167
rect 2513 16065 2547 16099
rect 2697 16065 2731 16099
rect 4169 16065 4203 16099
rect 5733 16065 5767 16099
rect 10149 16065 10183 16099
rect 10333 16065 10367 16099
rect 12265 16065 12299 16099
rect 13001 16065 13035 16099
rect 14565 16065 14599 16099
rect 16957 16065 16991 16099
rect 19073 16065 19107 16099
rect 22293 16065 22327 16099
rect 24317 16065 24351 16099
rect 24685 16065 24719 16099
rect 3985 15997 4019 16031
rect 6837 15997 6871 16031
rect 7093 15997 7127 16031
rect 8861 15997 8895 16031
rect 11253 15997 11287 16031
rect 12817 15997 12851 16031
rect 15025 15997 15059 16031
rect 15945 15997 15979 16031
rect 16865 15997 16899 16031
rect 21557 15997 21591 16031
rect 22017 15997 22051 16031
rect 25237 15997 25271 16031
rect 25789 15997 25823 16031
rect 26249 15997 26283 16031
rect 3065 15929 3099 15963
rect 4077 15929 4111 15963
rect 5549 15929 5583 15963
rect 9229 15929 9263 15963
rect 10057 15929 10091 15963
rect 12909 15929 12943 15963
rect 14473 15929 14507 15963
rect 16773 15929 16807 15963
rect 19318 15929 19352 15963
rect 22109 15929 22143 15963
rect 24133 15929 24167 15963
rect 25145 15929 25179 15963
rect 1961 15861 1995 15895
rect 2421 15861 2455 15895
rect 4721 15861 4755 15895
rect 5181 15861 5215 15895
rect 5641 15861 5675 15895
rect 6285 15861 6319 15895
rect 6561 15861 6595 15895
rect 13829 15861 13863 15895
rect 14381 15861 14415 15895
rect 15577 15861 15611 15895
rect 17417 15861 17451 15895
rect 18061 15861 18095 15895
rect 21649 15861 21683 15895
rect 24041 15861 24075 15895
rect 2145 15657 2179 15691
rect 3893 15657 3927 15691
rect 8033 15657 8067 15691
rect 10609 15657 10643 15691
rect 12173 15657 12207 15691
rect 12817 15657 12851 15691
rect 13645 15657 13679 15691
rect 14289 15657 14323 15691
rect 14657 15657 14691 15691
rect 17141 15657 17175 15691
rect 18705 15657 18739 15691
rect 19349 15657 19383 15691
rect 20361 15657 20395 15691
rect 20637 15657 20671 15691
rect 20913 15657 20947 15691
rect 21373 15657 21407 15691
rect 22017 15657 22051 15691
rect 22293 15657 22327 15691
rect 24777 15657 24811 15691
rect 25145 15657 25179 15691
rect 2789 15589 2823 15623
rect 4629 15589 4663 15623
rect 4988 15589 5022 15623
rect 6653 15589 6687 15623
rect 7113 15589 7147 15623
rect 8401 15589 8435 15623
rect 10241 15589 10275 15623
rect 11060 15589 11094 15623
rect 13185 15589 13219 15623
rect 19717 15589 19751 15623
rect 25513 15589 25547 15623
rect 1409 15521 1443 15555
rect 4721 15521 4755 15555
rect 8493 15521 8527 15555
rect 9689 15521 9723 15555
rect 10793 15521 10827 15555
rect 16028 15521 16062 15555
rect 18613 15521 18647 15555
rect 19809 15521 19843 15555
rect 21281 15521 21315 15555
rect 22733 15521 22767 15555
rect 24961 15521 24995 15555
rect 2881 15453 2915 15487
rect 3065 15453 3099 15487
rect 8585 15453 8619 15487
rect 8861 15453 8895 15487
rect 9413 15453 9447 15487
rect 13737 15453 13771 15487
rect 13921 15453 13955 15487
rect 15117 15453 15151 15487
rect 15761 15453 15795 15487
rect 18797 15453 18831 15487
rect 21465 15453 21499 15487
rect 22477 15453 22511 15487
rect 6101 15385 6135 15419
rect 7389 15385 7423 15419
rect 7757 15385 7791 15419
rect 9873 15385 9907 15419
rect 18245 15385 18279 15419
rect 1593 15317 1627 15351
rect 2421 15317 2455 15351
rect 3525 15317 3559 15351
rect 8861 15317 8895 15351
rect 9045 15317 9079 15351
rect 13277 15317 13311 15351
rect 15485 15317 15519 15351
rect 17693 15317 17727 15351
rect 18153 15317 18187 15351
rect 23857 15317 23891 15351
rect 24409 15317 24443 15351
rect 1961 15113 1995 15147
rect 7021 15113 7055 15147
rect 8125 15113 8159 15147
rect 8401 15113 8435 15147
rect 10885 15113 10919 15147
rect 12725 15113 12759 15147
rect 14473 15113 14507 15147
rect 17417 15113 17451 15147
rect 19533 15113 19567 15147
rect 21925 15113 21959 15147
rect 24961 15113 24995 15147
rect 25421 15113 25455 15147
rect 2421 15045 2455 15079
rect 6009 15045 6043 15079
rect 14197 15045 14231 15079
rect 18889 15045 18923 15079
rect 22385 15045 22419 15079
rect 23029 15045 23063 15079
rect 26249 15045 26283 15079
rect 2881 14977 2915 15011
rect 3065 14977 3099 15011
rect 7573 14977 7607 15011
rect 11069 14977 11103 15011
rect 13277 14977 13311 15011
rect 15301 14977 15335 15011
rect 15485 14977 15519 15011
rect 17785 14977 17819 15011
rect 18521 14977 18555 15011
rect 18613 14977 18647 15011
rect 1409 14909 1443 14943
rect 2789 14909 2823 14943
rect 3893 14909 3927 14943
rect 3985 14909 4019 14943
rect 7481 14909 7515 14943
rect 8585 14909 8619 14943
rect 13093 14909 13127 14943
rect 13185 14909 13219 14943
rect 14289 14909 14323 14943
rect 24133 14977 24167 15011
rect 24225 14977 24259 15011
rect 19993 14909 20027 14943
rect 22477 14909 22511 14943
rect 23489 14909 23523 14943
rect 25237 14909 25271 14943
rect 25789 14909 25823 14943
rect 4252 14841 4286 14875
rect 6653 14841 6687 14875
rect 8830 14841 8864 14875
rect 15025 14841 15059 14875
rect 15752 14841 15786 14875
rect 18889 14841 18923 14875
rect 19073 14841 19107 14875
rect 20260 14841 20294 14875
rect 1593 14773 1627 14807
rect 2329 14773 2363 14807
rect 3525 14773 3559 14807
rect 5365 14773 5399 14807
rect 7389 14773 7423 14807
rect 9965 14773 9999 14807
rect 10609 14773 10643 14807
rect 11621 14773 11655 14807
rect 12265 14773 12299 14807
rect 13829 14773 13863 14807
rect 16865 14773 16899 14807
rect 18061 14773 18095 14807
rect 18429 14773 18463 14807
rect 19809 14773 19843 14807
rect 21373 14773 21407 14807
rect 22661 14773 22695 14807
rect 23673 14773 23707 14807
rect 24041 14773 24075 14807
rect 1961 14569 1995 14603
rect 2421 14569 2455 14603
rect 3433 14569 3467 14603
rect 3893 14569 3927 14603
rect 6193 14569 6227 14603
rect 8033 14569 8067 14603
rect 8401 14569 8435 14603
rect 10241 14569 10275 14603
rect 10885 14569 10919 14603
rect 13369 14569 13403 14603
rect 13921 14569 13955 14603
rect 14289 14569 14323 14603
rect 15117 14569 15151 14603
rect 17877 14569 17911 14603
rect 18429 14569 18463 14603
rect 19257 14569 19291 14603
rect 19625 14569 19659 14603
rect 21097 14569 21131 14603
rect 21465 14569 21499 14603
rect 23673 14569 23707 14603
rect 24777 14569 24811 14603
rect 2881 14501 2915 14535
rect 7389 14501 7423 14535
rect 7849 14501 7883 14535
rect 8493 14501 8527 14535
rect 11897 14501 11931 14535
rect 12234 14501 12268 14535
rect 15945 14501 15979 14535
rect 16405 14501 16439 14535
rect 21925 14501 21959 14535
rect 1409 14433 1443 14467
rect 2789 14433 2823 14467
rect 4517 14433 4551 14467
rect 6745 14433 6779 14467
rect 11989 14433 12023 14467
rect 16497 14433 16531 14467
rect 16764 14433 16798 14467
rect 20913 14433 20947 14467
rect 22560 14433 22594 14467
rect 25145 14433 25179 14467
rect 2973 14365 3007 14399
rect 4261 14365 4295 14399
rect 8585 14365 8619 14399
rect 10333 14365 10367 14399
rect 10517 14365 10551 14399
rect 11253 14365 11287 14399
rect 15301 14365 15335 14399
rect 19717 14365 19751 14399
rect 19901 14365 19935 14399
rect 20637 14365 20671 14399
rect 22293 14365 22327 14399
rect 25237 14365 25271 14399
rect 25329 14365 25363 14399
rect 26249 14365 26283 14399
rect 2329 14297 2363 14331
rect 6929 14297 6963 14331
rect 9505 14297 9539 14331
rect 19165 14297 19199 14331
rect 24593 14297 24627 14331
rect 1593 14229 1627 14263
rect 5641 14229 5675 14263
rect 6561 14229 6595 14263
rect 9137 14229 9171 14263
rect 9873 14229 9907 14263
rect 14657 14229 14691 14263
rect 20361 14229 20395 14263
rect 24225 14229 24259 14263
rect 25789 14229 25823 14263
rect 2421 14025 2455 14059
rect 2697 14025 2731 14059
rect 3433 14025 3467 14059
rect 11253 14025 11287 14059
rect 12449 14025 12483 14059
rect 16957 14025 16991 14059
rect 17417 14025 17451 14059
rect 17785 14025 17819 14059
rect 18337 14025 18371 14059
rect 19073 14025 19107 14059
rect 19349 14025 19383 14059
rect 20821 14025 20855 14059
rect 21465 14025 21499 14059
rect 21925 14025 21959 14059
rect 22937 14025 22971 14059
rect 23489 14025 23523 14059
rect 23673 14025 23707 14059
rect 25421 14025 25455 14059
rect 26249 14025 26283 14059
rect 2237 13889 2271 13923
rect 1961 13753 1995 13787
rect 3341 13957 3375 13991
rect 4997 13957 5031 13991
rect 8401 13957 8435 13991
rect 11989 13957 12023 13991
rect 14013 13957 14047 13991
rect 15945 13957 15979 13991
rect 3893 13889 3927 13923
rect 3985 13889 4019 13923
rect 4905 13889 4939 13923
rect 5457 13889 5491 13923
rect 5641 13889 5675 13923
rect 6009 13889 6043 13923
rect 13093 13889 13127 13923
rect 13461 13889 13495 13923
rect 14473 13889 14507 13923
rect 14565 13889 14599 13923
rect 15393 13889 15427 13923
rect 16589 13889 16623 13923
rect 4537 13821 4571 13855
rect 5365 13821 5399 13855
rect 7021 13821 7055 13855
rect 7277 13821 7311 13855
rect 9045 13821 9079 13855
rect 9781 13821 9815 13855
rect 9873 13821 9907 13855
rect 12909 13821 12943 13855
rect 13921 13821 13955 13855
rect 15761 13821 15795 13855
rect 16405 13821 16439 13855
rect 19165 13957 19199 13991
rect 24777 13957 24811 13991
rect 22477 13889 22511 13923
rect 24133 13889 24167 13923
rect 24225 13889 24259 13923
rect 19165 13821 19199 13855
rect 19441 13821 19475 13855
rect 21741 13821 21775 13855
rect 25237 13821 25271 13855
rect 25789 13821 25823 13855
rect 9413 13753 9447 13787
rect 10118 13753 10152 13787
rect 12817 13753 12851 13787
rect 14381 13753 14415 13787
rect 18889 13753 18923 13787
rect 19073 13753 19107 13787
rect 19708 13753 19742 13787
rect 22293 13753 22327 13787
rect 1593 13685 1627 13719
rect 2053 13685 2087 13719
rect 2421 13685 2455 13719
rect 3801 13685 3835 13719
rect 6561 13685 6595 13719
rect 15025 13685 15059 13719
rect 16313 13685 16347 13719
rect 18429 13685 18463 13719
rect 22385 13685 22419 13719
rect 24041 13685 24075 13719
rect 2237 13481 2271 13515
rect 2329 13481 2363 13515
rect 3617 13481 3651 13515
rect 4813 13481 4847 13515
rect 5273 13481 5307 13515
rect 7757 13481 7791 13515
rect 8309 13481 8343 13515
rect 8677 13481 8711 13515
rect 9045 13481 9079 13515
rect 9505 13481 9539 13515
rect 9689 13481 9723 13515
rect 11253 13481 11287 13515
rect 11621 13481 11655 13515
rect 12725 13481 12759 13515
rect 13185 13481 13219 13515
rect 13921 13481 13955 13515
rect 14197 13481 14231 13515
rect 17049 13481 17083 13515
rect 19073 13481 19107 13515
rect 19533 13481 19567 13515
rect 22845 13481 22879 13515
rect 23305 13481 23339 13515
rect 23397 13481 23431 13515
rect 24501 13481 24535 13515
rect 25145 13481 25179 13515
rect 25881 13481 25915 13515
rect 26249 13481 26283 13515
rect 1685 13413 1719 13447
rect 3249 13413 3283 13447
rect 4353 13413 4387 13447
rect 11161 13413 11195 13447
rect 17325 13413 17359 13447
rect 20085 13413 20119 13447
rect 2881 13345 2915 13379
rect 5181 13345 5215 13379
rect 6633 13345 6667 13379
rect 10057 13345 10091 13379
rect 11713 13345 11747 13379
rect 16313 13345 16347 13379
rect 17877 13345 17911 13379
rect 19441 13345 19475 13379
rect 21180 13345 21214 13379
rect 23765 13345 23799 13379
rect 23857 13345 23891 13379
rect 24961 13345 24995 13379
rect 2421 13277 2455 13311
rect 5365 13277 5399 13311
rect 6377 13277 6411 13311
rect 10149 13277 10183 13311
rect 10241 13277 10275 13311
rect 10701 13277 10735 13311
rect 11805 13277 11839 13311
rect 12357 13277 12391 13311
rect 13277 13277 13311 13311
rect 13461 13277 13495 13311
rect 14933 13277 14967 13311
rect 16405 13277 16439 13311
rect 16497 13277 16531 13311
rect 17969 13277 18003 13311
rect 18153 13277 18187 13311
rect 18981 13277 19015 13311
rect 19717 13277 19751 13311
rect 20913 13277 20947 13311
rect 24041 13277 24075 13311
rect 4629 13209 4663 13243
rect 17509 13209 17543 13243
rect 18613 13209 18647 13243
rect 1869 13141 1903 13175
rect 5917 13141 5951 13175
rect 6193 13141 6227 13175
rect 12817 13141 12851 13175
rect 14657 13141 14691 13175
rect 15761 13141 15795 13175
rect 15945 13141 15979 13175
rect 20729 13141 20763 13175
rect 22293 13141 22327 13175
rect 24869 13141 24903 13175
rect 25513 13141 25547 13175
rect 1869 12937 1903 12971
rect 2053 12937 2087 12971
rect 3065 12937 3099 12971
rect 4721 12937 4755 12971
rect 9505 12937 9539 12971
rect 9965 12937 9999 12971
rect 11621 12937 11655 12971
rect 12909 12937 12943 12971
rect 14381 12937 14415 12971
rect 16129 12937 16163 12971
rect 18429 12937 18463 12971
rect 18797 12937 18831 12971
rect 21373 12937 21407 12971
rect 22753 12937 22787 12971
rect 23489 12937 23523 12971
rect 23673 12937 23707 12971
rect 25421 12937 25455 12971
rect 3433 12869 3467 12903
rect 3617 12869 3651 12903
rect 8401 12869 8435 12903
rect 15669 12869 15703 12903
rect 17509 12869 17543 12903
rect 21005 12869 21039 12903
rect 23029 12869 23063 12903
rect 23213 12869 23247 12903
rect 25053 12869 25087 12903
rect 2605 12801 2639 12835
rect 4169 12801 4203 12835
rect 5825 12801 5859 12835
rect 7389 12801 7423 12835
rect 8953 12801 8987 12835
rect 10609 12801 10643 12835
rect 13461 12801 13495 12835
rect 13645 12801 13679 12835
rect 15117 12801 15151 12835
rect 16681 12801 16715 12835
rect 16773 12801 16807 12835
rect 21833 12801 21867 12835
rect 21925 12801 21959 12835
rect 3985 12733 4019 12767
rect 5549 12733 5583 12767
rect 7849 12733 7883 12767
rect 8309 12733 8343 12767
rect 8769 12733 8803 12767
rect 12173 12733 12207 12767
rect 14013 12733 14047 12767
rect 15025 12733 15059 12767
rect 16589 12733 16623 12767
rect 18889 12733 18923 12767
rect 4077 12665 4111 12699
rect 5089 12665 5123 12699
rect 7205 12665 7239 12699
rect 9873 12665 9907 12699
rect 10425 12665 10459 12699
rect 11345 12665 11379 12699
rect 14933 12665 14967 12699
rect 19156 12665 19190 12699
rect 21741 12665 21775 12699
rect 24133 12801 24167 12835
rect 24225 12801 24259 12835
rect 25237 12733 25271 12767
rect 25789 12733 25823 12767
rect 2421 12597 2455 12631
rect 2513 12597 2547 12631
rect 5181 12597 5215 12631
rect 5641 12597 5675 12631
rect 6377 12597 6411 12631
rect 6837 12597 6871 12631
rect 7297 12597 7331 12631
rect 8861 12597 8895 12631
rect 10333 12597 10367 12631
rect 13001 12597 13035 12631
rect 13369 12597 13403 12631
rect 14565 12597 14599 12631
rect 16221 12597 16255 12631
rect 20269 12597 20303 12631
rect 23213 12597 23247 12631
rect 24041 12597 24075 12631
rect 2145 12393 2179 12427
rect 4261 12393 4295 12427
rect 6469 12393 6503 12427
rect 7021 12393 7055 12427
rect 9045 12393 9079 12427
rect 9413 12393 9447 12427
rect 10057 12393 10091 12427
rect 10333 12393 10367 12427
rect 11437 12393 11471 12427
rect 11713 12393 11747 12427
rect 14657 12393 14691 12427
rect 15117 12393 15151 12427
rect 16037 12393 16071 12427
rect 17601 12393 17635 12427
rect 18981 12393 19015 12427
rect 19073 12393 19107 12427
rect 19441 12393 19475 12427
rect 21373 12393 21407 12427
rect 21833 12393 21867 12427
rect 22845 12393 22879 12427
rect 23397 12393 23431 12427
rect 23765 12393 23799 12427
rect 23857 12393 23891 12427
rect 24501 12393 24535 12427
rect 25145 12393 25179 12427
rect 2789 12325 2823 12359
rect 2881 12325 2915 12359
rect 7481 12325 7515 12359
rect 20729 12325 20763 12359
rect 23305 12325 23339 12359
rect 3525 12257 3559 12291
rect 4077 12257 4111 12291
rect 5825 12257 5859 12291
rect 5917 12257 5951 12291
rect 6285 12257 6319 12291
rect 7389 12257 7423 12291
rect 10701 12257 10735 12291
rect 12164 12257 12198 12291
rect 16589 12257 16623 12291
rect 22201 12257 22235 12291
rect 24961 12257 24995 12291
rect 25605 12257 25639 12291
rect 1409 12189 1443 12223
rect 3065 12189 3099 12223
rect 6009 12189 6043 12223
rect 7573 12189 7607 12223
rect 8401 12189 8435 12223
rect 8585 12189 8619 12223
rect 10793 12189 10827 12223
rect 10977 12189 11011 12223
rect 11897 12189 11931 12223
rect 16681 12189 16715 12223
rect 16865 12189 16899 12223
rect 18061 12189 18095 12223
rect 19533 12189 19567 12223
rect 19717 12189 19751 12223
rect 22293 12189 22327 12223
rect 22477 12189 22511 12223
rect 24041 12189 24075 12223
rect 24869 12189 24903 12223
rect 2421 12121 2455 12155
rect 5181 12121 5215 12155
rect 5457 12121 5491 12155
rect 6285 12121 6319 12155
rect 17969 12121 18003 12155
rect 18613 12121 18647 12155
rect 3893 12053 3927 12087
rect 4629 12053 4663 12087
rect 6837 12053 6871 12087
rect 8033 12053 8067 12087
rect 13277 12053 13311 12087
rect 13829 12053 13863 12087
rect 14197 12053 14231 12087
rect 15577 12053 15611 12087
rect 16221 12053 16255 12087
rect 20361 12053 20395 12087
rect 2605 11849 2639 11883
rect 5825 11849 5859 11883
rect 8217 11849 8251 11883
rect 8769 11849 8803 11883
rect 9137 11849 9171 11883
rect 14933 11849 14967 11883
rect 15301 11849 15335 11883
rect 17877 11849 17911 11883
rect 20913 11849 20947 11883
rect 21833 11849 21867 11883
rect 22937 11849 22971 11883
rect 23489 11849 23523 11883
rect 24961 11849 24995 11883
rect 25421 11849 25455 11883
rect 25881 11849 25915 11883
rect 26249 11781 26283 11815
rect 2237 11713 2271 11747
rect 15485 11713 15519 11747
rect 18061 11713 18095 11747
rect 20453 11713 20487 11747
rect 21281 11713 21315 11747
rect 21649 11713 21683 11747
rect 22385 11713 22419 11747
rect 24225 11713 24259 11747
rect 1961 11645 1995 11679
rect 2053 11645 2087 11679
rect 3065 11645 3099 11679
rect 3157 11645 3191 11679
rect 5641 11645 5675 11679
rect 6653 11645 6687 11679
rect 6837 11645 6871 11679
rect 9873 11645 9907 11679
rect 10140 11645 10174 11679
rect 13001 11645 13035 11679
rect 20729 11645 20763 11679
rect 25237 11645 25271 11679
rect 3424 11577 3458 11611
rect 5089 11577 5123 11611
rect 7082 11577 7116 11611
rect 9781 11577 9815 11611
rect 13246 11577 13280 11611
rect 15730 11577 15764 11611
rect 18306 11577 18340 11611
rect 19993 11577 20027 11611
rect 22293 11577 22327 11611
rect 1593 11509 1627 11543
rect 4537 11509 4571 11543
rect 5549 11509 5583 11543
rect 6193 11509 6227 11543
rect 11253 11509 11287 11543
rect 11989 11509 12023 11543
rect 12909 11509 12943 11543
rect 14381 11509 14415 11543
rect 16865 11509 16899 11543
rect 17417 11509 17451 11543
rect 19441 11509 19475 11543
rect 22201 11509 22235 11543
rect 23673 11509 23707 11543
rect 24041 11509 24075 11543
rect 24133 11509 24167 11543
rect 1961 11305 1995 11339
rect 2237 11305 2271 11339
rect 2881 11305 2915 11339
rect 3433 11305 3467 11339
rect 4353 11305 4387 11339
rect 6377 11305 6411 11339
rect 6929 11305 6963 11339
rect 7205 11305 7239 11339
rect 7665 11305 7699 11339
rect 8217 11305 8251 11339
rect 9321 11305 9355 11339
rect 9873 11305 9907 11339
rect 10333 11305 10367 11339
rect 11805 11305 11839 11339
rect 12357 11305 12391 11339
rect 12725 11305 12759 11339
rect 13001 11305 13035 11339
rect 13369 11305 13403 11339
rect 14381 11305 14415 11339
rect 15485 11305 15519 11339
rect 16313 11305 16347 11339
rect 17877 11305 17911 11339
rect 18981 11305 19015 11339
rect 20913 11305 20947 11339
rect 21281 11305 21315 11339
rect 22017 11305 22051 11339
rect 22477 11305 22511 11339
rect 24041 11305 24075 11339
rect 24777 11305 24811 11339
rect 25145 11305 25179 11339
rect 2789 11237 2823 11271
rect 10692 11237 10726 11271
rect 15945 11237 15979 11271
rect 16764 11237 16798 11271
rect 22385 11237 22419 11271
rect 24409 11237 24443 11271
rect 4445 11169 4479 11203
rect 4701 11169 4735 11203
rect 8125 11169 8159 11203
rect 10425 11169 10459 11203
rect 15301 11169 15335 11203
rect 19349 11169 19383 11203
rect 20729 11169 20763 11203
rect 22845 11169 22879 11203
rect 24593 11169 24627 11203
rect 1409 11101 1443 11135
rect 3065 11101 3099 11135
rect 8309 11101 8343 11135
rect 13461 11101 13495 11135
rect 13645 11101 13679 11135
rect 14749 11101 14783 11135
rect 16497 11101 16531 11135
rect 19441 11101 19475 11135
rect 19533 11101 19567 11135
rect 21373 11101 21407 11135
rect 21557 11101 21591 11135
rect 22937 11101 22971 11135
rect 23121 11101 23155 11135
rect 23673 11101 23707 11135
rect 25513 11101 25547 11135
rect 2421 11033 2455 11067
rect 5825 11033 5859 11067
rect 7757 11033 7791 11067
rect 18889 11033 18923 11067
rect 3801 10965 3835 10999
rect 9045 10965 9079 10999
rect 14105 10965 14139 10999
rect 18429 10965 18463 10999
rect 20085 10965 20119 10999
rect 1593 10761 1627 10795
rect 2513 10761 2547 10795
rect 4537 10761 4571 10795
rect 4997 10761 5031 10795
rect 6193 10761 6227 10795
rect 6653 10761 6687 10795
rect 7297 10761 7331 10795
rect 10425 10761 10459 10795
rect 11621 10761 11655 10795
rect 11897 10761 11931 10795
rect 13001 10761 13035 10795
rect 13461 10761 13495 10795
rect 19073 10761 19107 10795
rect 19441 10761 19475 10795
rect 19625 10761 19659 10795
rect 22477 10761 22511 10795
rect 23305 10761 23339 10795
rect 23857 10761 23891 10795
rect 24777 10761 24811 10795
rect 25605 10761 25639 10795
rect 5181 10693 5215 10727
rect 8953 10693 8987 10727
rect 2605 10625 2639 10659
rect 5641 10625 5675 10659
rect 5825 10625 5859 10659
rect 7849 10625 7883 10659
rect 9597 10625 9631 10659
rect 10977 10625 11011 10659
rect 11161 10625 11195 10659
rect 13829 10625 13863 10659
rect 13921 10625 13955 10659
rect 16957 10625 16991 10659
rect 17417 10625 17451 10659
rect 18613 10625 18647 10659
rect 20085 10625 20119 10659
rect 20269 10625 20303 10659
rect 21649 10625 21683 10659
rect 21833 10625 21867 10659
rect 1409 10557 1443 10591
rect 2872 10557 2906 10591
rect 5549 10557 5583 10591
rect 7205 10557 7239 10591
rect 7757 10557 7791 10591
rect 10057 10557 10091 10591
rect 16221 10557 16255 10591
rect 16865 10557 16899 10591
rect 2053 10489 2087 10523
rect 9413 10489 9447 10523
rect 14188 10489 14222 10523
rect 15945 10489 15979 10523
rect 16773 10489 16807 10523
rect 17877 10489 17911 10523
rect 18521 10489 18555 10523
rect 21005 10489 21039 10523
rect 21557 10489 21591 10523
rect 22201 10489 22235 10523
rect 22661 10625 22695 10659
rect 22937 10557 22971 10591
rect 24593 10557 24627 10591
rect 25145 10557 25179 10591
rect 3985 10421 4019 10455
rect 7665 10421 7699 10455
rect 8401 10421 8435 10455
rect 8769 10421 8803 10455
rect 9321 10421 9355 10455
rect 10517 10421 10551 10455
rect 10885 10421 10919 10455
rect 12449 10421 12483 10455
rect 15301 10421 15335 10455
rect 16405 10421 16439 10455
rect 18061 10421 18095 10455
rect 18429 10421 18463 10455
rect 19993 10421 20027 10455
rect 21189 10421 21223 10455
rect 22477 10421 22511 10455
rect 24409 10421 24443 10455
rect 1869 10217 1903 10251
rect 2329 10217 2363 10251
rect 2789 10217 2823 10251
rect 5181 10217 5215 10251
rect 5917 10217 5951 10251
rect 6469 10217 6503 10251
rect 9413 10217 9447 10251
rect 9873 10217 9907 10251
rect 10333 10217 10367 10251
rect 11713 10217 11747 10251
rect 11897 10217 11931 10251
rect 13461 10217 13495 10251
rect 14841 10217 14875 10251
rect 15301 10217 15335 10251
rect 15761 10217 15795 10251
rect 16497 10217 16531 10251
rect 19993 10217 20027 10251
rect 20913 10217 20947 10251
rect 21925 10217 21959 10251
rect 22293 10217 22327 10251
rect 22477 10217 22511 10251
rect 23765 10217 23799 10251
rect 24409 10217 24443 10251
rect 24777 10217 24811 10251
rect 25053 10217 25087 10251
rect 25789 10217 25823 10251
rect 3433 10149 3467 10183
rect 3801 10149 3835 10183
rect 4445 10149 4479 10183
rect 10793 10149 10827 10183
rect 12357 10149 12391 10183
rect 13921 10149 13955 10183
rect 19717 10149 19751 10183
rect 20729 10149 20763 10183
rect 22937 10149 22971 10183
rect 2881 10081 2915 10115
rect 4537 10081 4571 10115
rect 5641 10081 5675 10115
rect 8033 10081 8067 10115
rect 10701 10081 10735 10115
rect 12265 10081 12299 10115
rect 13829 10081 13863 10115
rect 14473 10081 14507 10115
rect 15669 10081 15703 10115
rect 17233 10081 17267 10115
rect 18797 10081 18831 10115
rect 18889 10081 18923 10115
rect 21281 10081 21315 10115
rect 23581 10081 23615 10115
rect 24593 10081 24627 10115
rect 3065 10013 3099 10047
rect 4629 10013 4663 10047
rect 6561 10013 6595 10047
rect 6653 10013 6687 10047
rect 8125 10013 8159 10047
rect 8217 10013 8251 10047
rect 10977 10013 11011 10047
rect 12541 10013 12575 10047
rect 14013 10013 14047 10047
rect 15945 10013 15979 10047
rect 17325 10013 17359 10047
rect 17417 10013 17451 10047
rect 18981 10013 19015 10047
rect 21373 10013 21407 10047
rect 21557 10013 21591 10047
rect 23305 10013 23339 10047
rect 6101 9945 6135 9979
rect 7665 9945 7699 9979
rect 11345 9945 11379 9979
rect 13093 9945 13127 9979
rect 25421 9945 25455 9979
rect 2421 9877 2455 9911
rect 4077 9877 4111 9911
rect 7389 9877 7423 9911
rect 9045 9877 9079 9911
rect 16865 9877 16899 9911
rect 18061 9877 18095 9911
rect 18429 9877 18463 9911
rect 24041 9877 24075 9911
rect 2881 9673 2915 9707
rect 5273 9673 5307 9707
rect 5825 9673 5859 9707
rect 6469 9673 6503 9707
rect 10609 9673 10643 9707
rect 11989 9673 12023 9707
rect 17785 9673 17819 9707
rect 19073 9673 19107 9707
rect 20913 9673 20947 9707
rect 22293 9673 22327 9707
rect 22661 9673 22695 9707
rect 23489 9673 23523 9707
rect 23857 9673 23891 9707
rect 24685 9673 24719 9707
rect 1777 9605 1811 9639
rect 4721 9605 4755 9639
rect 11161 9605 11195 9639
rect 11529 9605 11563 9639
rect 12909 9605 12943 9639
rect 15853 9605 15887 9639
rect 19625 9605 19659 9639
rect 22937 9605 22971 9639
rect 24961 9605 24995 9639
rect 2421 9537 2455 9571
rect 7205 9537 7239 9571
rect 8217 9537 8251 9571
rect 15485 9537 15519 9571
rect 16497 9537 16531 9571
rect 18613 9537 18647 9571
rect 19441 9537 19475 9571
rect 20269 9537 20303 9571
rect 21741 9537 21775 9571
rect 22385 9537 22419 9571
rect 25329 9537 25363 9571
rect 1685 9469 1719 9503
rect 3249 9469 3283 9503
rect 3341 9469 3375 9503
rect 8033 9469 8067 9503
rect 9229 9469 9263 9503
rect 9496 9469 9530 9503
rect 13461 9469 13495 9503
rect 16405 9469 16439 9503
rect 18429 9469 18463 9503
rect 19993 9469 20027 9503
rect 21649 9469 21683 9503
rect 2145 9401 2179 9435
rect 3586 9401 3620 9435
rect 8125 9401 8159 9435
rect 8677 9401 8711 9435
rect 13706 9401 13740 9435
rect 17417 9401 17451 9435
rect 18521 9401 18555 9435
rect 20085 9401 20119 9435
rect 21557 9401 21591 9435
rect 23673 9469 23707 9503
rect 24133 9469 24167 9503
rect 25697 9469 25731 9503
rect 2237 9333 2271 9367
rect 6101 9333 6135 9367
rect 7481 9333 7515 9367
rect 7665 9333 7699 9367
rect 9045 9333 9079 9367
rect 12449 9333 12483 9367
rect 13277 9333 13311 9367
rect 14841 9333 14875 9367
rect 15945 9333 15979 9367
rect 16313 9333 16347 9367
rect 17049 9333 17083 9367
rect 18061 9333 18095 9367
rect 21189 9333 21223 9367
rect 22385 9333 22419 9367
rect 26065 9333 26099 9367
rect 26433 9333 26467 9367
rect 2421 9129 2455 9163
rect 4353 9129 4387 9163
rect 4905 9129 4939 9163
rect 8493 9129 8527 9163
rect 9321 9129 9355 9163
rect 9873 9129 9907 9163
rect 10333 9129 10367 9163
rect 10793 9129 10827 9163
rect 13185 9129 13219 9163
rect 14013 9129 14047 9163
rect 14105 9129 14139 9163
rect 15117 9129 15151 9163
rect 17325 9129 17359 9163
rect 18797 9129 18831 9163
rect 20269 9129 20303 9163
rect 20729 9129 20763 9163
rect 21925 9129 21959 9163
rect 23305 9129 23339 9163
rect 24317 9129 24351 9163
rect 25053 9129 25087 9163
rect 25421 9129 25455 9163
rect 25789 9129 25823 9163
rect 26249 9129 26283 9163
rect 4813 9061 4847 9095
rect 5825 9061 5859 9095
rect 8769 9061 8803 9095
rect 11152 9061 11186 9095
rect 15568 9061 15602 9095
rect 24685 9061 24719 9095
rect 1409 8993 1443 9027
rect 2789 8993 2823 9027
rect 6725 8993 6759 9027
rect 9689 8993 9723 9027
rect 18153 8993 18187 9027
rect 19165 8993 19199 9027
rect 19717 8993 19751 9027
rect 21281 8993 21315 9027
rect 22477 8993 22511 9027
rect 23489 8993 23523 9027
rect 2881 8925 2915 8959
rect 3065 8925 3099 8959
rect 3525 8925 3559 8959
rect 3893 8925 3927 8959
rect 5089 8925 5123 8959
rect 6469 8925 6503 8959
rect 10885 8925 10919 8959
rect 14197 8925 14231 8959
rect 15301 8925 15335 8959
rect 18245 8925 18279 8959
rect 18337 8925 18371 8959
rect 21373 8925 21407 8959
rect 21465 8925 21499 8959
rect 22201 8925 22235 8959
rect 1961 8857 1995 8891
rect 2329 8857 2363 8891
rect 13645 8857 13679 8891
rect 17785 8857 17819 8891
rect 19625 8857 19659 8891
rect 4445 8789 4479 8823
rect 5549 8789 5583 8823
rect 6285 8789 6319 8823
rect 7849 8789 7883 8823
rect 12265 8789 12299 8823
rect 13461 8789 13495 8823
rect 14749 8789 14783 8823
rect 16681 8789 16715 8823
rect 17601 8789 17635 8823
rect 19901 8789 19935 8823
rect 20913 8789 20947 8823
rect 22109 8789 22143 8823
rect 22293 8789 22327 8823
rect 22661 8789 22695 8823
rect 22937 8789 22971 8823
rect 23673 8789 23707 8823
rect 23949 8789 23983 8823
rect 1501 8585 1535 8619
rect 4169 8585 4203 8619
rect 5733 8585 5767 8619
rect 6009 8585 6043 8619
rect 9137 8585 9171 8619
rect 10241 8585 10275 8619
rect 12081 8585 12115 8619
rect 14657 8585 14691 8619
rect 15761 8585 15795 8619
rect 20085 8585 20119 8619
rect 20545 8585 20579 8619
rect 21557 8585 21591 8619
rect 22753 8585 22787 8619
rect 23029 8585 23063 8619
rect 23489 8585 23523 8619
rect 24133 8585 24167 8619
rect 25237 8585 25271 8619
rect 25697 8585 25731 8619
rect 25973 8585 26007 8619
rect 26341 8585 26375 8619
rect 2605 8517 2639 8551
rect 4629 8517 4663 8551
rect 19441 8517 19475 8551
rect 20453 8517 20487 8551
rect 22293 8517 22327 8551
rect 24961 8517 24995 8551
rect 1961 8449 1995 8483
rect 2053 8449 2087 8483
rect 3709 8449 3743 8483
rect 4537 8449 4571 8483
rect 5181 8449 5215 8483
rect 10701 8449 10735 8483
rect 10885 8449 10919 8483
rect 13093 8449 13127 8483
rect 13277 8449 13311 8483
rect 15669 8449 15703 8483
rect 16221 8449 16255 8483
rect 16313 8449 16347 8483
rect 21005 8449 21039 8483
rect 21097 8449 21131 8483
rect 1869 8381 1903 8415
rect 2973 8381 3007 8415
rect 3433 8381 3467 8415
rect 3525 8381 3559 8415
rect 4997 8381 5031 8415
rect 6561 8381 6595 8415
rect 7665 8381 7699 8415
rect 7757 8381 7791 8415
rect 9781 8381 9815 8415
rect 17785 8381 17819 8415
rect 18061 8381 18095 8415
rect 20913 8381 20947 8415
rect 22109 8381 22143 8415
rect 23673 8381 23707 8415
rect 24501 8381 24535 8415
rect 8002 8313 8036 8347
rect 10149 8313 10183 8347
rect 10609 8313 10643 8347
rect 12817 8313 12851 8347
rect 13544 8313 13578 8347
rect 15209 8313 15243 8347
rect 16129 8313 16163 8347
rect 18306 8313 18340 8347
rect 3065 8245 3099 8279
rect 5089 8245 5123 8279
rect 7021 8245 7055 8279
rect 11345 8245 11379 8279
rect 11713 8245 11747 8279
rect 16773 8245 16807 8279
rect 17417 8245 17451 8279
rect 21925 8245 21959 8279
rect 23857 8245 23891 8279
rect 2237 8041 2271 8075
rect 2789 8041 2823 8075
rect 4261 8041 4295 8075
rect 4721 8041 4755 8075
rect 5089 8041 5123 8075
rect 10517 8041 10551 8075
rect 11621 8041 11655 8075
rect 14105 8041 14139 8075
rect 15117 8041 15151 8075
rect 17785 8041 17819 8075
rect 19165 8041 19199 8075
rect 20729 8041 20763 8075
rect 22937 8041 22971 8075
rect 24593 8041 24627 8075
rect 25053 8041 25087 8075
rect 2881 7973 2915 8007
rect 5632 7973 5666 8007
rect 8493 7973 8527 8007
rect 10057 7973 10091 8007
rect 10885 7973 10919 8007
rect 15546 7973 15580 8007
rect 17601 7973 17635 8007
rect 18613 7973 18647 8007
rect 4077 7905 4111 7939
rect 5365 7905 5399 7939
rect 7481 7905 7515 7939
rect 8401 7905 8435 7939
rect 12337 7905 12371 7939
rect 18153 7905 18187 7939
rect 2973 7837 3007 7871
rect 3525 7837 3559 7871
rect 7849 7837 7883 7871
rect 8585 7837 8619 7871
rect 10333 7837 10367 7871
rect 10977 7837 11011 7871
rect 11069 7837 11103 7871
rect 12081 7837 12115 7871
rect 15301 7837 15335 7871
rect 18245 7837 18279 7871
rect 18337 7837 18371 7871
rect 1869 7769 1903 7803
rect 11897 7769 11931 7803
rect 19349 7905 19383 7939
rect 21281 7905 21315 7939
rect 22845 7905 22879 7939
rect 24041 7905 24075 7939
rect 25145 7905 25179 7939
rect 18797 7837 18831 7871
rect 20269 7837 20303 7871
rect 21373 7837 21407 7871
rect 21557 7837 21591 7871
rect 23029 7837 23063 7871
rect 26065 7837 26099 7871
rect 19901 7769 19935 7803
rect 22477 7769 22511 7803
rect 2421 7701 2455 7735
rect 3893 7701 3927 7735
rect 6745 7701 6779 7735
rect 8033 7701 8067 7735
rect 9321 7701 9355 7735
rect 13461 7701 13495 7735
rect 14473 7701 14507 7735
rect 16681 7701 16715 7735
rect 17233 7701 17267 7735
rect 18613 7701 18647 7735
rect 19533 7701 19567 7735
rect 20913 7701 20947 7735
rect 21925 7701 21959 7735
rect 22385 7701 22419 7735
rect 23489 7701 23523 7735
rect 23857 7701 23891 7735
rect 24225 7701 24259 7735
rect 25329 7701 25363 7735
rect 25697 7701 25731 7735
rect 3157 7497 3191 7531
rect 6101 7497 6135 7531
rect 8217 7497 8251 7531
rect 10793 7497 10827 7531
rect 11897 7497 11931 7531
rect 18061 7497 18095 7531
rect 19349 7497 19383 7531
rect 19625 7497 19659 7531
rect 21189 7497 21223 7531
rect 22937 7497 22971 7531
rect 24593 7497 24627 7531
rect 25329 7497 25363 7531
rect 25697 7497 25731 7531
rect 2697 7429 2731 7463
rect 3065 7429 3099 7463
rect 4537 7429 4571 7463
rect 7113 7429 7147 7463
rect 8585 7429 8619 7463
rect 12449 7429 12483 7463
rect 17141 7429 17175 7463
rect 21097 7429 21131 7463
rect 2053 7361 2087 7395
rect 2237 7361 2271 7395
rect 3709 7361 3743 7395
rect 5181 7361 5215 7395
rect 5273 7361 5307 7395
rect 6653 7361 6687 7395
rect 7757 7361 7791 7395
rect 9781 7361 9815 7395
rect 11345 7361 11379 7395
rect 13093 7361 13127 7395
rect 14565 7361 14599 7395
rect 16129 7361 16163 7395
rect 16589 7361 16623 7395
rect 18613 7361 18647 7395
rect 20177 7361 20211 7395
rect 21649 7361 21683 7395
rect 21741 7361 21775 7395
rect 24225 7361 24259 7395
rect 1961 7293 1995 7327
rect 3617 7293 3651 7327
rect 5825 7293 5859 7327
rect 7573 7293 7607 7327
rect 11161 7293 11195 7327
rect 14473 7293 14507 7327
rect 15117 7293 15151 7327
rect 16037 7293 16071 7327
rect 20085 7293 20119 7327
rect 21557 7293 21591 7327
rect 23673 7293 23707 7327
rect 24777 7293 24811 7327
rect 5089 7225 5123 7259
rect 7481 7225 7515 7259
rect 9137 7225 9171 7259
rect 9597 7225 9631 7259
rect 10333 7225 10367 7259
rect 12265 7225 12299 7259
rect 12817 7225 12851 7259
rect 15485 7225 15519 7259
rect 15945 7225 15979 7259
rect 17877 7225 17911 7259
rect 22569 7225 22603 7259
rect 1593 7157 1627 7191
rect 3525 7157 3559 7191
rect 4169 7157 4203 7191
rect 4721 7157 4755 7191
rect 9229 7157 9263 7191
rect 9689 7157 9723 7191
rect 10701 7157 10735 7191
rect 11253 7157 11287 7191
rect 12909 7157 12943 7191
rect 13461 7157 13495 7191
rect 13829 7157 13863 7191
rect 14013 7157 14047 7191
rect 14381 7157 14415 7191
rect 15577 7157 15611 7191
rect 17509 7157 17543 7191
rect 18429 7157 18463 7191
rect 18521 7157 18555 7191
rect 19993 7157 20027 7191
rect 20729 7157 20763 7191
rect 23305 7157 23339 7191
rect 23857 7157 23891 7191
rect 24961 7157 24995 7191
rect 26157 7157 26191 7191
rect 26433 7157 26467 7191
rect 1685 6953 1719 6987
rect 2789 6953 2823 6987
rect 4077 6953 4111 6987
rect 4445 6953 4479 6987
rect 6469 6953 6503 6987
rect 9321 6953 9355 6987
rect 11805 6953 11839 6987
rect 12541 6953 12575 6987
rect 14013 6953 14047 6987
rect 21281 6953 21315 6987
rect 22477 6953 22511 6987
rect 22845 6953 22879 6987
rect 24777 6953 24811 6987
rect 2881 6885 2915 6919
rect 13277 6885 13311 6919
rect 19441 6885 19475 6919
rect 19901 6885 19935 6919
rect 4537 6817 4571 6851
rect 7665 6817 7699 6851
rect 8125 6817 8159 6851
rect 8217 6817 8251 6851
rect 10333 6817 10367 6851
rect 10681 6817 10715 6851
rect 15025 6817 15059 6851
rect 15485 6817 15519 6851
rect 16497 6817 16531 6851
rect 16856 6817 16890 6851
rect 2973 6749 3007 6783
rect 4629 6749 4663 6783
rect 5273 6749 5307 6783
rect 6561 6749 6595 6783
rect 6653 6749 6687 6783
rect 8309 6749 8343 6783
rect 8769 6749 8803 6783
rect 10425 6749 10459 6783
rect 13369 6749 13403 6783
rect 13553 6749 13587 6783
rect 16589 6749 16623 6783
rect 18613 6749 18647 6783
rect 19533 6749 19567 6783
rect 19717 6749 19751 6783
rect 2421 6681 2455 6715
rect 3801 6681 3835 6715
rect 5917 6681 5951 6715
rect 6101 6681 6135 6715
rect 7757 6681 7791 6715
rect 14381 6681 14415 6715
rect 18889 6681 18923 6715
rect 24041 6817 24075 6851
rect 25145 6817 25179 6851
rect 21373 6749 21407 6783
rect 21465 6749 21499 6783
rect 22937 6749 22971 6783
rect 23121 6749 23155 6783
rect 25697 6749 25731 6783
rect 20913 6681 20947 6715
rect 21925 6681 21959 6715
rect 2329 6613 2363 6647
rect 3433 6613 3467 6647
rect 5549 6613 5583 6647
rect 7297 6613 7331 6647
rect 9873 6613 9907 6647
rect 12909 6613 12943 6647
rect 15669 6613 15703 6647
rect 16129 6613 16163 6647
rect 17969 6613 18003 6647
rect 19073 6613 19107 6647
rect 19901 6613 19935 6647
rect 20177 6613 20211 6647
rect 20729 6613 20763 6647
rect 22293 6613 22327 6647
rect 23765 6613 23799 6647
rect 24225 6613 24259 6647
rect 25329 6613 25363 6647
rect 26065 6613 26099 6647
rect 2237 6409 2271 6443
rect 3249 6409 3283 6443
rect 6101 6409 6135 6443
rect 6561 6409 6595 6443
rect 7757 6409 7791 6443
rect 10057 6409 10091 6443
rect 10609 6409 10643 6443
rect 15025 6409 15059 6443
rect 15853 6409 15887 6443
rect 16405 6409 16439 6443
rect 18061 6409 18095 6443
rect 22569 6409 22603 6443
rect 22845 6409 22879 6443
rect 24685 6409 24719 6443
rect 25053 6409 25087 6443
rect 25789 6409 25823 6443
rect 5825 6341 5859 6375
rect 10517 6341 10551 6375
rect 14473 6341 14507 6375
rect 17877 6341 17911 6375
rect 21005 6341 21039 6375
rect 1685 6273 1719 6307
rect 2881 6273 2915 6307
rect 6837 6273 6871 6307
rect 11161 6273 11195 6307
rect 11989 6273 12023 6307
rect 16313 6273 16347 6307
rect 17049 6273 17083 6307
rect 18521 6273 18555 6307
rect 18705 6273 18739 6307
rect 19165 6273 19199 6307
rect 20085 6273 20119 6307
rect 20269 6273 20303 6307
rect 21741 6273 21775 6307
rect 24225 6273 24259 6307
rect 2605 6205 2639 6239
rect 3709 6205 3743 6239
rect 3801 6205 3835 6239
rect 4068 6205 4102 6239
rect 7849 6205 7883 6239
rect 10977 6205 11011 6239
rect 13093 6205 13127 6239
rect 13360 6205 13394 6239
rect 16865 6205 16899 6239
rect 18429 6205 18463 6239
rect 21557 6205 21591 6239
rect 24133 6205 24167 6239
rect 25237 6205 25271 6239
rect 8116 6137 8150 6171
rect 11069 6137 11103 6171
rect 16773 6137 16807 6171
rect 19993 6137 20027 6171
rect 23489 6137 23523 6171
rect 24041 6137 24075 6171
rect 2145 6069 2179 6103
rect 2697 6069 2731 6103
rect 5181 6069 5215 6103
rect 7297 6069 7331 6103
rect 9229 6069 9263 6103
rect 11713 6069 11747 6103
rect 12909 6069 12943 6103
rect 15485 6069 15519 6103
rect 17417 6069 17451 6103
rect 19441 6069 19475 6103
rect 19625 6069 19659 6103
rect 21189 6069 21223 6103
rect 21649 6069 21683 6103
rect 23673 6069 23707 6103
rect 25421 6069 25455 6103
rect 26249 6069 26283 6103
rect 2421 5865 2455 5899
rect 2881 5865 2915 5899
rect 4261 5865 4295 5899
rect 4629 5865 4663 5899
rect 5365 5865 5399 5899
rect 5825 5865 5859 5899
rect 6837 5865 6871 5899
rect 8309 5865 8343 5899
rect 8861 5865 8895 5899
rect 11069 5865 11103 5899
rect 12633 5865 12667 5899
rect 14105 5865 14139 5899
rect 14657 5865 14691 5899
rect 15301 5865 15335 5899
rect 15761 5865 15795 5899
rect 16681 5865 16715 5899
rect 19165 5865 19199 5899
rect 21373 5865 21407 5899
rect 21925 5865 21959 5899
rect 22477 5865 22511 5899
rect 22937 5865 22971 5899
rect 24409 5865 24443 5899
rect 25053 5865 25087 5899
rect 5733 5797 5767 5831
rect 7196 5797 7230 5831
rect 9956 5797 9990 5831
rect 11897 5797 11931 5831
rect 12265 5797 12299 5831
rect 17132 5797 17166 5831
rect 19993 5797 20027 5831
rect 21281 5797 21315 5831
rect 23765 5797 23799 5831
rect 26249 5797 26283 5831
rect 2789 5729 2823 5763
rect 4077 5729 4111 5763
rect 12992 5729 13026 5763
rect 15669 5729 15703 5763
rect 16865 5729 16899 5763
rect 19349 5729 19383 5763
rect 20269 5729 20303 5763
rect 22845 5729 22879 5763
rect 24501 5729 24535 5763
rect 2973 5661 3007 5695
rect 3249 5661 3283 5695
rect 3525 5661 3559 5695
rect 5917 5661 5951 5695
rect 6929 5661 6963 5695
rect 9689 5661 9723 5695
rect 12725 5661 12759 5695
rect 15853 5661 15887 5695
rect 21465 5661 21499 5695
rect 23029 5661 23063 5695
rect 24593 5661 24627 5695
rect 4997 5593 5031 5627
rect 15025 5593 15059 5627
rect 18245 5593 18279 5627
rect 20913 5593 20947 5627
rect 22385 5593 22419 5627
rect 24041 5593 24075 5627
rect 25789 5593 25823 5627
rect 1777 5525 1811 5559
rect 2237 5525 2271 5559
rect 3249 5525 3283 5559
rect 3893 5525 3927 5559
rect 6377 5525 6411 5559
rect 9229 5525 9263 5559
rect 19533 5525 19567 5559
rect 20729 5525 20763 5559
rect 25421 5525 25455 5559
rect 2789 5321 2823 5355
rect 3157 5321 3191 5355
rect 6285 5321 6319 5355
rect 7113 5321 7147 5355
rect 7573 5321 7607 5355
rect 8677 5321 8711 5355
rect 10517 5321 10551 5355
rect 12449 5321 12483 5355
rect 13921 5321 13955 5355
rect 15025 5321 15059 5355
rect 16589 5321 16623 5355
rect 17509 5321 17543 5355
rect 19349 5321 19383 5355
rect 20637 5321 20671 5355
rect 21005 5321 21039 5355
rect 22569 5321 22603 5355
rect 22937 5321 22971 5355
rect 23673 5321 23707 5355
rect 24777 5321 24811 5355
rect 25053 5321 25087 5355
rect 25881 5321 25915 5355
rect 1685 5253 1719 5287
rect 7665 5253 7699 5287
rect 16865 5253 16899 5287
rect 17877 5253 17911 5287
rect 19625 5253 19659 5287
rect 2237 5185 2271 5219
rect 5733 5185 5767 5219
rect 8125 5185 8159 5219
rect 8309 5185 8343 5219
rect 10057 5185 10091 5219
rect 11161 5185 11195 5219
rect 11529 5185 11563 5219
rect 12265 5185 12299 5219
rect 13001 5185 13035 5219
rect 16037 5185 16071 5219
rect 18521 5185 18555 5219
rect 18613 5185 18647 5219
rect 20177 5185 20211 5219
rect 21649 5185 21683 5219
rect 21741 5185 21775 5219
rect 23397 5185 23431 5219
rect 24317 5185 24351 5219
rect 2053 5117 2087 5151
rect 2145 5117 2179 5151
rect 3249 5117 3283 5151
rect 3516 5117 3550 5151
rect 8033 5117 8067 5151
rect 12909 5117 12943 5151
rect 14381 5117 14415 5151
rect 15853 5117 15887 5151
rect 20085 5117 20119 5151
rect 21557 5117 21591 5151
rect 24041 5117 24075 5151
rect 25237 5117 25271 5151
rect 10885 5049 10919 5083
rect 12817 5049 12851 5083
rect 15945 5049 15979 5083
rect 19993 5049 20027 5083
rect 24133 5049 24167 5083
rect 26157 5049 26191 5083
rect 4629 4981 4663 5015
rect 5273 4981 5307 5015
rect 5549 4981 5583 5015
rect 6561 4981 6595 5015
rect 9321 4981 9355 5015
rect 9505 4981 9539 5015
rect 10425 4981 10459 5015
rect 10977 4981 11011 5015
rect 13461 4981 13495 5015
rect 14197 4981 14231 5015
rect 14565 4981 14599 5015
rect 15393 4981 15427 5015
rect 15485 4981 15519 5015
rect 18061 4981 18095 5015
rect 18429 4981 18463 5015
rect 21189 4981 21223 5015
rect 25421 4981 25455 5015
rect 2329 4777 2363 4811
rect 2421 4777 2455 4811
rect 2789 4777 2823 4811
rect 8953 4777 8987 4811
rect 10425 4777 10459 4811
rect 10885 4777 10919 4811
rect 11529 4777 11563 4811
rect 13645 4777 13679 4811
rect 14013 4777 14047 4811
rect 15117 4777 15151 4811
rect 18153 4777 18187 4811
rect 20729 4777 20763 4811
rect 21925 4777 21959 4811
rect 22385 4777 22419 4811
rect 23765 4777 23799 4811
rect 24133 4777 24167 4811
rect 3893 4709 3927 4743
rect 4344 4709 4378 4743
rect 6101 4709 6135 4743
rect 9965 4709 9999 4743
rect 13185 4709 13219 4743
rect 19073 4709 19107 4743
rect 22937 4709 22971 4743
rect 25053 4709 25087 4743
rect 2881 4641 2915 4675
rect 6817 4641 6851 4675
rect 10793 4641 10827 4675
rect 12449 4641 12483 4675
rect 13553 4641 13587 4675
rect 16396 4641 16430 4675
rect 18429 4641 18463 4675
rect 18981 4641 19015 4675
rect 21281 4641 21315 4675
rect 22845 4641 22879 4675
rect 24501 4641 24535 4675
rect 3065 4573 3099 4607
rect 4077 4573 4111 4607
rect 6561 4573 6595 4607
rect 11069 4573 11103 4607
rect 12541 4573 12575 4607
rect 12725 4573 12759 4607
rect 14105 4573 14139 4607
rect 14289 4573 14323 4607
rect 16129 4573 16163 4607
rect 19165 4573 19199 4607
rect 19625 4573 19659 4607
rect 21373 4573 21407 4607
rect 21465 4573 21499 4607
rect 23029 4573 23063 4607
rect 6377 4505 6411 4539
rect 11989 4505 12023 4539
rect 25789 4505 25823 4539
rect 1961 4437 1995 4471
rect 3525 4437 3559 4471
rect 5457 4437 5491 4471
rect 7941 4437 7975 4471
rect 8585 4437 8619 4471
rect 9413 4437 9447 4471
rect 10333 4437 10367 4471
rect 12081 4437 12115 4471
rect 14749 4437 14783 4471
rect 15577 4437 15611 4471
rect 16037 4437 16071 4471
rect 17509 4437 17543 4471
rect 18613 4437 18647 4471
rect 19993 4437 20027 4471
rect 20913 4437 20947 4471
rect 22477 4437 22511 4471
rect 24685 4437 24719 4471
rect 25421 4437 25455 4471
rect 26249 4437 26283 4471
rect 2973 4233 3007 4267
rect 3433 4233 3467 4267
rect 19073 4233 19107 4267
rect 19625 4233 19659 4267
rect 22569 4233 22603 4267
rect 24685 4233 24719 4267
rect 24869 4233 24903 4267
rect 1777 4165 1811 4199
rect 14197 4165 14231 4199
rect 2421 4097 2455 4131
rect 3985 4097 4019 4131
rect 4997 4097 5031 4131
rect 5825 4097 5859 4131
rect 9137 4097 9171 4131
rect 9781 4097 9815 4131
rect 9873 4097 9907 4131
rect 11529 4097 11563 4131
rect 13185 4097 13219 4131
rect 13369 4097 13403 4131
rect 14933 4097 14967 4131
rect 15301 4097 15335 4131
rect 16129 4097 16163 4131
rect 16681 4097 16715 4131
rect 16865 4097 16899 4131
rect 17785 4097 17819 4131
rect 18521 4097 18555 4131
rect 18613 4097 18647 4131
rect 20177 4097 20211 4131
rect 21741 4097 21775 4131
rect 24225 4097 24259 4131
rect 2237 4029 2271 4063
rect 2329 4029 2363 4063
rect 5549 4029 5583 4063
rect 6837 4029 6871 4063
rect 9689 4029 9723 4063
rect 12173 4029 12207 4063
rect 13093 4029 13127 4063
rect 13829 4029 13863 4063
rect 14657 4029 14691 4063
rect 16589 4029 16623 4063
rect 17417 4029 17451 4063
rect 18429 4029 18463 4063
rect 20085 4029 20119 4063
rect 21557 4029 21591 4063
rect 24869 4029 24903 4063
rect 25053 4029 25087 4063
rect 25237 4029 25271 4063
rect 25789 4029 25823 4063
rect 3341 3961 3375 3995
rect 3893 3961 3927 3995
rect 5641 3961 5675 3995
rect 7104 3961 7138 3995
rect 14749 3961 14783 3995
rect 21097 3961 21131 3995
rect 21649 3961 21683 3995
rect 24133 3961 24167 3995
rect 26249 3961 26283 3995
rect 1869 3893 1903 3927
rect 3801 3893 3835 3927
rect 4537 3893 4571 3927
rect 5181 3893 5215 3927
rect 6193 3893 6227 3927
rect 6561 3893 6595 3927
rect 8217 3893 8251 3927
rect 8861 3893 8895 3927
rect 9321 3893 9355 3927
rect 10517 3893 10551 3927
rect 10885 3893 10919 3927
rect 11897 3893 11931 3927
rect 12725 3893 12759 3927
rect 14289 3893 14323 3927
rect 15669 3893 15703 3927
rect 16221 3893 16255 3927
rect 18061 3893 18095 3927
rect 19441 3893 19475 3927
rect 19993 3893 20027 3927
rect 20729 3893 20763 3927
rect 21189 3893 21223 3927
rect 22845 3893 22879 3927
rect 23397 3893 23431 3927
rect 23673 3893 23707 3927
rect 24041 3893 24075 3927
rect 25421 3893 25455 3927
rect 2421 3689 2455 3723
rect 3525 3689 3559 3723
rect 4077 3689 4111 3723
rect 4537 3689 4571 3723
rect 5273 3689 5307 3723
rect 9321 3689 9355 3723
rect 9689 3689 9723 3723
rect 10149 3689 10183 3723
rect 10793 3689 10827 3723
rect 13093 3689 13127 3723
rect 13737 3689 13771 3723
rect 14197 3689 14231 3723
rect 15025 3689 15059 3723
rect 16313 3689 16347 3723
rect 17877 3689 17911 3723
rect 18613 3689 18647 3723
rect 18981 3689 19015 3723
rect 19441 3689 19475 3723
rect 20913 3689 20947 3723
rect 21373 3689 21407 3723
rect 24409 3689 24443 3723
rect 2329 3621 2363 3655
rect 5641 3621 5675 3655
rect 11529 3621 11563 3655
rect 14105 3621 14139 3655
rect 17233 3621 17267 3655
rect 17785 3621 17819 3655
rect 19349 3621 19383 3655
rect 23489 3621 23523 3655
rect 25421 3621 25455 3655
rect 1409 3553 1443 3587
rect 1961 3553 1995 3587
rect 2789 3553 2823 3587
rect 4445 3553 4479 3587
rect 5825 3553 5859 3587
rect 6081 3553 6115 3587
rect 8585 3553 8619 3587
rect 10057 3553 10091 3587
rect 11161 3553 11195 3587
rect 11980 3553 12014 3587
rect 16221 3553 16255 3587
rect 21281 3553 21315 3587
rect 22845 3553 22879 3587
rect 24501 3553 24535 3587
rect 26249 3553 26283 3587
rect 2881 3485 2915 3519
rect 2973 3485 3007 3519
rect 3893 3485 3927 3519
rect 4721 3485 4755 3519
rect 10333 3485 10367 3519
rect 11713 3485 11747 3519
rect 14749 3485 14783 3519
rect 16497 3485 16531 3519
rect 16957 3485 16991 3519
rect 17969 3485 18003 3519
rect 19625 3485 19659 3519
rect 21465 3485 21499 3519
rect 21925 3485 21959 3519
rect 22937 3485 22971 3519
rect 23121 3485 23155 3519
rect 24685 3485 24719 3519
rect 7205 3417 7239 3451
rect 22385 3417 22419 3451
rect 24041 3417 24075 3451
rect 25053 3417 25087 3451
rect 1593 3349 1627 3383
rect 7757 3349 7791 3383
rect 8493 3349 8527 3383
rect 8769 3349 8803 3383
rect 15577 3349 15611 3383
rect 15853 3349 15887 3383
rect 17417 3349 17451 3383
rect 19993 3349 20027 3383
rect 20637 3349 20671 3383
rect 22477 3349 22511 3383
rect 23857 3349 23891 3383
rect 25789 3349 25823 3383
rect 2053 3145 2087 3179
rect 3617 3145 3651 3179
rect 4997 3145 5031 3179
rect 5181 3145 5215 3179
rect 10333 3145 10367 3179
rect 11161 3145 11195 3179
rect 12265 3145 12299 3179
rect 14381 3145 14415 3179
rect 16221 3145 16255 3179
rect 17785 3145 17819 3179
rect 19625 3145 19659 3179
rect 21189 3145 21223 3179
rect 22293 3145 22327 3179
rect 23673 3145 23707 3179
rect 24685 3145 24719 3179
rect 4629 3077 4663 3111
rect 6837 3077 6871 3111
rect 10701 3077 10735 3111
rect 17141 3077 17175 3111
rect 23489 3077 23523 3111
rect 1961 3009 1995 3043
rect 2605 3009 2639 3043
rect 3157 3009 3191 3043
rect 4169 3009 4203 3043
rect 5825 3009 5859 3043
rect 7481 3009 7515 3043
rect 13185 3009 13219 3043
rect 13829 3009 13863 3043
rect 18613 3009 18647 3043
rect 19073 3009 19107 3043
rect 20085 3009 20119 3043
rect 20177 3009 20211 3043
rect 21741 3009 21775 3043
rect 22937 3009 22971 3043
rect 24133 3009 24167 3043
rect 24317 3009 24351 3043
rect 26249 3009 26283 3043
rect 2513 2941 2547 2975
rect 3249 2941 3283 2975
rect 3525 2941 3559 2975
rect 4077 2941 4111 2975
rect 6285 2941 6319 2975
rect 7205 2941 7239 2975
rect 8401 2941 8435 2975
rect 8668 2941 8702 2975
rect 11253 2941 11287 2975
rect 14841 2941 14875 2975
rect 15108 2941 15142 2975
rect 16865 2941 16899 2975
rect 18429 2941 18463 2975
rect 18521 2941 18555 2975
rect 19533 2941 19567 2975
rect 19993 2941 20027 2975
rect 21649 2941 21683 2975
rect 25237 2941 25271 2975
rect 25789 2941 25823 2975
rect 2421 2873 2455 2907
rect 5549 2873 5583 2907
rect 7297 2873 7331 2907
rect 12817 2873 12851 2907
rect 13737 2873 13771 2907
rect 20729 2873 20763 2907
rect 21097 2873 21131 2907
rect 21557 2873 21591 2907
rect 3249 2805 3283 2839
rect 3985 2805 4019 2839
rect 5641 2805 5675 2839
rect 6653 2805 6687 2839
rect 7941 2805 7975 2839
rect 8217 2805 8251 2839
rect 9781 2805 9815 2839
rect 11437 2805 11471 2839
rect 11805 2805 11839 2839
rect 13277 2805 13311 2839
rect 13645 2805 13679 2839
rect 14657 2805 14691 2839
rect 18061 2805 18095 2839
rect 22661 2805 22695 2839
rect 24041 2805 24075 2839
rect 25053 2805 25087 2839
rect 25421 2805 25455 2839
rect 2421 2601 2455 2635
rect 2881 2601 2915 2635
rect 5733 2601 5767 2635
rect 6653 2601 6687 2635
rect 8309 2601 8343 2635
rect 14289 2601 14323 2635
rect 14933 2601 14967 2635
rect 18061 2601 18095 2635
rect 18797 2601 18831 2635
rect 21189 2601 21223 2635
rect 22293 2601 22327 2635
rect 24041 2601 24075 2635
rect 2789 2533 2823 2567
rect 3709 2533 3743 2567
rect 7196 2533 7230 2567
rect 10048 2533 10082 2567
rect 12081 2533 12115 2567
rect 13176 2533 13210 2567
rect 15730 2533 15764 2567
rect 21649 2533 21683 2567
rect 24409 2533 24443 2567
rect 1409 2465 1443 2499
rect 4353 2465 4387 2499
rect 4620 2465 4654 2499
rect 6285 2465 6319 2499
rect 6929 2465 6963 2499
rect 8861 2465 8895 2499
rect 9505 2465 9539 2499
rect 9781 2465 9815 2499
rect 12357 2465 12391 2499
rect 12909 2465 12943 2499
rect 15209 2465 15243 2499
rect 15485 2465 15519 2499
rect 18705 2465 18739 2499
rect 19717 2465 19751 2499
rect 19901 2465 19935 2499
rect 21557 2465 21591 2499
rect 22753 2465 22787 2499
rect 23397 2465 23431 2499
rect 23673 2465 23707 2499
rect 24501 2465 24535 2499
rect 25605 2465 25639 2499
rect 26065 2465 26099 2499
rect 26433 2465 26467 2499
rect 2329 2397 2363 2431
rect 2973 2397 3007 2431
rect 18889 2397 18923 2431
rect 21741 2397 21775 2431
rect 22569 2397 22603 2431
rect 24593 2397 24627 2431
rect 25053 2397 25087 2431
rect 17693 2329 17727 2363
rect 20545 2329 20579 2363
rect 25421 2329 25455 2363
rect 1593 2261 1627 2295
rect 1961 2261 1995 2295
rect 11161 2261 11195 2295
rect 16865 2261 16899 2295
rect 18337 2261 18371 2295
rect 20085 2261 20119 2295
rect 20913 2261 20947 2295
rect 22937 2261 22971 2295
rect 25789 2261 25823 2295
<< metal1 >>
rect 20714 26800 20720 26852
rect 20772 26840 20778 26852
rect 23750 26840 23756 26852
rect 20772 26812 23756 26840
rect 20772 26800 20778 26812
rect 23750 26800 23756 26812
rect 23808 26800 23814 26852
rect 18506 26664 18512 26716
rect 18564 26704 18570 26716
rect 24762 26704 24768 26716
rect 18564 26676 24768 26704
rect 18564 26664 18570 26676
rect 24762 26664 24768 26676
rect 24820 26664 24826 26716
rect 2685 26571 2743 26577
rect 2685 26537 2697 26571
rect 2731 26568 2743 26571
rect 20346 26568 20352 26580
rect 2731 26540 20352 26568
rect 2731 26537 2743 26540
rect 2685 26531 2743 26537
rect 20346 26528 20352 26540
rect 20404 26528 20410 26580
rect 13538 26460 13544 26512
rect 13596 26500 13602 26512
rect 23290 26500 23296 26512
rect 13596 26472 23296 26500
rect 13596 26460 13602 26472
rect 23290 26460 23296 26472
rect 23348 26460 23354 26512
rect 19337 26367 19395 26373
rect 19337 26364 19349 26367
rect 10684 26336 19349 26364
rect 7374 26120 7380 26172
rect 7432 26160 7438 26172
rect 10684 26160 10712 26336
rect 19337 26333 19349 26336
rect 19383 26333 19395 26367
rect 19337 26327 19395 26333
rect 20438 26256 20444 26308
rect 20496 26296 20502 26308
rect 23750 26296 23756 26308
rect 20496 26268 23756 26296
rect 20496 26256 20502 26268
rect 23750 26256 23756 26268
rect 23808 26256 23814 26308
rect 10778 26188 10784 26240
rect 10836 26228 10842 26240
rect 21358 26228 21364 26240
rect 10836 26200 21364 26228
rect 10836 26188 10842 26200
rect 21358 26188 21364 26200
rect 21416 26188 21422 26240
rect 7432 26132 10712 26160
rect 16853 26163 16911 26169
rect 7432 26120 7438 26132
rect 16853 26129 16865 26163
rect 16899 26160 16911 26163
rect 25038 26160 25044 26172
rect 16899 26132 25044 26160
rect 16899 26129 16911 26132
rect 16853 26123 16911 26129
rect 25038 26120 25044 26132
rect 25096 26120 25102 26172
rect 2682 26092 2688 26104
rect 2643 26064 2688 26092
rect 2682 26052 2688 26064
rect 2740 26052 2746 26104
rect 5166 26052 5172 26104
rect 5224 26092 5230 26104
rect 11425 26095 11483 26101
rect 11425 26092 11437 26095
rect 5224 26064 11437 26092
rect 5224 26052 5230 26064
rect 11425 26061 11437 26064
rect 11471 26061 11483 26095
rect 11425 26055 11483 26061
rect 11514 26052 11520 26104
rect 11572 26092 11578 26104
rect 16669 26095 16727 26101
rect 16669 26092 16681 26095
rect 11572 26064 16681 26092
rect 11572 26052 11578 26064
rect 16669 26061 16681 26064
rect 16715 26061 16727 26095
rect 22922 26092 22928 26104
rect 16669 26055 16727 26061
rect 16776 26064 22928 26092
rect 10870 25984 10876 26036
rect 10928 26024 10934 26036
rect 16776 26024 16804 26064
rect 22922 26052 22928 26064
rect 22980 26052 22986 26104
rect 10928 25996 16804 26024
rect 10928 25984 10934 25996
rect 18414 25984 18420 26036
rect 18472 26024 18478 26036
rect 26602 26024 26608 26036
rect 18472 25996 26608 26024
rect 18472 25984 18478 25996
rect 26602 25984 26608 25996
rect 26660 25984 26666 26036
rect 5074 25916 5080 25968
rect 5132 25956 5138 25968
rect 16853 25959 16911 25965
rect 16853 25956 16865 25959
rect 5132 25928 16865 25956
rect 5132 25916 5138 25928
rect 16853 25925 16865 25928
rect 16899 25925 16911 25959
rect 16853 25919 16911 25925
rect 16942 25916 16948 25968
rect 17000 25956 17006 25968
rect 18230 25956 18236 25968
rect 17000 25928 18236 25956
rect 17000 25916 17006 25928
rect 18230 25916 18236 25928
rect 18288 25916 18294 25968
rect 18322 25916 18328 25968
rect 18380 25956 18386 25968
rect 19242 25956 19248 25968
rect 18380 25928 19248 25956
rect 18380 25916 18386 25928
rect 19242 25916 19248 25928
rect 19300 25916 19306 25968
rect 19337 25959 19395 25965
rect 19337 25925 19349 25959
rect 19383 25956 19395 25959
rect 20898 25956 20904 25968
rect 19383 25928 20904 25956
rect 19383 25925 19395 25928
rect 19337 25919 19395 25925
rect 20898 25916 20904 25928
rect 20956 25916 20962 25968
rect 20990 25916 20996 25968
rect 21048 25956 21054 25968
rect 22738 25956 22744 25968
rect 21048 25928 22744 25956
rect 21048 25916 21054 25928
rect 22738 25916 22744 25928
rect 22796 25916 22802 25968
rect 6822 25848 6828 25900
rect 6880 25888 6886 25900
rect 11698 25888 11704 25900
rect 6880 25860 11704 25888
rect 6880 25848 6886 25860
rect 11698 25848 11704 25860
rect 11756 25848 11762 25900
rect 11793 25891 11851 25897
rect 11793 25857 11805 25891
rect 11839 25888 11851 25891
rect 23750 25888 23756 25900
rect 11839 25860 23756 25888
rect 11839 25857 11851 25860
rect 11793 25851 11851 25857
rect 23750 25848 23756 25860
rect 23808 25848 23814 25900
rect 11330 25780 11336 25832
rect 11388 25820 11394 25832
rect 15381 25823 15439 25829
rect 15381 25820 15393 25823
rect 11388 25792 15393 25820
rect 11388 25780 11394 25792
rect 15381 25789 15393 25792
rect 15427 25789 15439 25823
rect 15381 25783 15439 25789
rect 15562 25780 15568 25832
rect 15620 25820 15626 25832
rect 15620 25792 19012 25820
rect 15620 25780 15626 25792
rect 18874 25752 18880 25764
rect 15120 25724 18880 25752
rect 9950 25644 9956 25696
rect 10008 25684 10014 25696
rect 15120 25684 15148 25724
rect 18874 25712 18880 25724
rect 18932 25712 18938 25764
rect 18984 25752 19012 25792
rect 19978 25780 19984 25832
rect 20036 25820 20042 25832
rect 20714 25820 20720 25832
rect 20036 25792 20720 25820
rect 20036 25780 20042 25792
rect 20714 25780 20720 25792
rect 20772 25780 20778 25832
rect 24578 25752 24584 25764
rect 18984 25724 24584 25752
rect 24578 25712 24584 25724
rect 24636 25712 24642 25764
rect 10008 25656 15148 25684
rect 15381 25687 15439 25693
rect 10008 25644 10014 25656
rect 15381 25653 15393 25687
rect 15427 25684 15439 25687
rect 16666 25684 16672 25696
rect 15427 25656 16672 25684
rect 15427 25653 15439 25656
rect 15381 25647 15439 25653
rect 16666 25644 16672 25656
rect 16724 25644 16730 25696
rect 16761 25687 16819 25693
rect 16761 25653 16773 25687
rect 16807 25684 16819 25687
rect 23474 25684 23480 25696
rect 16807 25656 23480 25684
rect 16807 25653 16819 25656
rect 16761 25647 16819 25653
rect 23474 25644 23480 25656
rect 23532 25644 23538 25696
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 5534 25440 5540 25492
rect 5592 25480 5598 25492
rect 9490 25480 9496 25492
rect 5592 25452 9496 25480
rect 5592 25440 5598 25452
rect 9490 25440 9496 25452
rect 9548 25440 9554 25492
rect 9950 25480 9956 25492
rect 9911 25452 9956 25480
rect 9950 25440 9956 25452
rect 10008 25440 10014 25492
rect 10060 25452 11652 25480
rect 1486 25372 1492 25424
rect 1544 25412 1550 25424
rect 5169 25415 5227 25421
rect 5169 25412 5181 25415
rect 1544 25384 5181 25412
rect 1544 25372 1550 25384
rect 5169 25381 5181 25384
rect 5215 25381 5227 25415
rect 5169 25375 5227 25381
rect 5258 25372 5264 25424
rect 5316 25412 5322 25424
rect 10060 25412 10088 25452
rect 5316 25384 10088 25412
rect 10505 25415 10563 25421
rect 5316 25372 5322 25384
rect 10505 25381 10517 25415
rect 10551 25412 10563 25415
rect 11624 25412 11652 25452
rect 11698 25440 11704 25492
rect 11756 25480 11762 25492
rect 12802 25480 12808 25492
rect 11756 25452 12808 25480
rect 11756 25440 11762 25452
rect 12802 25440 12808 25452
rect 12860 25440 12866 25492
rect 12894 25440 12900 25492
rect 12952 25480 12958 25492
rect 14182 25480 14188 25492
rect 12952 25452 14188 25480
rect 12952 25440 12958 25452
rect 14182 25440 14188 25452
rect 14240 25440 14246 25492
rect 14369 25483 14427 25489
rect 14369 25449 14381 25483
rect 14415 25449 14427 25483
rect 14369 25443 14427 25449
rect 14553 25483 14611 25489
rect 14553 25449 14565 25483
rect 14599 25480 14611 25483
rect 15470 25480 15476 25492
rect 14599 25452 15476 25480
rect 14599 25449 14611 25452
rect 14553 25443 14611 25449
rect 14090 25412 14096 25424
rect 10551 25384 11560 25412
rect 11624 25384 14096 25412
rect 10551 25381 10563 25384
rect 10505 25375 10563 25381
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 2130 25344 2136 25356
rect 1443 25316 2136 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 2130 25304 2136 25316
rect 2188 25304 2194 25356
rect 2498 25344 2504 25356
rect 2459 25316 2504 25344
rect 2498 25304 2504 25316
rect 2556 25304 2562 25356
rect 4062 25344 4068 25356
rect 4023 25316 4068 25344
rect 4062 25304 4068 25316
rect 4120 25304 4126 25356
rect 6546 25304 6552 25356
rect 6604 25344 6610 25356
rect 7929 25347 7987 25353
rect 7929 25344 7941 25347
rect 6604 25316 7941 25344
rect 6604 25304 6610 25316
rect 7929 25313 7941 25316
rect 7975 25313 7987 25347
rect 9766 25344 9772 25356
rect 9727 25316 9772 25344
rect 7929 25307 7987 25313
rect 9766 25304 9772 25316
rect 9824 25304 9830 25356
rect 11330 25344 11336 25356
rect 10796 25316 11336 25344
rect 2222 25236 2228 25288
rect 2280 25276 2286 25288
rect 3789 25279 3847 25285
rect 3789 25276 3801 25279
rect 2280 25248 3801 25276
rect 2280 25236 2286 25248
rect 3789 25245 3801 25248
rect 3835 25245 3847 25279
rect 8021 25279 8079 25285
rect 8021 25276 8033 25279
rect 3789 25239 3847 25245
rect 7392 25248 8033 25276
rect 4338 25168 4344 25220
rect 4396 25208 4402 25220
rect 5166 25208 5172 25220
rect 4396 25180 5172 25208
rect 4396 25168 4402 25180
rect 5166 25168 5172 25180
rect 5224 25168 5230 25220
rect 566 25100 572 25152
rect 624 25140 630 25152
rect 1581 25143 1639 25149
rect 1581 25140 1593 25143
rect 624 25112 1593 25140
rect 624 25100 630 25112
rect 1581 25109 1593 25112
rect 1627 25109 1639 25143
rect 2038 25140 2044 25152
rect 1999 25112 2044 25140
rect 1581 25103 1639 25109
rect 2038 25100 2044 25112
rect 2096 25100 2102 25152
rect 2314 25140 2320 25152
rect 2275 25112 2320 25140
rect 2314 25100 2320 25112
rect 2372 25100 2378 25152
rect 2685 25143 2743 25149
rect 2685 25109 2697 25143
rect 2731 25140 2743 25143
rect 2866 25140 2872 25152
rect 2731 25112 2872 25140
rect 2731 25109 2743 25112
rect 2685 25103 2743 25109
rect 2866 25100 2872 25112
rect 2924 25100 2930 25152
rect 3142 25140 3148 25152
rect 3103 25112 3148 25140
rect 3142 25100 3148 25112
rect 3200 25100 3206 25152
rect 3418 25140 3424 25152
rect 3379 25112 3424 25140
rect 3418 25100 3424 25112
rect 3476 25100 3482 25152
rect 3694 25100 3700 25152
rect 3752 25140 3758 25152
rect 4249 25143 4307 25149
rect 4249 25140 4261 25143
rect 3752 25112 4261 25140
rect 3752 25100 3758 25112
rect 4249 25109 4261 25112
rect 4295 25109 4307 25143
rect 4706 25140 4712 25152
rect 4667 25112 4712 25140
rect 4249 25103 4307 25109
rect 4706 25100 4712 25112
rect 4764 25100 4770 25152
rect 4982 25140 4988 25152
rect 4943 25112 4988 25140
rect 4982 25100 4988 25112
rect 5040 25100 5046 25152
rect 6454 25100 6460 25152
rect 6512 25140 6518 25152
rect 7392 25149 7420 25248
rect 8021 25245 8033 25248
rect 8067 25245 8079 25279
rect 8021 25239 8079 25245
rect 8113 25279 8171 25285
rect 8113 25245 8125 25279
rect 8159 25245 8171 25279
rect 8113 25239 8171 25245
rect 7926 25168 7932 25220
rect 7984 25208 7990 25220
rect 8128 25208 8156 25239
rect 10796 25217 10824 25316
rect 11330 25304 11336 25316
rect 11388 25304 11394 25356
rect 11054 25236 11060 25288
rect 11112 25276 11118 25288
rect 11532 25285 11560 25384
rect 14090 25372 14096 25384
rect 14148 25372 14154 25424
rect 14384 25412 14412 25443
rect 15470 25440 15476 25452
rect 15528 25440 15534 25492
rect 15749 25483 15807 25489
rect 15749 25449 15761 25483
rect 15795 25480 15807 25483
rect 19518 25480 19524 25492
rect 15795 25452 19524 25480
rect 15795 25449 15807 25452
rect 15749 25443 15807 25449
rect 19518 25440 19524 25452
rect 19576 25440 19582 25492
rect 19705 25483 19763 25489
rect 19705 25449 19717 25483
rect 19751 25480 19763 25483
rect 19978 25480 19984 25492
rect 19751 25452 19984 25480
rect 19751 25449 19763 25452
rect 19705 25443 19763 25449
rect 19978 25440 19984 25452
rect 20036 25440 20042 25492
rect 20073 25483 20131 25489
rect 20073 25449 20085 25483
rect 20119 25480 20131 25483
rect 20622 25480 20628 25492
rect 20119 25452 20628 25480
rect 20119 25449 20131 25452
rect 20073 25443 20131 25449
rect 20622 25440 20628 25452
rect 20680 25440 20686 25492
rect 21361 25483 21419 25489
rect 21361 25449 21373 25483
rect 21407 25480 21419 25483
rect 23014 25480 23020 25492
rect 21407 25452 23020 25480
rect 21407 25449 21419 25452
rect 21361 25443 21419 25449
rect 23014 25440 23020 25452
rect 23072 25440 23078 25492
rect 21266 25412 21272 25424
rect 14384 25384 21272 25412
rect 21266 25372 21272 25384
rect 21324 25372 21330 25424
rect 12066 25304 12072 25356
rect 12124 25344 12130 25356
rect 12989 25347 13047 25353
rect 12989 25344 13001 25347
rect 12124 25316 13001 25344
rect 12124 25304 12130 25316
rect 12989 25313 13001 25316
rect 13035 25313 13047 25347
rect 12989 25307 13047 25313
rect 14185 25347 14243 25353
rect 14185 25313 14197 25347
rect 14231 25344 14243 25347
rect 14231 25316 14265 25344
rect 14231 25313 14243 25316
rect 14185 25307 14243 25313
rect 11425 25279 11483 25285
rect 11425 25276 11437 25279
rect 11112 25248 11437 25276
rect 11112 25236 11118 25248
rect 11425 25245 11437 25248
rect 11471 25245 11483 25279
rect 11425 25239 11483 25245
rect 11517 25279 11575 25285
rect 11517 25245 11529 25279
rect 11563 25276 11575 25279
rect 12894 25276 12900 25288
rect 11563 25248 12900 25276
rect 11563 25245 11575 25248
rect 11517 25239 11575 25245
rect 12894 25236 12900 25248
rect 12952 25236 12958 25288
rect 13078 25276 13084 25288
rect 13039 25248 13084 25276
rect 13078 25236 13084 25248
rect 13136 25236 13142 25288
rect 13265 25279 13323 25285
rect 13265 25245 13277 25279
rect 13311 25276 13323 25279
rect 13998 25276 14004 25288
rect 13311 25248 14004 25276
rect 13311 25245 13323 25248
rect 13265 25239 13323 25245
rect 13998 25236 14004 25248
rect 14056 25236 14062 25288
rect 14093 25279 14151 25285
rect 14093 25245 14105 25279
rect 14139 25276 14151 25279
rect 14200 25276 14228 25307
rect 14366 25304 14372 25356
rect 14424 25344 14430 25356
rect 15565 25347 15623 25353
rect 14424 25316 15516 25344
rect 14424 25304 14430 25316
rect 14553 25279 14611 25285
rect 14553 25276 14565 25279
rect 14139 25248 14565 25276
rect 14139 25245 14151 25248
rect 14093 25239 14151 25245
rect 14553 25245 14565 25248
rect 14599 25245 14611 25279
rect 15488 25276 15516 25316
rect 15565 25313 15577 25347
rect 15611 25344 15623 25347
rect 15930 25344 15936 25356
rect 15611 25316 15936 25344
rect 15611 25313 15623 25316
rect 15565 25307 15623 25313
rect 15930 25304 15936 25316
rect 15988 25304 15994 25356
rect 16850 25344 16856 25356
rect 16040 25316 16856 25344
rect 16040 25276 16068 25316
rect 16850 25304 16856 25316
rect 16908 25304 16914 25356
rect 16942 25304 16948 25356
rect 17000 25344 17006 25356
rect 17037 25347 17095 25353
rect 17037 25344 17049 25347
rect 17000 25316 17049 25344
rect 17000 25304 17006 25316
rect 17037 25313 17049 25316
rect 17083 25313 17095 25347
rect 17037 25307 17095 25313
rect 17129 25347 17187 25353
rect 17129 25313 17141 25347
rect 17175 25344 17187 25347
rect 17494 25344 17500 25356
rect 17175 25316 17500 25344
rect 17175 25313 17187 25316
rect 17129 25307 17187 25313
rect 17494 25304 17500 25316
rect 17552 25304 17558 25356
rect 17589 25347 17647 25353
rect 17589 25313 17601 25347
rect 17635 25344 17647 25347
rect 17773 25347 17831 25353
rect 17773 25344 17785 25347
rect 17635 25316 17785 25344
rect 17635 25313 17647 25316
rect 17589 25307 17647 25313
rect 17773 25313 17785 25316
rect 17819 25344 17831 25347
rect 18598 25344 18604 25356
rect 17819 25316 18604 25344
rect 17819 25313 17831 25316
rect 17773 25307 17831 25313
rect 18598 25304 18604 25316
rect 18656 25304 18662 25356
rect 18690 25304 18696 25356
rect 18748 25344 18754 25356
rect 18748 25316 18793 25344
rect 18748 25304 18754 25316
rect 19058 25304 19064 25356
rect 19116 25344 19122 25356
rect 19889 25347 19947 25353
rect 19889 25344 19901 25347
rect 19116 25316 19901 25344
rect 19116 25304 19122 25316
rect 19889 25313 19901 25316
rect 19935 25344 19947 25347
rect 20714 25344 20720 25356
rect 19935 25316 20720 25344
rect 19935 25313 19947 25316
rect 19889 25307 19947 25313
rect 20714 25304 20720 25316
rect 20772 25304 20778 25356
rect 21174 25344 21180 25356
rect 21135 25316 21180 25344
rect 21174 25304 21180 25316
rect 21232 25304 21238 25356
rect 22281 25347 22339 25353
rect 22281 25313 22293 25347
rect 22327 25344 22339 25347
rect 22370 25344 22376 25356
rect 22327 25316 22376 25344
rect 22327 25313 22339 25316
rect 22281 25307 22339 25313
rect 22370 25304 22376 25316
rect 22428 25304 22434 25356
rect 24029 25347 24087 25353
rect 24029 25313 24041 25347
rect 24075 25344 24087 25347
rect 24210 25344 24216 25356
rect 24075 25316 24216 25344
rect 24075 25313 24087 25316
rect 24029 25307 24087 25313
rect 24210 25304 24216 25316
rect 24268 25304 24274 25356
rect 15488 25248 16068 25276
rect 16485 25279 16543 25285
rect 14553 25239 14611 25245
rect 16485 25245 16497 25279
rect 16531 25276 16543 25279
rect 17310 25276 17316 25288
rect 16531 25248 17316 25276
rect 16531 25245 16543 25248
rect 16485 25239 16543 25245
rect 17310 25236 17316 25248
rect 17368 25236 17374 25288
rect 18785 25279 18843 25285
rect 18785 25276 18797 25279
rect 18156 25248 18797 25276
rect 10781 25211 10839 25217
rect 10781 25208 10793 25211
rect 7984 25180 8156 25208
rect 8588 25180 10793 25208
rect 7984 25168 7990 25180
rect 7377 25143 7435 25149
rect 7377 25140 7389 25143
rect 6512 25112 7389 25140
rect 6512 25100 6518 25112
rect 7377 25109 7389 25112
rect 7423 25109 7435 25143
rect 7377 25103 7435 25109
rect 7561 25143 7619 25149
rect 7561 25109 7573 25143
rect 7607 25140 7619 25143
rect 7650 25140 7656 25152
rect 7607 25112 7656 25140
rect 7607 25109 7619 25112
rect 7561 25103 7619 25109
rect 7650 25100 7656 25112
rect 7708 25100 7714 25152
rect 7834 25100 7840 25152
rect 7892 25140 7898 25152
rect 8588 25140 8616 25180
rect 10781 25177 10793 25180
rect 10827 25177 10839 25211
rect 10781 25171 10839 25177
rect 10965 25211 11023 25217
rect 10965 25177 10977 25211
rect 11011 25208 11023 25211
rect 18156 25208 18184 25248
rect 18785 25245 18797 25248
rect 18831 25245 18843 25279
rect 18966 25276 18972 25288
rect 18927 25248 18972 25276
rect 18785 25239 18843 25245
rect 11011 25180 18184 25208
rect 18800 25208 18828 25239
rect 18966 25236 18972 25248
rect 19024 25236 19030 25288
rect 19242 25236 19248 25288
rect 19300 25276 19306 25288
rect 21545 25279 21603 25285
rect 19300 25248 20944 25276
rect 19300 25236 19306 25248
rect 20441 25211 20499 25217
rect 20441 25208 20453 25211
rect 18800 25180 20453 25208
rect 11011 25177 11023 25180
rect 10965 25171 11023 25177
rect 20441 25177 20453 25180
rect 20487 25177 20499 25211
rect 20916 25208 20944 25248
rect 21545 25245 21557 25279
rect 21591 25276 21603 25279
rect 23198 25276 23204 25288
rect 21591 25248 23204 25276
rect 21591 25245 21603 25248
rect 21545 25239 21603 25245
rect 23198 25236 23204 25248
rect 23256 25236 23262 25288
rect 22465 25211 22523 25217
rect 22465 25208 22477 25211
rect 20916 25180 22477 25208
rect 20441 25171 20499 25177
rect 22465 25177 22477 25180
rect 22511 25177 22523 25211
rect 22465 25171 22523 25177
rect 7892 25112 8616 25140
rect 8665 25143 8723 25149
rect 7892 25100 7898 25112
rect 8665 25109 8677 25143
rect 8711 25140 8723 25143
rect 8754 25140 8760 25152
rect 8711 25112 8760 25140
rect 8711 25109 8723 25112
rect 8665 25103 8723 25109
rect 8754 25100 8760 25112
rect 8812 25100 8818 25152
rect 9585 25143 9643 25149
rect 9585 25109 9597 25143
rect 9631 25140 9643 25143
rect 9766 25140 9772 25152
rect 9631 25112 9772 25140
rect 9631 25109 9643 25112
rect 9585 25103 9643 25109
rect 9766 25100 9772 25112
rect 9824 25100 9830 25152
rect 11974 25140 11980 25152
rect 11935 25112 11980 25140
rect 11974 25100 11980 25112
rect 12032 25100 12038 25152
rect 12434 25100 12440 25152
rect 12492 25140 12498 25152
rect 12621 25143 12679 25149
rect 12492 25112 12537 25140
rect 12492 25100 12498 25112
rect 12621 25109 12633 25143
rect 12667 25140 12679 25143
rect 12986 25140 12992 25152
rect 12667 25112 12992 25140
rect 12667 25109 12679 25112
rect 12621 25103 12679 25109
rect 12986 25100 12992 25112
rect 13044 25100 13050 25152
rect 13170 25100 13176 25152
rect 13228 25140 13234 25152
rect 13633 25143 13691 25149
rect 13633 25140 13645 25143
rect 13228 25112 13645 25140
rect 13228 25100 13234 25112
rect 13633 25109 13645 25112
rect 13679 25109 13691 25143
rect 14826 25140 14832 25152
rect 14787 25112 14832 25140
rect 13633 25103 13691 25109
rect 14826 25100 14832 25112
rect 14884 25100 14890 25152
rect 15197 25143 15255 25149
rect 15197 25109 15209 25143
rect 15243 25140 15255 25143
rect 15286 25140 15292 25152
rect 15243 25112 15292 25140
rect 15243 25109 15255 25112
rect 15197 25103 15255 25109
rect 15286 25100 15292 25112
rect 15344 25100 15350 25152
rect 16666 25140 16672 25152
rect 16627 25112 16672 25140
rect 16666 25100 16672 25112
rect 16724 25100 16730 25152
rect 17310 25100 17316 25152
rect 17368 25140 17374 25152
rect 17589 25143 17647 25149
rect 17589 25140 17601 25143
rect 17368 25112 17601 25140
rect 17368 25100 17374 25112
rect 17589 25109 17601 25112
rect 17635 25109 17647 25143
rect 18138 25140 18144 25152
rect 18099 25112 18144 25140
rect 17589 25103 17647 25109
rect 18138 25100 18144 25112
rect 18196 25100 18202 25152
rect 18230 25100 18236 25152
rect 18288 25140 18294 25152
rect 18325 25143 18383 25149
rect 18325 25140 18337 25143
rect 18288 25112 18337 25140
rect 18288 25100 18294 25112
rect 18325 25109 18337 25112
rect 18371 25109 18383 25143
rect 18325 25103 18383 25109
rect 18782 25100 18788 25152
rect 18840 25140 18846 25152
rect 21545 25143 21603 25149
rect 21545 25140 21557 25143
rect 18840 25112 21557 25140
rect 18840 25100 18846 25112
rect 21545 25109 21557 25112
rect 21591 25109 21603 25143
rect 21726 25140 21732 25152
rect 21687 25112 21732 25140
rect 21545 25103 21603 25109
rect 21726 25100 21732 25112
rect 21784 25100 21790 25152
rect 24213 25143 24271 25149
rect 24213 25109 24225 25143
rect 24259 25140 24271 25143
rect 26050 25140 26056 25152
rect 24259 25112 26056 25140
rect 24259 25109 24271 25112
rect 24213 25103 24271 25109
rect 26050 25100 26056 25112
rect 26108 25100 26114 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 6730 24896 6736 24948
rect 6788 24936 6794 24948
rect 6788 24908 12940 24936
rect 6788 24896 6794 24908
rect 3418 24828 3424 24880
rect 3476 24868 3482 24880
rect 4525 24871 4583 24877
rect 4525 24868 4537 24871
rect 3476 24840 4537 24868
rect 3476 24828 3482 24840
rect 4525 24837 4537 24840
rect 4571 24837 4583 24871
rect 4525 24831 4583 24837
rect 4706 24828 4712 24880
rect 4764 24868 4770 24880
rect 4764 24840 5120 24868
rect 4764 24828 4770 24840
rect 5092 24809 5120 24840
rect 7926 24828 7932 24880
rect 7984 24868 7990 24880
rect 11054 24868 11060 24880
rect 7984 24840 8708 24868
rect 7984 24828 7990 24840
rect 8680 24809 8708 24840
rect 8772 24840 10916 24868
rect 11015 24840 11060 24868
rect 5077 24803 5135 24809
rect 5077 24769 5089 24803
rect 5123 24769 5135 24803
rect 5077 24763 5135 24769
rect 8665 24803 8723 24809
rect 8665 24769 8677 24803
rect 8711 24769 8723 24803
rect 8665 24763 8723 24769
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 1578 24732 1584 24744
rect 1443 24704 1584 24732
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 1578 24692 1584 24704
rect 1636 24732 1642 24744
rect 2317 24735 2375 24741
rect 2317 24732 2329 24735
rect 1636 24704 2329 24732
rect 1636 24692 1642 24704
rect 2317 24701 2329 24704
rect 2363 24701 2375 24735
rect 2317 24695 2375 24701
rect 2406 24692 2412 24744
rect 2464 24732 2470 24744
rect 2501 24735 2559 24741
rect 2501 24732 2513 24735
rect 2464 24704 2513 24732
rect 2464 24692 2470 24704
rect 2501 24701 2513 24704
rect 2547 24732 2559 24735
rect 3053 24735 3111 24741
rect 3053 24732 3065 24735
rect 2547 24704 3065 24732
rect 2547 24701 2559 24704
rect 2501 24695 2559 24701
rect 3053 24701 3065 24704
rect 3099 24701 3111 24735
rect 3053 24695 3111 24701
rect 4893 24735 4951 24741
rect 4893 24701 4905 24735
rect 4939 24732 4951 24735
rect 4982 24732 4988 24744
rect 4939 24704 4988 24732
rect 4939 24701 4951 24704
rect 4893 24695 4951 24701
rect 4982 24692 4988 24704
rect 5040 24692 5046 24744
rect 7466 24692 7472 24744
rect 7524 24732 7530 24744
rect 8772 24732 8800 24840
rect 10226 24800 10232 24812
rect 10187 24772 10232 24800
rect 10226 24760 10232 24772
rect 10284 24760 10290 24812
rect 10888 24800 10916 24840
rect 11054 24828 11060 24840
rect 11112 24828 11118 24880
rect 11514 24868 11520 24880
rect 11164 24840 11520 24868
rect 11164 24800 11192 24840
rect 11514 24828 11520 24840
rect 11572 24828 11578 24880
rect 10888 24772 11192 24800
rect 12250 24760 12256 24812
rect 12308 24800 12314 24812
rect 12308 24772 12848 24800
rect 12308 24760 12314 24772
rect 7524 24704 8800 24732
rect 7524 24692 7530 24704
rect 9490 24692 9496 24744
rect 9548 24732 9554 24744
rect 10137 24735 10195 24741
rect 10137 24732 10149 24735
rect 9548 24704 10149 24732
rect 9548 24692 9554 24704
rect 10137 24701 10149 24704
rect 10183 24701 10195 24735
rect 10137 24695 10195 24701
rect 11241 24735 11299 24741
rect 11241 24701 11253 24735
rect 11287 24732 11299 24735
rect 12342 24732 12348 24744
rect 11287 24704 12348 24732
rect 11287 24701 11299 24704
rect 11241 24695 11299 24701
rect 12342 24692 12348 24704
rect 12400 24692 12406 24744
rect 12820 24741 12848 24772
rect 12805 24735 12863 24741
rect 12805 24701 12817 24735
rect 12851 24701 12863 24735
rect 12912 24732 12940 24908
rect 13078 24896 13084 24948
rect 13136 24936 13142 24948
rect 13449 24939 13507 24945
rect 13449 24936 13461 24939
rect 13136 24908 13461 24936
rect 13136 24896 13142 24908
rect 13449 24905 13461 24908
rect 13495 24905 13507 24939
rect 13449 24899 13507 24905
rect 14090 24896 14096 24948
rect 14148 24936 14154 24948
rect 14148 24908 24992 24936
rect 14148 24896 14154 24908
rect 12986 24828 12992 24880
rect 13044 24868 13050 24880
rect 15654 24868 15660 24880
rect 13044 24840 15660 24868
rect 13044 24828 13050 24840
rect 15654 24828 15660 24840
rect 15712 24828 15718 24880
rect 15746 24828 15752 24880
rect 15804 24868 15810 24880
rect 18874 24868 18880 24880
rect 15804 24840 18880 24868
rect 15804 24828 15810 24840
rect 18874 24828 18880 24840
rect 18932 24828 18938 24880
rect 20622 24868 20628 24880
rect 20088 24840 20628 24868
rect 13081 24803 13139 24809
rect 13081 24769 13093 24803
rect 13127 24800 13139 24803
rect 13446 24800 13452 24812
rect 13127 24772 13452 24800
rect 13127 24769 13139 24772
rect 13081 24763 13139 24769
rect 13446 24760 13452 24772
rect 13504 24760 13510 24812
rect 13998 24760 14004 24812
rect 14056 24800 14062 24812
rect 14185 24803 14243 24809
rect 14185 24800 14197 24803
rect 14056 24772 14197 24800
rect 14056 24760 14062 24772
rect 14185 24769 14197 24772
rect 14231 24769 14243 24803
rect 14826 24800 14832 24812
rect 14787 24772 14832 24800
rect 14185 24763 14243 24769
rect 14826 24760 14832 24772
rect 14884 24760 14890 24812
rect 14921 24803 14979 24809
rect 14921 24769 14933 24803
rect 14967 24769 14979 24803
rect 14921 24763 14979 24769
rect 17037 24803 17095 24809
rect 17037 24769 17049 24803
rect 17083 24800 17095 24803
rect 17310 24800 17316 24812
rect 17083 24772 17316 24800
rect 17083 24769 17095 24772
rect 17037 24763 17095 24769
rect 14366 24732 14372 24744
rect 12912 24704 14372 24732
rect 12805 24695 12863 24701
rect 14366 24692 14372 24704
rect 14424 24692 14430 24744
rect 14458 24692 14464 24744
rect 14516 24732 14522 24744
rect 14936 24732 14964 24763
rect 17310 24760 17316 24772
rect 17368 24760 17374 24812
rect 17402 24760 17408 24812
rect 17460 24800 17466 24812
rect 18230 24800 18236 24812
rect 17460 24772 18236 24800
rect 17460 24760 17466 24772
rect 18230 24760 18236 24772
rect 18288 24760 18294 24812
rect 18598 24800 18604 24812
rect 18559 24772 18604 24800
rect 18598 24760 18604 24772
rect 18656 24800 18662 24812
rect 18966 24800 18972 24812
rect 18656 24772 18972 24800
rect 18656 24760 18662 24772
rect 18966 24760 18972 24772
rect 19024 24760 19030 24812
rect 20088 24809 20116 24840
rect 20622 24828 20628 24840
rect 20680 24868 20686 24880
rect 24762 24868 24768 24880
rect 20680 24840 24768 24868
rect 20680 24828 20686 24840
rect 24762 24828 24768 24840
rect 24820 24828 24826 24880
rect 19521 24803 19579 24809
rect 19521 24769 19533 24803
rect 19567 24800 19579 24803
rect 20073 24803 20131 24809
rect 20073 24800 20085 24803
rect 19567 24772 20085 24800
rect 19567 24769 19579 24772
rect 19521 24763 19579 24769
rect 20073 24769 20085 24772
rect 20119 24769 20131 24803
rect 20073 24763 20131 24769
rect 20257 24803 20315 24809
rect 20257 24769 20269 24803
rect 20303 24800 20315 24803
rect 20346 24800 20352 24812
rect 20303 24772 20352 24800
rect 20303 24769 20315 24772
rect 20257 24763 20315 24769
rect 20346 24760 20352 24772
rect 20404 24760 20410 24812
rect 20714 24800 20720 24812
rect 20675 24772 20720 24800
rect 20714 24760 20720 24772
rect 20772 24760 20778 24812
rect 24964 24809 24992 24908
rect 24949 24803 25007 24809
rect 24949 24769 24961 24803
rect 24995 24769 25007 24803
rect 24949 24763 25007 24769
rect 14516 24704 14964 24732
rect 14516 24692 14522 24704
rect 18138 24692 18144 24744
rect 18196 24732 18202 24744
rect 18417 24735 18475 24741
rect 18417 24732 18429 24735
rect 18196 24704 18429 24732
rect 18196 24692 18202 24704
rect 18417 24701 18429 24704
rect 18463 24732 18475 24735
rect 19978 24732 19984 24744
rect 18463 24704 19984 24732
rect 18463 24701 18475 24704
rect 18417 24695 18475 24701
rect 19978 24692 19984 24704
rect 20036 24692 20042 24744
rect 21637 24735 21695 24741
rect 21637 24701 21649 24735
rect 21683 24732 21695 24735
rect 21726 24732 21732 24744
rect 21683 24704 21732 24732
rect 21683 24701 21695 24704
rect 21637 24695 21695 24701
rect 21726 24692 21732 24704
rect 21784 24692 21790 24744
rect 23845 24735 23903 24741
rect 23845 24732 23857 24735
rect 23584 24704 23857 24732
rect 7101 24667 7159 24673
rect 3712 24636 5028 24664
rect 1394 24556 1400 24608
rect 1452 24596 1458 24608
rect 1581 24599 1639 24605
rect 1581 24596 1593 24599
rect 1452 24568 1593 24596
rect 1452 24556 1458 24568
rect 1581 24565 1593 24568
rect 1627 24565 1639 24599
rect 1581 24559 1639 24565
rect 2041 24599 2099 24605
rect 2041 24565 2053 24599
rect 2087 24596 2099 24599
rect 2130 24596 2136 24608
rect 2087 24568 2136 24596
rect 2087 24565 2099 24568
rect 2041 24559 2099 24565
rect 2130 24556 2136 24568
rect 2188 24556 2194 24608
rect 2406 24556 2412 24608
rect 2464 24596 2470 24608
rect 2685 24599 2743 24605
rect 2685 24596 2697 24599
rect 2464 24568 2697 24596
rect 2464 24556 2470 24568
rect 2685 24565 2697 24568
rect 2731 24565 2743 24599
rect 2685 24559 2743 24565
rect 3050 24556 3056 24608
rect 3108 24596 3114 24608
rect 3712 24605 3740 24636
rect 3697 24599 3755 24605
rect 3697 24596 3709 24599
rect 3108 24568 3709 24596
rect 3108 24556 3114 24568
rect 3697 24565 3709 24568
rect 3743 24565 3755 24599
rect 3697 24559 3755 24565
rect 3786 24556 3792 24608
rect 3844 24596 3850 24608
rect 4062 24596 4068 24608
rect 3844 24568 4068 24596
rect 3844 24556 3850 24568
rect 4062 24556 4068 24568
rect 4120 24556 4126 24608
rect 5000 24605 5028 24636
rect 7101 24633 7113 24667
rect 7147 24664 7159 24667
rect 9125 24667 9183 24673
rect 9125 24664 9137 24667
rect 7147 24636 9137 24664
rect 7147 24633 7159 24636
rect 7101 24627 7159 24633
rect 9125 24633 9137 24636
rect 9171 24664 9183 24667
rect 10045 24667 10103 24673
rect 10045 24664 10057 24667
rect 9171 24636 10057 24664
rect 9171 24633 9183 24636
rect 9125 24627 9183 24633
rect 10045 24633 10057 24636
rect 10091 24633 10103 24667
rect 10045 24627 10103 24633
rect 11885 24667 11943 24673
rect 11885 24633 11897 24667
rect 11931 24664 11943 24667
rect 12897 24667 12955 24673
rect 12897 24664 12909 24667
rect 11931 24636 12909 24664
rect 11931 24633 11943 24636
rect 11885 24627 11943 24633
rect 12897 24633 12909 24636
rect 12943 24664 12955 24667
rect 14737 24667 14795 24673
rect 12943 24636 14688 24664
rect 12943 24633 12955 24636
rect 12897 24627 12955 24633
rect 4985 24599 5043 24605
rect 4985 24565 4997 24599
rect 5031 24565 5043 24599
rect 4985 24559 5043 24565
rect 5994 24556 6000 24608
rect 6052 24596 6058 24608
rect 6546 24596 6552 24608
rect 6052 24568 6552 24596
rect 6052 24556 6058 24568
rect 6546 24556 6552 24568
rect 6604 24556 6610 24608
rect 7653 24599 7711 24605
rect 7653 24565 7665 24599
rect 7699 24596 7711 24599
rect 7926 24596 7932 24608
rect 7699 24568 7932 24596
rect 7699 24565 7711 24568
rect 7653 24559 7711 24565
rect 7926 24556 7932 24568
rect 7984 24556 7990 24608
rect 8110 24596 8116 24608
rect 8071 24568 8116 24596
rect 8110 24556 8116 24568
rect 8168 24556 8174 24608
rect 8202 24556 8208 24608
rect 8260 24596 8266 24608
rect 8481 24599 8539 24605
rect 8481 24596 8493 24599
rect 8260 24568 8493 24596
rect 8260 24556 8266 24568
rect 8481 24565 8493 24568
rect 8527 24565 8539 24599
rect 8481 24559 8539 24565
rect 8573 24599 8631 24605
rect 8573 24565 8585 24599
rect 8619 24596 8631 24599
rect 8754 24596 8760 24608
rect 8619 24568 8760 24596
rect 8619 24565 8631 24568
rect 8573 24559 8631 24565
rect 8754 24556 8760 24568
rect 8812 24556 8818 24608
rect 9490 24596 9496 24608
rect 9451 24568 9496 24596
rect 9490 24556 9496 24568
rect 9548 24556 9554 24608
rect 9674 24596 9680 24608
rect 9635 24568 9680 24596
rect 9674 24556 9680 24568
rect 9732 24556 9738 24608
rect 11422 24596 11428 24608
rect 11383 24568 11428 24596
rect 11422 24556 11428 24568
rect 11480 24556 11486 24608
rect 12250 24596 12256 24608
rect 12211 24568 12256 24596
rect 12250 24556 12256 24568
rect 12308 24556 12314 24608
rect 12437 24599 12495 24605
rect 12437 24565 12449 24599
rect 12483 24596 12495 24599
rect 12710 24596 12716 24608
rect 12483 24568 12716 24596
rect 12483 24565 12495 24568
rect 12437 24559 12495 24565
rect 12710 24556 12716 24568
rect 12768 24556 12774 24608
rect 13446 24556 13452 24608
rect 13504 24596 13510 24608
rect 13817 24599 13875 24605
rect 13817 24596 13829 24599
rect 13504 24568 13829 24596
rect 13504 24556 13510 24568
rect 13817 24565 13829 24568
rect 13863 24565 13875 24599
rect 13817 24559 13875 24565
rect 14369 24599 14427 24605
rect 14369 24565 14381 24599
rect 14415 24596 14427 24599
rect 14550 24596 14556 24608
rect 14415 24568 14556 24596
rect 14415 24565 14427 24568
rect 14369 24559 14427 24565
rect 14550 24556 14556 24568
rect 14608 24556 14614 24608
rect 14660 24596 14688 24636
rect 14737 24633 14749 24667
rect 14783 24664 14795 24667
rect 14918 24664 14924 24676
rect 14783 24636 14924 24664
rect 14783 24633 14795 24636
rect 14737 24627 14795 24633
rect 14918 24624 14924 24636
rect 14976 24624 14982 24676
rect 16298 24664 16304 24676
rect 16259 24636 16304 24664
rect 16298 24624 16304 24636
rect 16356 24664 16362 24676
rect 16853 24667 16911 24673
rect 16853 24664 16865 24667
rect 16356 24636 16865 24664
rect 16356 24624 16362 24636
rect 16853 24633 16865 24636
rect 16899 24633 16911 24667
rect 16853 24627 16911 24633
rect 17586 24624 17592 24676
rect 17644 24664 17650 24676
rect 17865 24667 17923 24673
rect 17865 24664 17877 24667
rect 17644 24636 17877 24664
rect 17644 24624 17650 24636
rect 17865 24633 17877 24636
rect 17911 24664 17923 24667
rect 18506 24664 18512 24676
rect 17911 24636 18512 24664
rect 17911 24633 17923 24636
rect 17865 24627 17923 24633
rect 18506 24624 18512 24636
rect 18564 24624 18570 24676
rect 18690 24624 18696 24676
rect 18748 24664 18754 24676
rect 19061 24667 19119 24673
rect 19061 24664 19073 24667
rect 18748 24636 19073 24664
rect 18748 24624 18754 24636
rect 19061 24633 19073 24636
rect 19107 24633 19119 24667
rect 20530 24664 20536 24676
rect 19061 24627 19119 24633
rect 19628 24636 20536 24664
rect 15378 24596 15384 24608
rect 14660 24568 15384 24596
rect 15378 24556 15384 24568
rect 15436 24556 15442 24608
rect 15657 24599 15715 24605
rect 15657 24565 15669 24599
rect 15703 24596 15715 24599
rect 15930 24596 15936 24608
rect 15703 24568 15936 24596
rect 15703 24565 15715 24568
rect 15657 24559 15715 24565
rect 15930 24556 15936 24568
rect 15988 24556 15994 24608
rect 16390 24596 16396 24608
rect 16351 24568 16396 24596
rect 16390 24556 16396 24568
rect 16448 24556 16454 24608
rect 16482 24556 16488 24608
rect 16540 24596 16546 24608
rect 16761 24599 16819 24605
rect 16761 24596 16773 24599
rect 16540 24568 16773 24596
rect 16540 24556 16546 24568
rect 16761 24565 16773 24568
rect 16807 24565 16819 24599
rect 17494 24596 17500 24608
rect 17455 24568 17500 24596
rect 16761 24559 16819 24565
rect 17494 24556 17500 24568
rect 17552 24556 17558 24608
rect 17954 24556 17960 24608
rect 18012 24596 18018 24608
rect 19628 24605 19656 24636
rect 20530 24624 20536 24636
rect 20588 24624 20594 24676
rect 23584 24608 23612 24704
rect 23845 24701 23857 24704
rect 23891 24701 23903 24735
rect 23845 24695 23903 24701
rect 18049 24599 18107 24605
rect 18049 24596 18061 24599
rect 18012 24568 18061 24596
rect 18012 24556 18018 24568
rect 18049 24565 18061 24568
rect 18095 24565 18107 24599
rect 18049 24559 18107 24565
rect 19613 24599 19671 24605
rect 19613 24565 19625 24599
rect 19659 24565 19671 24599
rect 19613 24559 19671 24565
rect 21174 24556 21180 24608
rect 21232 24596 21238 24608
rect 21269 24599 21327 24605
rect 21269 24596 21281 24599
rect 21232 24568 21281 24596
rect 21232 24556 21238 24568
rect 21269 24565 21281 24568
rect 21315 24596 21327 24599
rect 21634 24596 21640 24608
rect 21315 24568 21640 24596
rect 21315 24565 21327 24568
rect 21269 24559 21327 24565
rect 21634 24556 21640 24568
rect 21692 24556 21698 24608
rect 21818 24596 21824 24608
rect 21779 24568 21824 24596
rect 21818 24556 21824 24568
rect 21876 24556 21882 24608
rect 22370 24596 22376 24608
rect 22331 24568 22376 24596
rect 22370 24556 22376 24568
rect 22428 24556 22434 24608
rect 23477 24599 23535 24605
rect 23477 24565 23489 24599
rect 23523 24596 23535 24599
rect 23566 24596 23572 24608
rect 23523 24568 23572 24596
rect 23523 24565 23535 24568
rect 23477 24559 23535 24565
rect 23566 24556 23572 24568
rect 23624 24556 23630 24608
rect 24026 24596 24032 24608
rect 23987 24568 24032 24596
rect 24026 24556 24032 24568
rect 24084 24556 24090 24608
rect 24394 24596 24400 24608
rect 24355 24568 24400 24596
rect 24394 24556 24400 24568
rect 24452 24556 24458 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 4801 24395 4859 24401
rect 4801 24361 4813 24395
rect 4847 24392 4859 24395
rect 4982 24392 4988 24404
rect 4847 24364 4988 24392
rect 4847 24361 4859 24364
rect 4801 24355 4859 24361
rect 4982 24352 4988 24364
rect 5040 24352 5046 24404
rect 5169 24395 5227 24401
rect 5169 24361 5181 24395
rect 5215 24392 5227 24395
rect 5258 24392 5264 24404
rect 5215 24364 5264 24392
rect 5215 24361 5227 24364
rect 5169 24355 5227 24361
rect 5258 24352 5264 24364
rect 5316 24352 5322 24404
rect 14826 24352 14832 24404
rect 14884 24392 14890 24404
rect 15289 24395 15347 24401
rect 15289 24392 15301 24395
rect 14884 24364 15301 24392
rect 14884 24352 14890 24364
rect 15289 24361 15301 24364
rect 15335 24361 15347 24395
rect 15289 24355 15347 24361
rect 15657 24395 15715 24401
rect 15657 24361 15669 24395
rect 15703 24392 15715 24395
rect 15746 24392 15752 24404
rect 15703 24364 15752 24392
rect 15703 24361 15715 24364
rect 15657 24355 15715 24361
rect 15746 24352 15752 24364
rect 15804 24352 15810 24404
rect 16482 24392 16488 24404
rect 16443 24364 16488 24392
rect 16482 24352 16488 24364
rect 16540 24352 16546 24404
rect 18782 24352 18788 24404
rect 18840 24392 18846 24404
rect 19153 24395 19211 24401
rect 19153 24392 19165 24395
rect 18840 24364 19165 24392
rect 18840 24352 18846 24364
rect 19153 24361 19165 24364
rect 19199 24361 19211 24395
rect 20622 24392 20628 24404
rect 20583 24364 20628 24392
rect 19153 24355 19211 24361
rect 20622 24352 20628 24364
rect 20680 24352 20686 24404
rect 22649 24395 22707 24401
rect 22649 24361 22661 24395
rect 22695 24392 22707 24395
rect 24118 24392 24124 24404
rect 22695 24364 24124 24392
rect 22695 24361 22707 24364
rect 22649 24355 22707 24361
rect 24118 24352 24124 24364
rect 24176 24352 24182 24404
rect 24670 24392 24676 24404
rect 24631 24364 24676 24392
rect 24670 24352 24676 24364
rect 24728 24352 24734 24404
rect 1118 24284 1124 24336
rect 1176 24324 1182 24336
rect 6178 24324 6184 24336
rect 1176 24296 5304 24324
rect 6139 24296 6184 24324
rect 1176 24284 1182 24296
rect 1854 24216 1860 24268
rect 1912 24256 1918 24268
rect 2041 24259 2099 24265
rect 2041 24256 2053 24259
rect 1912 24228 2053 24256
rect 1912 24216 1918 24228
rect 2041 24225 2053 24228
rect 2087 24256 2099 24259
rect 2222 24256 2228 24268
rect 2087 24228 2228 24256
rect 2087 24225 2099 24228
rect 2041 24219 2099 24225
rect 2222 24216 2228 24228
rect 2280 24216 2286 24268
rect 5276 24265 5304 24296
rect 6178 24284 6184 24296
rect 6236 24284 6242 24336
rect 7098 24284 7104 24336
rect 7156 24324 7162 24336
rect 9398 24324 9404 24336
rect 7156 24296 9404 24324
rect 7156 24284 7162 24296
rect 9398 24284 9404 24296
rect 9456 24284 9462 24336
rect 14182 24284 14188 24336
rect 14240 24324 14246 24336
rect 15013 24327 15071 24333
rect 15013 24324 15025 24327
rect 14240 24296 15025 24324
rect 14240 24284 14246 24296
rect 15013 24293 15025 24296
rect 15059 24324 15071 24327
rect 15378 24324 15384 24336
rect 15059 24296 15384 24324
rect 15059 24293 15071 24296
rect 15013 24287 15071 24293
rect 15378 24284 15384 24296
rect 15436 24284 15442 24336
rect 20990 24324 20996 24336
rect 15764 24296 20996 24324
rect 5261 24259 5319 24265
rect 5261 24225 5273 24259
rect 5307 24256 5319 24259
rect 5534 24256 5540 24268
rect 5307 24228 5540 24256
rect 5307 24225 5319 24228
rect 5261 24219 5319 24225
rect 5534 24216 5540 24228
rect 5592 24216 5598 24268
rect 6908 24259 6966 24265
rect 6908 24225 6920 24259
rect 6954 24256 6966 24259
rect 7190 24256 7196 24268
rect 6954 24228 7196 24256
rect 6954 24225 6966 24228
rect 6908 24219 6966 24225
rect 7190 24216 7196 24228
rect 7248 24216 7254 24268
rect 10134 24216 10140 24268
rect 10192 24256 10198 24268
rect 10669 24259 10727 24265
rect 10669 24256 10681 24259
rect 10192 24228 10681 24256
rect 10192 24216 10198 24228
rect 10669 24225 10681 24228
rect 10715 24225 10727 24259
rect 10669 24219 10727 24225
rect 12986 24216 12992 24268
rect 13044 24256 13050 24268
rect 13265 24259 13323 24265
rect 13265 24256 13277 24259
rect 13044 24228 13277 24256
rect 13044 24216 13050 24228
rect 13265 24225 13277 24228
rect 13311 24225 13323 24259
rect 13265 24219 13323 24225
rect 1946 24148 1952 24200
rect 2004 24188 2010 24200
rect 2130 24188 2136 24200
rect 2004 24160 2136 24188
rect 2004 24148 2010 24160
rect 2130 24148 2136 24160
rect 2188 24148 2194 24200
rect 2317 24191 2375 24197
rect 2317 24157 2329 24191
rect 2363 24188 2375 24191
rect 2958 24188 2964 24200
rect 2363 24160 2964 24188
rect 2363 24157 2375 24160
rect 2317 24151 2375 24157
rect 2958 24148 2964 24160
rect 3016 24148 3022 24200
rect 4709 24191 4767 24197
rect 4709 24157 4721 24191
rect 4755 24188 4767 24191
rect 5074 24188 5080 24200
rect 4755 24160 5080 24188
rect 4755 24157 4767 24160
rect 4709 24151 4767 24157
rect 5074 24148 5080 24160
rect 5132 24188 5138 24200
rect 5445 24191 5503 24197
rect 5445 24188 5457 24191
rect 5132 24160 5457 24188
rect 5132 24148 5138 24160
rect 5445 24157 5457 24160
rect 5491 24188 5503 24191
rect 6638 24188 6644 24200
rect 5491 24160 5948 24188
rect 6599 24160 6644 24188
rect 5491 24157 5503 24160
rect 5445 24151 5503 24157
rect 3329 24123 3387 24129
rect 3329 24089 3341 24123
rect 3375 24120 3387 24123
rect 3878 24120 3884 24132
rect 3375 24092 3884 24120
rect 3375 24089 3387 24092
rect 3329 24083 3387 24089
rect 3878 24080 3884 24092
rect 3936 24080 3942 24132
rect 1673 24055 1731 24061
rect 1673 24021 1685 24055
rect 1719 24052 1731 24055
rect 2222 24052 2228 24064
rect 1719 24024 2228 24052
rect 1719 24021 1731 24024
rect 1673 24015 1731 24021
rect 2222 24012 2228 24024
rect 2280 24012 2286 24064
rect 2498 24012 2504 24064
rect 2556 24052 2562 24064
rect 2777 24055 2835 24061
rect 2777 24052 2789 24055
rect 2556 24024 2789 24052
rect 2556 24012 2562 24024
rect 2777 24021 2789 24024
rect 2823 24021 2835 24055
rect 2777 24015 2835 24021
rect 3697 24055 3755 24061
rect 3697 24021 3709 24055
rect 3743 24052 3755 24055
rect 4062 24052 4068 24064
rect 3743 24024 4068 24052
rect 3743 24021 3755 24024
rect 3697 24015 3755 24021
rect 4062 24012 4068 24024
rect 4120 24012 4126 24064
rect 4338 24052 4344 24064
rect 4299 24024 4344 24052
rect 4338 24012 4344 24024
rect 4396 24012 4402 24064
rect 5920 24061 5948 24160
rect 6638 24148 6644 24160
rect 6696 24148 6702 24200
rect 10410 24188 10416 24200
rect 10371 24160 10416 24188
rect 10410 24148 10416 24160
rect 10468 24148 10474 24200
rect 11422 24148 11428 24200
rect 11480 24188 11486 24200
rect 12158 24188 12164 24200
rect 11480 24160 12164 24188
rect 11480 24148 11486 24160
rect 12158 24148 12164 24160
rect 12216 24188 12222 24200
rect 13354 24188 13360 24200
rect 12216 24160 13360 24188
rect 12216 24148 12222 24160
rect 13354 24148 13360 24160
rect 13412 24148 13418 24200
rect 13446 24148 13452 24200
rect 13504 24188 13510 24200
rect 13504 24160 13549 24188
rect 13504 24148 13510 24160
rect 14090 24148 14096 24200
rect 14148 24188 14154 24200
rect 15102 24188 15108 24200
rect 14148 24160 15108 24188
rect 14148 24148 14154 24160
rect 15102 24148 15108 24160
rect 15160 24148 15166 24200
rect 15286 24148 15292 24200
rect 15344 24188 15350 24200
rect 15764 24197 15792 24296
rect 20990 24284 20996 24296
rect 21048 24284 21054 24336
rect 16666 24216 16672 24268
rect 16724 24256 16730 24268
rect 17497 24259 17555 24265
rect 17497 24256 17509 24259
rect 16724 24228 17509 24256
rect 16724 24216 16730 24228
rect 17497 24225 17509 24228
rect 17543 24256 17555 24259
rect 17678 24256 17684 24268
rect 17543 24228 17684 24256
rect 17543 24225 17555 24228
rect 17497 24219 17555 24225
rect 17678 24216 17684 24228
rect 17736 24216 17742 24268
rect 19061 24259 19119 24265
rect 19061 24225 19073 24259
rect 19107 24256 19119 24259
rect 20438 24256 20444 24268
rect 19107 24228 20444 24256
rect 19107 24225 19119 24228
rect 19061 24219 19119 24225
rect 20438 24216 20444 24228
rect 20496 24216 20502 24268
rect 21266 24256 21272 24268
rect 21227 24228 21272 24256
rect 21266 24216 21272 24228
rect 21324 24216 21330 24268
rect 22465 24259 22523 24265
rect 22465 24225 22477 24259
rect 22511 24256 22523 24259
rect 22646 24256 22652 24268
rect 22511 24228 22652 24256
rect 22511 24225 22523 24228
rect 22465 24219 22523 24225
rect 22646 24216 22652 24228
rect 22704 24216 22710 24268
rect 24118 24216 24124 24268
rect 24176 24256 24182 24268
rect 24489 24259 24547 24265
rect 24489 24256 24501 24259
rect 24176 24228 24501 24256
rect 24176 24216 24182 24228
rect 24489 24225 24501 24228
rect 24535 24225 24547 24259
rect 24489 24219 24547 24225
rect 15749 24191 15807 24197
rect 15749 24188 15761 24191
rect 15344 24160 15761 24188
rect 15344 24148 15350 24160
rect 15749 24157 15761 24160
rect 15795 24157 15807 24191
rect 15749 24151 15807 24157
rect 15841 24191 15899 24197
rect 15841 24157 15853 24191
rect 15887 24157 15899 24191
rect 15841 24151 15899 24157
rect 16853 24191 16911 24197
rect 16853 24157 16865 24191
rect 16899 24188 16911 24191
rect 16942 24188 16948 24200
rect 16899 24160 16948 24188
rect 16899 24157 16911 24160
rect 16853 24151 16911 24157
rect 6362 24080 6368 24132
rect 6420 24120 6426 24132
rect 6546 24120 6552 24132
rect 6420 24092 6552 24120
rect 6420 24080 6426 24092
rect 6546 24080 6552 24092
rect 6604 24080 6610 24132
rect 8202 24080 8208 24132
rect 8260 24120 8266 24132
rect 8941 24123 8999 24129
rect 8941 24120 8953 24123
rect 8260 24092 8953 24120
rect 8260 24080 8266 24092
rect 8941 24089 8953 24092
rect 8987 24089 8999 24123
rect 8941 24083 8999 24089
rect 13998 24080 14004 24132
rect 14056 24120 14062 24132
rect 14826 24120 14832 24132
rect 14056 24092 14832 24120
rect 14056 24080 14062 24092
rect 14826 24080 14832 24092
rect 14884 24120 14890 24132
rect 15856 24120 15884 24151
rect 16942 24148 16948 24160
rect 17000 24148 17006 24200
rect 17402 24148 17408 24200
rect 17460 24188 17466 24200
rect 17589 24191 17647 24197
rect 17589 24188 17601 24191
rect 17460 24160 17601 24188
rect 17460 24148 17466 24160
rect 17589 24157 17601 24160
rect 17635 24157 17647 24191
rect 17589 24151 17647 24157
rect 17773 24191 17831 24197
rect 17773 24157 17785 24191
rect 17819 24188 17831 24191
rect 17862 24188 17868 24200
rect 17819 24160 17868 24188
rect 17819 24157 17831 24160
rect 17773 24151 17831 24157
rect 17862 24148 17868 24160
rect 17920 24148 17926 24200
rect 18233 24191 18291 24197
rect 18233 24157 18245 24191
rect 18279 24188 18291 24191
rect 18598 24188 18604 24200
rect 18279 24160 18604 24188
rect 18279 24157 18291 24160
rect 18233 24151 18291 24157
rect 18598 24148 18604 24160
rect 18656 24188 18662 24200
rect 19245 24191 19303 24197
rect 19245 24188 19257 24191
rect 18656 24160 19257 24188
rect 18656 24148 18662 24160
rect 19245 24157 19257 24160
rect 19291 24188 19303 24191
rect 20714 24188 20720 24200
rect 19291 24160 20720 24188
rect 19291 24157 19303 24160
rect 19245 24151 19303 24157
rect 20714 24148 20720 24160
rect 20772 24148 20778 24200
rect 21358 24188 21364 24200
rect 21319 24160 21364 24188
rect 21358 24148 21364 24160
rect 21416 24148 21422 24200
rect 21453 24191 21511 24197
rect 21453 24157 21465 24191
rect 21499 24157 21511 24191
rect 21453 24151 21511 24157
rect 14884 24092 15884 24120
rect 14884 24080 14890 24092
rect 16666 24080 16672 24132
rect 16724 24120 16730 24132
rect 18414 24120 18420 24132
rect 16724 24092 18420 24120
rect 16724 24080 16730 24092
rect 18414 24080 18420 24092
rect 18472 24080 18478 24132
rect 21468 24120 21496 24151
rect 20364 24092 21496 24120
rect 20364 24064 20392 24092
rect 5905 24055 5963 24061
rect 5905 24021 5917 24055
rect 5951 24052 5963 24055
rect 6086 24052 6092 24064
rect 5951 24024 6092 24052
rect 5951 24021 5963 24024
rect 5905 24015 5963 24021
rect 6086 24012 6092 24024
rect 6144 24052 6150 24064
rect 7558 24052 7564 24064
rect 6144 24024 7564 24052
rect 6144 24012 6150 24024
rect 7558 24012 7564 24024
rect 7616 24052 7622 24064
rect 8021 24055 8079 24061
rect 8021 24052 8033 24055
rect 7616 24024 8033 24052
rect 7616 24012 7622 24024
rect 8021 24021 8033 24024
rect 8067 24021 8079 24055
rect 8662 24052 8668 24064
rect 8623 24024 8668 24052
rect 8021 24015 8079 24021
rect 8662 24012 8668 24024
rect 8720 24012 8726 24064
rect 9953 24055 10011 24061
rect 9953 24021 9965 24055
rect 9999 24052 10011 24055
rect 10134 24052 10140 24064
rect 9999 24024 10140 24052
rect 9999 24021 10011 24024
rect 9953 24015 10011 24021
rect 10134 24012 10140 24024
rect 10192 24012 10198 24064
rect 10318 24052 10324 24064
rect 10279 24024 10324 24052
rect 10318 24012 10324 24024
rect 10376 24012 10382 24064
rect 11790 24052 11796 24064
rect 11751 24024 11796 24052
rect 11790 24012 11796 24024
rect 11848 24012 11854 24064
rect 12066 24012 12072 24064
rect 12124 24052 12130 24064
rect 12621 24055 12679 24061
rect 12621 24052 12633 24055
rect 12124 24024 12633 24052
rect 12124 24012 12130 24024
rect 12621 24021 12633 24024
rect 12667 24021 12679 24055
rect 12894 24052 12900 24064
rect 12855 24024 12900 24052
rect 12621 24015 12679 24021
rect 12894 24012 12900 24024
rect 12952 24012 12958 24064
rect 13722 24012 13728 24064
rect 13780 24052 13786 24064
rect 13909 24055 13967 24061
rect 13909 24052 13921 24055
rect 13780 24024 13921 24052
rect 13780 24012 13786 24024
rect 13909 24021 13921 24024
rect 13955 24021 13967 24055
rect 14458 24052 14464 24064
rect 14419 24024 14464 24052
rect 13909 24015 13967 24021
rect 14458 24012 14464 24024
rect 14516 24012 14522 24064
rect 17129 24055 17187 24061
rect 17129 24021 17141 24055
rect 17175 24052 17187 24055
rect 18046 24052 18052 24064
rect 17175 24024 18052 24052
rect 17175 24021 17187 24024
rect 17129 24015 17187 24021
rect 18046 24012 18052 24024
rect 18104 24012 18110 24064
rect 18693 24055 18751 24061
rect 18693 24021 18705 24055
rect 18739 24052 18751 24055
rect 19242 24052 19248 24064
rect 18739 24024 19248 24052
rect 18739 24021 18751 24024
rect 18693 24015 18751 24021
rect 19242 24012 19248 24024
rect 19300 24012 19306 24064
rect 19797 24055 19855 24061
rect 19797 24021 19809 24055
rect 19843 24052 19855 24055
rect 20257 24055 20315 24061
rect 20257 24052 20269 24055
rect 19843 24024 20269 24052
rect 19843 24021 19855 24024
rect 19797 24015 19855 24021
rect 20257 24021 20269 24024
rect 20303 24052 20315 24055
rect 20346 24052 20352 24064
rect 20303 24024 20352 24052
rect 20303 24021 20315 24024
rect 20257 24015 20315 24021
rect 20346 24012 20352 24024
rect 20404 24012 20410 24064
rect 20901 24055 20959 24061
rect 20901 24021 20913 24055
rect 20947 24052 20959 24055
rect 21542 24052 21548 24064
rect 20947 24024 21548 24052
rect 20947 24021 20959 24024
rect 20901 24015 20959 24021
rect 21542 24012 21548 24024
rect 21600 24012 21606 24064
rect 21818 24012 21824 24064
rect 21876 24052 21882 24064
rect 21913 24055 21971 24061
rect 21913 24052 21925 24055
rect 21876 24024 21925 24052
rect 21876 24012 21882 24024
rect 21913 24021 21925 24024
rect 21959 24021 21971 24055
rect 21913 24015 21971 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 3142 23808 3148 23860
rect 3200 23848 3206 23860
rect 3605 23851 3663 23857
rect 3605 23848 3617 23851
rect 3200 23820 3617 23848
rect 3200 23808 3206 23820
rect 3605 23817 3617 23820
rect 3651 23817 3663 23851
rect 3605 23811 3663 23817
rect 5534 23808 5540 23860
rect 5592 23848 5598 23860
rect 6181 23851 6239 23857
rect 6181 23848 6193 23851
rect 5592 23820 6193 23848
rect 5592 23808 5598 23820
rect 6181 23817 6193 23820
rect 6227 23817 6239 23851
rect 7466 23848 7472 23860
rect 7427 23820 7472 23848
rect 6181 23811 6239 23817
rect 7466 23808 7472 23820
rect 7524 23808 7530 23860
rect 12158 23848 12164 23860
rect 12119 23820 12164 23848
rect 12158 23808 12164 23820
rect 12216 23808 12222 23860
rect 14734 23848 14740 23860
rect 12452 23820 14596 23848
rect 14647 23820 14740 23848
rect 5169 23783 5227 23789
rect 5169 23780 5181 23783
rect 2240 23752 2820 23780
rect 2038 23672 2044 23724
rect 2096 23712 2102 23724
rect 2240 23721 2268 23752
rect 2133 23715 2191 23721
rect 2133 23712 2145 23715
rect 2096 23684 2145 23712
rect 2096 23672 2102 23684
rect 2133 23681 2145 23684
rect 2179 23681 2191 23715
rect 2133 23675 2191 23681
rect 2225 23715 2283 23721
rect 2225 23681 2237 23715
rect 2271 23681 2283 23715
rect 2225 23675 2283 23681
rect 2041 23579 2099 23585
rect 2041 23545 2053 23579
rect 2087 23576 2099 23579
rect 2314 23576 2320 23588
rect 2087 23548 2320 23576
rect 2087 23545 2099 23548
rect 2041 23539 2099 23545
rect 2314 23536 2320 23548
rect 2372 23536 2378 23588
rect 2792 23585 2820 23752
rect 4080 23752 5181 23780
rect 4080 23724 4108 23752
rect 5169 23749 5181 23752
rect 5215 23749 5227 23783
rect 5169 23743 5227 23749
rect 10962 23740 10968 23792
rect 11020 23780 11026 23792
rect 11020 23752 11468 23780
rect 11020 23740 11026 23752
rect 4062 23712 4068 23724
rect 4023 23684 4068 23712
rect 4062 23672 4068 23684
rect 4120 23672 4126 23724
rect 4249 23715 4307 23721
rect 4249 23681 4261 23715
rect 4295 23712 4307 23715
rect 4522 23712 4528 23724
rect 4295 23684 4528 23712
rect 4295 23681 4307 23684
rect 4249 23675 4307 23681
rect 3878 23604 3884 23656
rect 3936 23644 3942 23656
rect 3973 23647 4031 23653
rect 3973 23644 3985 23647
rect 3936 23616 3985 23644
rect 3936 23604 3942 23616
rect 3973 23613 3985 23616
rect 4019 23613 4031 23647
rect 4264 23644 4292 23675
rect 4522 23672 4528 23684
rect 4580 23712 4586 23724
rect 4706 23712 4712 23724
rect 4580 23684 4712 23712
rect 4580 23672 4586 23684
rect 4706 23672 4712 23684
rect 4764 23672 4770 23724
rect 5442 23672 5448 23724
rect 5500 23712 5506 23724
rect 5629 23715 5687 23721
rect 5629 23712 5641 23715
rect 5500 23684 5641 23712
rect 5500 23672 5506 23684
rect 5629 23681 5641 23684
rect 5675 23681 5687 23715
rect 5629 23675 5687 23681
rect 5813 23715 5871 23721
rect 5813 23681 5825 23715
rect 5859 23712 5871 23715
rect 6086 23712 6092 23724
rect 5859 23684 6092 23712
rect 5859 23681 5871 23684
rect 5813 23675 5871 23681
rect 6086 23672 6092 23684
rect 6144 23672 6150 23724
rect 10318 23672 10324 23724
rect 10376 23712 10382 23724
rect 11440 23721 11468 23752
rect 11698 23740 11704 23792
rect 11756 23780 11762 23792
rect 12452 23780 12480 23820
rect 11756 23752 12480 23780
rect 14568 23780 14596 23820
rect 14734 23808 14740 23820
rect 14792 23848 14798 23860
rect 15838 23848 15844 23860
rect 14792 23820 15844 23848
rect 14792 23808 14798 23820
rect 15838 23808 15844 23820
rect 15896 23808 15902 23860
rect 16577 23851 16635 23857
rect 16577 23817 16589 23851
rect 16623 23848 16635 23851
rect 16758 23848 16764 23860
rect 16623 23820 16764 23848
rect 16623 23817 16635 23820
rect 16577 23811 16635 23817
rect 16758 23808 16764 23820
rect 16816 23848 16822 23860
rect 17221 23851 17279 23857
rect 17221 23848 17233 23851
rect 16816 23820 17233 23848
rect 16816 23808 16822 23820
rect 17221 23817 17233 23820
rect 17267 23848 17279 23851
rect 17310 23848 17316 23860
rect 17267 23820 17316 23848
rect 17267 23817 17279 23820
rect 17221 23811 17279 23817
rect 17310 23808 17316 23820
rect 17368 23808 17374 23860
rect 20349 23851 20407 23857
rect 20349 23848 20361 23851
rect 17788 23820 20361 23848
rect 15013 23783 15071 23789
rect 15013 23780 15025 23783
rect 14568 23752 15025 23780
rect 11756 23740 11762 23752
rect 15013 23749 15025 23752
rect 15059 23780 15071 23783
rect 15194 23780 15200 23792
rect 15059 23752 15200 23780
rect 15059 23749 15071 23752
rect 15013 23743 15071 23749
rect 15194 23740 15200 23752
rect 15252 23740 15258 23792
rect 11241 23715 11299 23721
rect 11241 23712 11253 23715
rect 10376 23684 11253 23712
rect 10376 23672 10382 23684
rect 11241 23681 11253 23684
rect 11287 23681 11299 23715
rect 11241 23675 11299 23681
rect 11425 23715 11483 23721
rect 11425 23681 11437 23715
rect 11471 23712 11483 23715
rect 11790 23712 11796 23724
rect 11471 23684 11796 23712
rect 11471 23681 11483 23684
rect 11425 23675 11483 23681
rect 3973 23607 4031 23613
rect 4080 23616 4292 23644
rect 4617 23647 4675 23653
rect 2777 23579 2835 23585
rect 2777 23545 2789 23579
rect 2823 23576 2835 23579
rect 2958 23576 2964 23588
rect 2823 23548 2964 23576
rect 2823 23545 2835 23548
rect 2777 23539 2835 23545
rect 2958 23536 2964 23548
rect 3016 23576 3022 23588
rect 3053 23579 3111 23585
rect 3053 23576 3065 23579
rect 3016 23548 3065 23576
rect 3016 23536 3022 23548
rect 3053 23545 3065 23548
rect 3099 23545 3111 23579
rect 3053 23539 3111 23545
rect 3513 23579 3571 23585
rect 3513 23545 3525 23579
rect 3559 23576 3571 23579
rect 4080 23576 4108 23616
rect 4617 23613 4629 23647
rect 4663 23644 4675 23647
rect 5460 23644 5488 23672
rect 4663 23616 5488 23644
rect 5537 23647 5595 23653
rect 4663 23613 4675 23616
rect 4617 23607 4675 23613
rect 5537 23613 5549 23647
rect 5583 23644 5595 23647
rect 6362 23644 6368 23656
rect 5583 23616 6368 23644
rect 5583 23613 5595 23616
rect 5537 23607 5595 23613
rect 3559 23548 4108 23576
rect 5077 23579 5135 23585
rect 3559 23545 3571 23548
rect 3513 23539 3571 23545
rect 5077 23545 5089 23579
rect 5123 23576 5135 23579
rect 5552 23576 5580 23607
rect 6362 23604 6368 23616
rect 6420 23604 6426 23656
rect 6825 23647 6883 23653
rect 6825 23613 6837 23647
rect 6871 23644 6883 23647
rect 7466 23644 7472 23656
rect 6871 23616 7472 23644
rect 6871 23613 6883 23616
rect 6825 23607 6883 23613
rect 7466 23604 7472 23616
rect 7524 23604 7530 23656
rect 8021 23647 8079 23653
rect 8021 23613 8033 23647
rect 8067 23644 8079 23647
rect 8113 23647 8171 23653
rect 8113 23644 8125 23647
rect 8067 23616 8125 23644
rect 8067 23613 8079 23616
rect 8021 23607 8079 23613
rect 8113 23613 8125 23616
rect 8159 23613 8171 23647
rect 8113 23607 8171 23613
rect 8380 23647 8438 23653
rect 8380 23613 8392 23647
rect 8426 23644 8438 23647
rect 8662 23644 8668 23656
rect 8426 23616 8668 23644
rect 8426 23613 8438 23616
rect 8380 23607 8438 23613
rect 5123 23548 5580 23576
rect 5123 23545 5135 23548
rect 5077 23539 5135 23545
rect 5626 23536 5632 23588
rect 5684 23576 5690 23588
rect 6638 23576 6644 23588
rect 5684 23548 6644 23576
rect 5684 23536 5690 23548
rect 6638 23536 6644 23548
rect 6696 23576 6702 23588
rect 8036 23576 8064 23607
rect 8662 23604 8668 23616
rect 8720 23604 8726 23656
rect 11256 23644 11284 23675
rect 11790 23672 11796 23684
rect 11848 23672 11854 23724
rect 13630 23672 13636 23724
rect 13688 23712 13694 23724
rect 13688 23684 15332 23712
rect 13688 23672 13694 23684
rect 12342 23644 12348 23656
rect 11256 23616 12348 23644
rect 12342 23604 12348 23616
rect 12400 23604 12406 23656
rect 12437 23647 12495 23653
rect 12437 23613 12449 23647
rect 12483 23644 12495 23647
rect 15194 23644 15200 23656
rect 12483 23616 15200 23644
rect 12483 23613 12495 23616
rect 12437 23607 12495 23613
rect 6696 23548 8064 23576
rect 6696 23536 6702 23548
rect 10410 23536 10416 23588
rect 10468 23576 10474 23588
rect 10505 23579 10563 23585
rect 10505 23576 10517 23579
rect 10468 23548 10517 23576
rect 10468 23536 10474 23548
rect 10505 23545 10517 23548
rect 10551 23576 10563 23579
rect 11885 23579 11943 23585
rect 11885 23576 11897 23579
rect 10551 23548 11897 23576
rect 10551 23545 10563 23548
rect 10505 23539 10563 23545
rect 11885 23545 11897 23548
rect 11931 23576 11943 23579
rect 12452 23576 12480 23607
rect 15194 23604 15200 23616
rect 15252 23604 15258 23656
rect 15304 23644 15332 23684
rect 17788 23644 17816 23820
rect 20349 23817 20361 23820
rect 20395 23848 20407 23851
rect 21266 23848 21272 23860
rect 20395 23820 21272 23848
rect 20395 23817 20407 23820
rect 20349 23811 20407 23817
rect 21266 23808 21272 23820
rect 21324 23808 21330 23860
rect 21910 23808 21916 23860
rect 21968 23848 21974 23860
rect 22281 23851 22339 23857
rect 22281 23848 22293 23851
rect 21968 23820 22293 23848
rect 21968 23808 21974 23820
rect 22281 23817 22293 23820
rect 22327 23817 22339 23851
rect 24762 23848 24768 23860
rect 24723 23820 24768 23848
rect 22281 23811 22339 23817
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 19334 23740 19340 23792
rect 19392 23780 19398 23792
rect 19392 23752 25360 23780
rect 19392 23740 19398 23752
rect 20622 23672 20628 23724
rect 20680 23672 20686 23724
rect 20714 23672 20720 23724
rect 20772 23712 20778 23724
rect 21177 23715 21235 23721
rect 21177 23712 21189 23715
rect 20772 23684 21189 23712
rect 20772 23672 20778 23684
rect 21177 23681 21189 23684
rect 21223 23712 21235 23715
rect 21818 23712 21824 23724
rect 21223 23684 21824 23712
rect 21223 23681 21235 23684
rect 21177 23675 21235 23681
rect 21818 23672 21824 23684
rect 21876 23672 21882 23724
rect 24118 23672 24124 23724
rect 24176 23712 24182 23724
rect 25133 23715 25191 23721
rect 25133 23712 25145 23715
rect 24176 23684 25145 23712
rect 24176 23672 24182 23684
rect 25133 23681 25145 23684
rect 25179 23681 25191 23715
rect 25133 23675 25191 23681
rect 15304 23616 17816 23644
rect 17865 23647 17923 23653
rect 17865 23613 17877 23647
rect 17911 23644 17923 23647
rect 18049 23647 18107 23653
rect 18049 23644 18061 23647
rect 17911 23616 18061 23644
rect 17911 23613 17923 23616
rect 17865 23607 17923 23613
rect 18049 23613 18061 23616
rect 18095 23644 18107 23647
rect 18138 23644 18144 23656
rect 18095 23616 18144 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 18138 23604 18144 23616
rect 18196 23604 18202 23656
rect 19518 23604 19524 23656
rect 19576 23644 19582 23656
rect 20640 23644 20668 23672
rect 25332 23656 25360 23752
rect 20901 23647 20959 23653
rect 20901 23644 20913 23647
rect 19576 23616 20913 23644
rect 19576 23604 19582 23616
rect 20901 23613 20913 23616
rect 20947 23613 20959 23647
rect 21910 23644 21916 23656
rect 21871 23616 21916 23644
rect 20901 23607 20959 23613
rect 21910 23604 21916 23616
rect 21968 23644 21974 23656
rect 22097 23647 22155 23653
rect 22097 23644 22109 23647
rect 21968 23616 22109 23644
rect 21968 23604 21974 23616
rect 22097 23613 22109 23616
rect 22143 23613 22155 23647
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 22097 23607 22155 23613
rect 24412 23616 24593 23644
rect 11931 23548 12480 23576
rect 11931 23545 11943 23548
rect 11885 23539 11943 23545
rect 12526 23536 12532 23588
rect 12584 23576 12590 23588
rect 12682 23579 12740 23585
rect 12682 23576 12694 23579
rect 12584 23548 12694 23576
rect 12584 23536 12590 23548
rect 12682 23545 12694 23548
rect 12728 23576 12740 23579
rect 13446 23576 13452 23588
rect 12728 23548 13452 23576
rect 12728 23545 12740 23548
rect 12682 23539 12740 23545
rect 13446 23536 13452 23548
rect 13504 23576 13510 23588
rect 13906 23576 13912 23588
rect 13504 23548 13912 23576
rect 13504 23536 13510 23548
rect 13906 23536 13912 23548
rect 13964 23536 13970 23588
rect 15378 23536 15384 23588
rect 15436 23585 15442 23588
rect 15436 23579 15500 23585
rect 15436 23545 15454 23579
rect 15488 23545 15500 23579
rect 18294 23579 18352 23585
rect 18294 23576 18306 23579
rect 15436 23539 15500 23545
rect 17880 23548 18306 23576
rect 15436 23536 15442 23539
rect 17880 23520 17908 23548
rect 18294 23545 18306 23548
rect 18340 23545 18352 23579
rect 18294 23539 18352 23545
rect 20073 23579 20131 23585
rect 20073 23545 20085 23579
rect 20119 23576 20131 23579
rect 20438 23576 20444 23588
rect 20119 23548 20444 23576
rect 20119 23545 20131 23548
rect 20073 23539 20131 23545
rect 20438 23536 20444 23548
rect 20496 23536 20502 23588
rect 20548 23548 21128 23576
rect 1673 23511 1731 23517
rect 1673 23477 1685 23511
rect 1719 23508 1731 23511
rect 1946 23508 1952 23520
rect 1719 23480 1952 23508
rect 1719 23477 1731 23480
rect 1673 23471 1731 23477
rect 1946 23468 1952 23480
rect 2004 23468 2010 23520
rect 7006 23508 7012 23520
rect 6967 23480 7012 23508
rect 7006 23468 7012 23480
rect 7064 23468 7070 23520
rect 9490 23508 9496 23520
rect 9451 23480 9496 23508
rect 9490 23468 9496 23480
rect 9548 23468 9554 23520
rect 10134 23508 10140 23520
rect 10095 23480 10140 23508
rect 10134 23468 10140 23480
rect 10192 23468 10198 23520
rect 10778 23508 10784 23520
rect 10739 23480 10784 23508
rect 10778 23468 10784 23480
rect 10836 23468 10842 23520
rect 11146 23508 11152 23520
rect 11107 23480 11152 23508
rect 11146 23468 11152 23480
rect 11204 23468 11210 23520
rect 13814 23508 13820 23520
rect 13775 23480 13820 23508
rect 13814 23468 13820 23480
rect 13872 23468 13878 23520
rect 13998 23468 14004 23520
rect 14056 23508 14062 23520
rect 16482 23508 16488 23520
rect 14056 23480 16488 23508
rect 14056 23468 14062 23480
rect 16482 23468 16488 23480
rect 16540 23468 16546 23520
rect 17862 23468 17868 23520
rect 17920 23468 17926 23520
rect 19426 23508 19432 23520
rect 19387 23480 19432 23508
rect 19426 23468 19432 23480
rect 19484 23468 19490 23520
rect 20162 23468 20168 23520
rect 20220 23508 20226 23520
rect 20548 23517 20576 23548
rect 20533 23511 20591 23517
rect 20533 23508 20545 23511
rect 20220 23480 20545 23508
rect 20220 23468 20226 23480
rect 20533 23477 20545 23480
rect 20579 23477 20591 23511
rect 20990 23508 20996 23520
rect 20951 23480 20996 23508
rect 20533 23471 20591 23477
rect 20990 23468 20996 23480
rect 21048 23468 21054 23520
rect 21100 23508 21128 23548
rect 21358 23536 21364 23588
rect 21416 23576 21422 23588
rect 21637 23579 21695 23585
rect 21637 23576 21649 23579
rect 21416 23548 21649 23576
rect 21416 23536 21422 23548
rect 21637 23545 21649 23548
rect 21683 23576 21695 23579
rect 22002 23576 22008 23588
rect 21683 23548 22008 23576
rect 21683 23545 21695 23548
rect 21637 23539 21695 23545
rect 22002 23536 22008 23548
rect 22060 23536 22066 23588
rect 22462 23508 22468 23520
rect 21100 23480 22468 23508
rect 22462 23468 22468 23480
rect 22520 23468 22526 23520
rect 22646 23508 22652 23520
rect 22607 23480 22652 23508
rect 22646 23468 22652 23480
rect 22704 23468 22710 23520
rect 24026 23468 24032 23520
rect 24084 23508 24090 23520
rect 24412 23517 24440 23616
rect 24581 23613 24593 23616
rect 24627 23613 24639 23647
rect 24581 23607 24639 23613
rect 25314 23604 25320 23656
rect 25372 23604 25378 23656
rect 24397 23511 24455 23517
rect 24397 23508 24409 23511
rect 24084 23480 24409 23508
rect 24084 23468 24090 23480
rect 24397 23477 24409 23480
rect 24443 23477 24455 23511
rect 24397 23471 24455 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1578 23304 1584 23316
rect 1539 23276 1584 23304
rect 1578 23264 1584 23276
rect 1636 23264 1642 23316
rect 2409 23307 2467 23313
rect 2409 23273 2421 23307
rect 2455 23304 2467 23307
rect 3050 23304 3056 23316
rect 2455 23276 3056 23304
rect 2455 23273 2467 23276
rect 2409 23267 2467 23273
rect 3050 23264 3056 23276
rect 3108 23264 3114 23316
rect 4801 23307 4859 23313
rect 4801 23273 4813 23307
rect 4847 23304 4859 23307
rect 5258 23304 5264 23316
rect 4847 23276 5264 23304
rect 4847 23273 4859 23276
rect 4801 23267 4859 23273
rect 5258 23264 5264 23276
rect 5316 23264 5322 23316
rect 7190 23304 7196 23316
rect 7151 23276 7196 23304
rect 7190 23264 7196 23276
rect 7248 23304 7254 23316
rect 7837 23307 7895 23313
rect 7837 23304 7849 23307
rect 7248 23276 7849 23304
rect 7248 23264 7254 23276
rect 7837 23273 7849 23276
rect 7883 23273 7895 23307
rect 7837 23267 7895 23273
rect 9125 23307 9183 23313
rect 9125 23273 9137 23307
rect 9171 23304 9183 23307
rect 9674 23304 9680 23316
rect 9171 23276 9680 23304
rect 9171 23273 9183 23276
rect 9125 23267 9183 23273
rect 3510 23236 3516 23248
rect 1412 23208 3516 23236
rect 1412 23177 1440 23208
rect 3510 23196 3516 23208
rect 3568 23196 3574 23248
rect 4433 23239 4491 23245
rect 4433 23205 4445 23239
rect 4479 23236 4491 23239
rect 5074 23236 5080 23248
rect 4479 23208 5080 23236
rect 4479 23205 4491 23208
rect 4433 23199 4491 23205
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23137 1455 23171
rect 2774 23168 2780 23180
rect 2735 23140 2780 23168
rect 1397 23131 1455 23137
rect 2774 23128 2780 23140
rect 2832 23128 2838 23180
rect 2869 23171 2927 23177
rect 2869 23137 2881 23171
rect 2915 23168 2927 23171
rect 3234 23168 3240 23180
rect 2915 23140 3240 23168
rect 2915 23137 2927 23140
rect 2869 23131 2927 23137
rect 3234 23128 3240 23140
rect 3292 23128 3298 23180
rect 2317 23103 2375 23109
rect 2317 23069 2329 23103
rect 2363 23100 2375 23103
rect 3053 23103 3111 23109
rect 3053 23100 3065 23103
rect 2363 23072 3065 23100
rect 2363 23069 2375 23072
rect 2317 23063 2375 23069
rect 3053 23069 3065 23072
rect 3099 23100 3111 23103
rect 4448 23100 4476 23199
rect 5074 23196 5080 23208
rect 5132 23245 5138 23248
rect 5132 23239 5196 23245
rect 5132 23205 5150 23239
rect 5184 23205 5196 23239
rect 7852 23236 7880 23267
rect 9674 23264 9680 23276
rect 9732 23304 9738 23316
rect 10045 23307 10103 23313
rect 10045 23304 10057 23307
rect 9732 23276 10057 23304
rect 9732 23264 9738 23276
rect 10045 23273 10057 23276
rect 10091 23273 10103 23307
rect 10045 23267 10103 23273
rect 10873 23307 10931 23313
rect 10873 23273 10885 23307
rect 10919 23304 10931 23307
rect 10962 23304 10968 23316
rect 10919 23276 10968 23304
rect 10919 23273 10931 23276
rect 10873 23267 10931 23273
rect 9490 23236 9496 23248
rect 7852 23208 9496 23236
rect 5132 23199 5196 23205
rect 5132 23196 5138 23199
rect 4893 23171 4951 23177
rect 4893 23137 4905 23171
rect 4939 23168 4951 23171
rect 5442 23168 5448 23180
rect 4939 23140 5448 23168
rect 4939 23137 4951 23140
rect 4893 23131 4951 23137
rect 5442 23128 5448 23140
rect 5500 23168 5506 23180
rect 5626 23168 5632 23180
rect 5500 23140 5632 23168
rect 5500 23128 5506 23140
rect 5626 23128 5632 23140
rect 5684 23128 5690 23180
rect 5994 23128 6000 23180
rect 6052 23128 6058 23180
rect 8389 23171 8447 23177
rect 8389 23168 8401 23171
rect 8312 23140 8401 23168
rect 3099 23072 4476 23100
rect 3099 23069 3111 23072
rect 3053 23063 3111 23069
rect 3510 23032 3516 23044
rect 3471 23004 3516 23032
rect 3510 22992 3516 23004
rect 3568 22992 3574 23044
rect 6012 22976 6040 23128
rect 8018 23032 8024 23044
rect 7979 23004 8024 23032
rect 8018 22992 8024 23004
rect 8076 22992 8082 23044
rect 8312 23032 8340 23140
rect 8389 23137 8401 23140
rect 8435 23137 8447 23171
rect 8389 23131 8447 23137
rect 8478 23100 8484 23112
rect 8439 23072 8484 23100
rect 8478 23060 8484 23072
rect 8536 23060 8542 23112
rect 8588 23109 8616 23208
rect 9490 23196 9496 23208
rect 9548 23196 9554 23248
rect 9674 23128 9680 23180
rect 9732 23168 9738 23180
rect 10137 23171 10195 23177
rect 10137 23168 10149 23171
rect 9732 23140 10149 23168
rect 9732 23128 9738 23140
rect 10137 23137 10149 23140
rect 10183 23137 10195 23171
rect 10137 23131 10195 23137
rect 8573 23103 8631 23109
rect 8573 23069 8585 23103
rect 8619 23069 8631 23103
rect 8573 23063 8631 23069
rect 9030 23032 9036 23044
rect 8312 23004 9036 23032
rect 9030 22992 9036 23004
rect 9088 23032 9094 23044
rect 9677 23035 9735 23041
rect 9677 23032 9689 23035
rect 9088 23004 9689 23032
rect 9088 22992 9094 23004
rect 9677 23001 9689 23004
rect 9723 23001 9735 23035
rect 10152 23032 10180 23131
rect 10318 23100 10324 23112
rect 10231 23072 10324 23100
rect 10318 23060 10324 23072
rect 10376 23100 10382 23112
rect 10888 23100 10916 23267
rect 10962 23264 10968 23276
rect 11020 23264 11026 23316
rect 12345 23307 12403 23313
rect 12345 23273 12357 23307
rect 12391 23304 12403 23307
rect 12526 23304 12532 23316
rect 12391 23276 12532 23304
rect 12391 23273 12403 23276
rect 12345 23267 12403 23273
rect 12526 23264 12532 23276
rect 12584 23264 12590 23316
rect 13078 23264 13084 23316
rect 13136 23304 13142 23316
rect 13173 23307 13231 23313
rect 13173 23304 13185 23307
rect 13136 23276 13185 23304
rect 13136 23264 13142 23276
rect 13173 23273 13185 23276
rect 13219 23273 13231 23307
rect 13173 23267 13231 23273
rect 13265 23307 13323 23313
rect 13265 23273 13277 23307
rect 13311 23304 13323 23307
rect 13722 23304 13728 23316
rect 13311 23276 13728 23304
rect 13311 23273 13323 23276
rect 13265 23267 13323 23273
rect 13722 23264 13728 23276
rect 13780 23264 13786 23316
rect 13906 23304 13912 23316
rect 13867 23276 13912 23304
rect 13906 23264 13912 23276
rect 13964 23264 13970 23316
rect 14826 23264 14832 23316
rect 14884 23304 14890 23316
rect 15013 23307 15071 23313
rect 15013 23304 15025 23307
rect 14884 23276 15025 23304
rect 14884 23264 14890 23276
rect 15013 23273 15025 23276
rect 15059 23273 15071 23307
rect 15013 23267 15071 23273
rect 15473 23307 15531 23313
rect 15473 23273 15485 23307
rect 15519 23304 15531 23307
rect 15562 23304 15568 23316
rect 15519 23276 15568 23304
rect 15519 23273 15531 23276
rect 15473 23267 15531 23273
rect 15562 23264 15568 23276
rect 15620 23264 15626 23316
rect 19429 23307 19487 23313
rect 15672 23276 17080 23304
rect 12802 23196 12808 23248
rect 12860 23236 12866 23248
rect 15672 23236 15700 23276
rect 16758 23245 16764 23248
rect 16752 23236 16764 23245
rect 12860 23208 15700 23236
rect 16719 23208 16764 23236
rect 12860 23196 12866 23208
rect 16752 23199 16764 23208
rect 16758 23196 16764 23199
rect 16816 23196 16822 23248
rect 17052 23236 17080 23276
rect 19429 23273 19441 23307
rect 19475 23304 19487 23307
rect 20162 23304 20168 23316
rect 19475 23276 20168 23304
rect 19475 23273 19487 23276
rect 19429 23267 19487 23273
rect 20162 23264 20168 23276
rect 20220 23264 20226 23316
rect 20438 23264 20444 23316
rect 20496 23304 20502 23316
rect 21818 23304 21824 23316
rect 20496 23276 21824 23304
rect 20496 23264 20502 23276
rect 21818 23264 21824 23276
rect 21876 23304 21882 23316
rect 21913 23307 21971 23313
rect 21913 23304 21925 23307
rect 21876 23276 21925 23304
rect 21876 23264 21882 23276
rect 21913 23273 21925 23276
rect 21959 23273 21971 23307
rect 21913 23267 21971 23273
rect 22002 23264 22008 23316
rect 22060 23304 22066 23316
rect 22646 23304 22652 23316
rect 22060 23276 22652 23304
rect 22060 23264 22066 23276
rect 22646 23264 22652 23276
rect 22704 23264 22710 23316
rect 22738 23264 22744 23316
rect 22796 23304 22802 23316
rect 22925 23307 22983 23313
rect 22925 23304 22937 23307
rect 22796 23276 22937 23304
rect 22796 23264 22802 23276
rect 22925 23273 22937 23276
rect 22971 23273 22983 23307
rect 24762 23304 24768 23316
rect 24723 23276 24768 23304
rect 22925 23267 22983 23273
rect 24762 23264 24768 23276
rect 24820 23264 24826 23316
rect 19886 23236 19892 23248
rect 17052 23208 19892 23236
rect 19886 23196 19892 23208
rect 19944 23196 19950 23248
rect 20254 23196 20260 23248
rect 20312 23236 20318 23248
rect 22278 23236 22284 23248
rect 20312 23208 21496 23236
rect 22239 23208 22284 23236
rect 20312 23196 20318 23208
rect 21468 23180 21496 23208
rect 22278 23196 22284 23208
rect 22336 23196 22342 23248
rect 11054 23128 11060 23180
rect 11112 23168 11118 23180
rect 11609 23171 11667 23177
rect 11609 23168 11621 23171
rect 11112 23140 11621 23168
rect 11112 23128 11118 23140
rect 11609 23137 11621 23140
rect 11655 23137 11667 23171
rect 11609 23131 11667 23137
rect 11701 23171 11759 23177
rect 11701 23137 11713 23171
rect 11747 23168 11759 23171
rect 11882 23168 11888 23180
rect 11747 23140 11888 23168
rect 11747 23137 11759 23140
rect 11701 23131 11759 23137
rect 11882 23128 11888 23140
rect 11940 23128 11946 23180
rect 12894 23128 12900 23180
rect 12952 23168 12958 23180
rect 14553 23171 14611 23177
rect 14553 23168 14565 23171
rect 12952 23140 14565 23168
rect 12952 23128 12958 23140
rect 14553 23137 14565 23140
rect 14599 23137 14611 23171
rect 14553 23131 14611 23137
rect 14734 23128 14740 23180
rect 14792 23168 14798 23180
rect 15289 23171 15347 23177
rect 15289 23168 15301 23171
rect 14792 23140 15301 23168
rect 14792 23128 14798 23140
rect 15289 23137 15301 23140
rect 15335 23168 15347 23171
rect 16206 23168 16212 23180
rect 15335 23140 16212 23168
rect 15335 23137 15347 23140
rect 15289 23131 15347 23137
rect 16206 23128 16212 23140
rect 16264 23128 16270 23180
rect 19334 23128 19340 23180
rect 19392 23168 19398 23180
rect 21266 23168 21272 23180
rect 19392 23140 19437 23168
rect 21227 23140 21272 23168
rect 19392 23128 19398 23140
rect 21266 23128 21272 23140
rect 21324 23128 21330 23180
rect 21450 23168 21456 23180
rect 21363 23140 21456 23168
rect 21450 23128 21456 23140
rect 21508 23168 21514 23180
rect 22830 23168 22836 23180
rect 21508 23140 21588 23168
rect 22791 23140 22836 23168
rect 21508 23128 21514 23140
rect 11790 23100 11796 23112
rect 10376 23072 10916 23100
rect 11751 23072 11796 23100
rect 10376 23060 10382 23072
rect 11790 23060 11796 23072
rect 11848 23060 11854 23112
rect 13354 23100 13360 23112
rect 13315 23072 13360 23100
rect 13354 23060 13360 23072
rect 13412 23100 13418 23112
rect 13814 23100 13820 23112
rect 13412 23072 13820 23100
rect 13412 23060 13418 23072
rect 13814 23060 13820 23072
rect 13872 23100 13878 23112
rect 14185 23103 14243 23109
rect 14185 23100 14197 23103
rect 13872 23072 14197 23100
rect 13872 23060 13878 23072
rect 14185 23069 14197 23072
rect 14231 23069 14243 23103
rect 14185 23063 14243 23069
rect 15194 23060 15200 23112
rect 15252 23100 15258 23112
rect 15933 23103 15991 23109
rect 15933 23100 15945 23103
rect 15252 23072 15945 23100
rect 15252 23060 15258 23072
rect 15933 23069 15945 23072
rect 15979 23100 15991 23103
rect 16482 23100 16488 23112
rect 15979 23072 16488 23100
rect 15979 23069 15991 23072
rect 15933 23063 15991 23069
rect 16482 23060 16488 23072
rect 16540 23060 16546 23112
rect 19521 23103 19579 23109
rect 19521 23100 19533 23103
rect 17880 23072 19533 23100
rect 17880 23044 17908 23072
rect 19521 23069 19533 23072
rect 19567 23100 19579 23103
rect 20162 23100 20168 23112
rect 19567 23072 20168 23100
rect 19567 23069 19579 23072
rect 19521 23063 19579 23069
rect 20162 23060 20168 23072
rect 20220 23060 20226 23112
rect 20714 23060 20720 23112
rect 20772 23100 20778 23112
rect 21560 23109 21588 23140
rect 22830 23128 22836 23140
rect 22888 23128 22894 23180
rect 24581 23171 24639 23177
rect 24581 23137 24593 23171
rect 24627 23168 24639 23171
rect 24670 23168 24676 23180
rect 24627 23140 24676 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 21361 23103 21419 23109
rect 21361 23100 21373 23103
rect 20772 23072 21373 23100
rect 20772 23060 20778 23072
rect 21361 23069 21373 23072
rect 21407 23069 21419 23103
rect 21361 23063 21419 23069
rect 21545 23103 21603 23109
rect 21545 23069 21557 23103
rect 21591 23069 21603 23103
rect 21545 23063 21603 23069
rect 23109 23103 23167 23109
rect 23109 23069 23121 23103
rect 23155 23100 23167 23103
rect 23198 23100 23204 23112
rect 23155 23072 23204 23100
rect 23155 23069 23167 23072
rect 23109 23063 23167 23069
rect 23198 23060 23204 23072
rect 23256 23060 23262 23112
rect 11241 23035 11299 23041
rect 11241 23032 11253 23035
rect 10152 23004 11253 23032
rect 9677 22995 9735 23001
rect 11241 23001 11253 23004
rect 11287 23001 11299 23035
rect 11241 22995 11299 23001
rect 12713 23035 12771 23041
rect 12713 23001 12725 23035
rect 12759 23032 12771 23035
rect 12986 23032 12992 23044
rect 12759 23004 12992 23032
rect 12759 23001 12771 23004
rect 12713 22995 12771 23001
rect 12986 22992 12992 23004
rect 13044 22992 13050 23044
rect 13078 22992 13084 23044
rect 13136 23032 13142 23044
rect 13446 23032 13452 23044
rect 13136 23004 13452 23032
rect 13136 22992 13142 23004
rect 13446 22992 13452 23004
rect 13504 22992 13510 23044
rect 17862 23032 17868 23044
rect 17775 23004 17868 23032
rect 17862 22992 17868 23004
rect 17920 22992 17926 23044
rect 1854 22964 1860 22976
rect 1815 22936 1860 22964
rect 1854 22924 1860 22936
rect 1912 22924 1918 22976
rect 3881 22967 3939 22973
rect 3881 22933 3893 22967
rect 3927 22964 3939 22967
rect 4154 22964 4160 22976
rect 3927 22936 4160 22964
rect 3927 22933 3939 22936
rect 3881 22927 3939 22933
rect 4154 22924 4160 22936
rect 4212 22924 4218 22976
rect 5994 22924 6000 22976
rect 6052 22924 6058 22976
rect 6270 22964 6276 22976
rect 6231 22936 6276 22964
rect 6270 22924 6276 22936
rect 6328 22924 6334 22976
rect 6914 22964 6920 22976
rect 6875 22936 6920 22964
rect 6914 22924 6920 22936
rect 6972 22924 6978 22976
rect 9490 22964 9496 22976
rect 9451 22936 9496 22964
rect 9490 22924 9496 22936
rect 9548 22924 9554 22976
rect 12802 22964 12808 22976
rect 12763 22936 12808 22964
rect 12802 22924 12808 22936
rect 12860 22924 12866 22976
rect 16393 22967 16451 22973
rect 16393 22933 16405 22967
rect 16439 22964 16451 22967
rect 17880 22964 17908 22992
rect 16439 22936 17908 22964
rect 16439 22933 16451 22936
rect 16393 22927 16451 22933
rect 18598 22924 18604 22976
rect 18656 22964 18662 22976
rect 18693 22967 18751 22973
rect 18693 22964 18705 22967
rect 18656 22936 18705 22964
rect 18656 22924 18662 22936
rect 18693 22933 18705 22936
rect 18739 22964 18751 22967
rect 18782 22964 18788 22976
rect 18739 22936 18788 22964
rect 18739 22933 18751 22936
rect 18693 22927 18751 22933
rect 18782 22924 18788 22936
rect 18840 22924 18846 22976
rect 18966 22964 18972 22976
rect 18927 22936 18972 22964
rect 18966 22924 18972 22936
rect 19024 22924 19030 22976
rect 20254 22964 20260 22976
rect 20215 22936 20260 22964
rect 20254 22924 20260 22936
rect 20312 22924 20318 22976
rect 20438 22924 20444 22976
rect 20496 22964 20502 22976
rect 20533 22967 20591 22973
rect 20533 22964 20545 22967
rect 20496 22936 20545 22964
rect 20496 22924 20502 22936
rect 20533 22933 20545 22936
rect 20579 22933 20591 22967
rect 20533 22927 20591 22933
rect 20901 22967 20959 22973
rect 20901 22933 20913 22967
rect 20947 22964 20959 22967
rect 22002 22964 22008 22976
rect 20947 22936 22008 22964
rect 20947 22933 20959 22936
rect 20901 22927 20959 22933
rect 22002 22924 22008 22936
rect 22060 22924 22066 22976
rect 22094 22924 22100 22976
rect 22152 22964 22158 22976
rect 22465 22967 22523 22973
rect 22465 22964 22477 22967
rect 22152 22936 22477 22964
rect 22152 22924 22158 22936
rect 22465 22933 22477 22936
rect 22511 22933 22523 22967
rect 23474 22964 23480 22976
rect 23435 22936 23480 22964
rect 22465 22927 22523 22933
rect 23474 22924 23480 22936
rect 23532 22924 23538 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2041 22763 2099 22769
rect 2041 22760 2053 22763
rect 1412 22732 2053 22760
rect 1412 22565 1440 22732
rect 2041 22729 2053 22732
rect 2087 22760 2099 22763
rect 3878 22760 3884 22772
rect 2087 22732 3884 22760
rect 2087 22729 2099 22732
rect 2041 22723 2099 22729
rect 3878 22720 3884 22732
rect 3936 22720 3942 22772
rect 4982 22720 4988 22772
rect 5040 22760 5046 22772
rect 5350 22760 5356 22772
rect 5040 22732 5356 22760
rect 5040 22720 5046 22732
rect 5350 22720 5356 22732
rect 5408 22720 5414 22772
rect 6822 22760 6828 22772
rect 6783 22732 6828 22760
rect 6822 22720 6828 22732
rect 6880 22720 6886 22772
rect 9398 22720 9404 22772
rect 9456 22760 9462 22772
rect 10318 22760 10324 22772
rect 9456 22732 10324 22760
rect 9456 22720 9462 22732
rect 10318 22720 10324 22732
rect 10376 22720 10382 22772
rect 11054 22760 11060 22772
rect 11015 22732 11060 22760
rect 11054 22720 11060 22732
rect 11112 22720 11118 22772
rect 11422 22760 11428 22772
rect 11383 22732 11428 22760
rect 11422 22720 11428 22732
rect 11480 22720 11486 22772
rect 12434 22720 12440 22772
rect 12492 22760 12498 22772
rect 12492 22732 12537 22760
rect 12492 22720 12498 22732
rect 15378 22720 15384 22772
rect 15436 22760 15442 22772
rect 15657 22763 15715 22769
rect 15657 22760 15669 22763
rect 15436 22732 15669 22760
rect 15436 22720 15442 22732
rect 15657 22729 15669 22732
rect 15703 22729 15715 22763
rect 16206 22760 16212 22772
rect 16167 22732 16212 22760
rect 15657 22723 15715 22729
rect 16206 22720 16212 22732
rect 16264 22720 16270 22772
rect 19518 22760 19524 22772
rect 19479 22732 19524 22760
rect 19518 22720 19524 22732
rect 19576 22760 19582 22772
rect 20070 22760 20076 22772
rect 19576 22732 20076 22760
rect 19576 22720 19582 22732
rect 20070 22720 20076 22732
rect 20128 22720 20134 22772
rect 20990 22760 20996 22772
rect 20951 22732 20996 22760
rect 20990 22720 20996 22732
rect 21048 22720 21054 22772
rect 22830 22760 22836 22772
rect 22791 22732 22836 22760
rect 22830 22720 22836 22732
rect 22888 22720 22894 22772
rect 23842 22760 23848 22772
rect 23803 22732 23848 22760
rect 23842 22720 23848 22732
rect 23900 22720 23906 22772
rect 1581 22695 1639 22701
rect 1581 22661 1593 22695
rect 1627 22692 1639 22695
rect 3050 22692 3056 22704
rect 1627 22664 3056 22692
rect 1627 22661 1639 22664
rect 1581 22655 1639 22661
rect 3050 22652 3056 22664
rect 3108 22652 3114 22704
rect 10134 22652 10140 22704
rect 10192 22692 10198 22704
rect 10781 22695 10839 22701
rect 10781 22692 10793 22695
rect 10192 22664 10793 22692
rect 10192 22652 10198 22664
rect 10781 22661 10793 22664
rect 10827 22692 10839 22695
rect 11790 22692 11796 22704
rect 10827 22664 11796 22692
rect 10827 22661 10839 22664
rect 10781 22655 10839 22661
rect 11790 22652 11796 22664
rect 11848 22692 11854 22704
rect 12253 22695 12311 22701
rect 12253 22692 12265 22695
rect 11848 22664 12265 22692
rect 11848 22652 11854 22664
rect 12253 22661 12265 22664
rect 12299 22692 12311 22695
rect 13354 22692 13360 22704
rect 12299 22664 13360 22692
rect 12299 22661 12311 22664
rect 12253 22655 12311 22661
rect 2774 22584 2780 22636
rect 2832 22624 2838 22636
rect 3142 22624 3148 22636
rect 2832 22596 3004 22624
rect 3103 22596 3148 22624
rect 2832 22584 2838 22596
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22525 1455 22559
rect 1397 22519 1455 22525
rect 2593 22559 2651 22565
rect 2593 22525 2605 22559
rect 2639 22556 2651 22559
rect 2639 22528 2912 22556
rect 2639 22525 2651 22528
rect 2593 22519 2651 22525
rect 1486 22420 1492 22432
rect 1044 22392 1492 22420
rect 1044 22148 1072 22392
rect 1486 22380 1492 22392
rect 1544 22380 1550 22432
rect 1578 22380 1584 22432
rect 1636 22420 1642 22432
rect 2685 22423 2743 22429
rect 2685 22420 2697 22423
rect 1636 22392 2697 22420
rect 1636 22380 1642 22392
rect 2685 22389 2697 22392
rect 2731 22389 2743 22423
rect 2884 22420 2912 22528
rect 2976 22488 3004 22596
rect 3142 22584 3148 22596
rect 3200 22584 3206 22636
rect 3326 22624 3332 22636
rect 3287 22596 3332 22624
rect 3326 22584 3332 22596
rect 3384 22584 3390 22636
rect 6181 22627 6239 22633
rect 6181 22593 6193 22627
rect 6227 22624 6239 22627
rect 7469 22627 7527 22633
rect 7469 22624 7481 22627
rect 6227 22596 7481 22624
rect 6227 22593 6239 22596
rect 6181 22587 6239 22593
rect 7469 22593 7481 22596
rect 7515 22624 7527 22627
rect 7558 22624 7564 22636
rect 7515 22596 7564 22624
rect 7515 22593 7527 22596
rect 7469 22587 7527 22593
rect 7558 22584 7564 22596
rect 7616 22584 7622 22636
rect 8573 22627 8631 22633
rect 8573 22593 8585 22627
rect 8619 22624 8631 22627
rect 8665 22627 8723 22633
rect 8665 22624 8677 22627
rect 8619 22596 8677 22624
rect 8619 22593 8631 22596
rect 8573 22587 8631 22593
rect 8665 22593 8677 22596
rect 8711 22593 8723 22627
rect 11054 22624 11060 22636
rect 8665 22587 8723 22593
rect 9876 22596 11060 22624
rect 3053 22559 3111 22565
rect 3053 22525 3065 22559
rect 3099 22556 3111 22559
rect 3418 22556 3424 22568
rect 3099 22528 3424 22556
rect 3099 22525 3111 22528
rect 3053 22519 3111 22525
rect 3418 22516 3424 22528
rect 3476 22516 3482 22568
rect 4522 22565 4528 22568
rect 4157 22559 4215 22565
rect 4157 22525 4169 22559
rect 4203 22556 4215 22559
rect 4249 22559 4307 22565
rect 4249 22556 4261 22559
rect 4203 22528 4261 22556
rect 4203 22525 4215 22528
rect 4157 22519 4215 22525
rect 4249 22525 4261 22528
rect 4295 22525 4307 22559
rect 4516 22556 4528 22565
rect 4435 22528 4528 22556
rect 4249 22519 4307 22525
rect 4516 22519 4528 22528
rect 4580 22556 4586 22568
rect 6270 22556 6276 22568
rect 4580 22528 6276 22556
rect 3142 22488 3148 22500
rect 2976 22460 3148 22488
rect 3142 22448 3148 22460
rect 3200 22488 3206 22500
rect 3697 22491 3755 22497
rect 3697 22488 3709 22491
rect 3200 22460 3709 22488
rect 3200 22448 3206 22460
rect 3697 22457 3709 22460
rect 3743 22457 3755 22491
rect 4264 22488 4292 22519
rect 4522 22516 4528 22519
rect 4580 22516 4586 22528
rect 6270 22516 6276 22528
rect 6328 22516 6334 22568
rect 6914 22516 6920 22568
rect 6972 22556 6978 22568
rect 7190 22556 7196 22568
rect 6972 22528 7196 22556
rect 6972 22516 6978 22528
rect 7190 22516 7196 22528
rect 7248 22516 7254 22568
rect 8680 22556 8708 22587
rect 9876 22556 9904 22596
rect 11054 22584 11060 22596
rect 11112 22584 11118 22636
rect 12894 22624 12900 22636
rect 12855 22596 12900 22624
rect 12894 22584 12900 22596
rect 12952 22584 12958 22636
rect 13004 22633 13032 22664
rect 13354 22652 13360 22664
rect 13412 22652 13418 22704
rect 17034 22692 17040 22704
rect 16995 22664 17040 22692
rect 17034 22652 17040 22664
rect 17092 22652 17098 22704
rect 17586 22652 17592 22704
rect 17644 22692 17650 22704
rect 17862 22692 17868 22704
rect 17644 22664 17868 22692
rect 17644 22652 17650 22664
rect 17862 22652 17868 22664
rect 17920 22652 17926 22704
rect 19610 22692 19616 22704
rect 19571 22664 19616 22692
rect 19610 22652 19616 22664
rect 19668 22652 19674 22704
rect 19886 22652 19892 22704
rect 19944 22692 19950 22704
rect 20714 22692 20720 22704
rect 19944 22664 20576 22692
rect 20675 22664 20720 22692
rect 19944 22652 19950 22664
rect 12989 22627 13047 22633
rect 12989 22593 13001 22627
rect 13035 22593 13047 22627
rect 12989 22587 13047 22593
rect 14200 22596 14412 22624
rect 10042 22556 10048 22568
rect 8680 22528 9904 22556
rect 9968 22528 10048 22556
rect 9968 22500 9996 22528
rect 10042 22516 10048 22528
rect 10100 22516 10106 22568
rect 11238 22556 11244 22568
rect 11151 22528 11244 22556
rect 11238 22516 11244 22528
rect 11296 22556 11302 22568
rect 11974 22556 11980 22568
rect 11296 22528 11980 22556
rect 11296 22516 11302 22528
rect 11974 22516 11980 22528
rect 12032 22516 12038 22568
rect 12710 22516 12716 22568
rect 12768 22556 12774 22568
rect 12805 22559 12863 22565
rect 12805 22556 12817 22559
rect 12768 22528 12817 22556
rect 12768 22516 12774 22528
rect 12805 22525 12817 22528
rect 12851 22525 12863 22559
rect 12805 22519 12863 22525
rect 13354 22516 13360 22568
rect 13412 22556 13418 22568
rect 13538 22556 13544 22568
rect 13412 22528 13544 22556
rect 13412 22516 13418 22528
rect 13538 22516 13544 22528
rect 13596 22516 13602 22568
rect 4706 22488 4712 22500
rect 4264 22460 4712 22488
rect 3697 22451 3755 22457
rect 4706 22448 4712 22460
rect 4764 22448 4770 22500
rect 6641 22491 6699 22497
rect 6641 22457 6653 22491
rect 6687 22488 6699 22491
rect 7006 22488 7012 22500
rect 6687 22460 7012 22488
rect 6687 22457 6699 22460
rect 6641 22451 6699 22457
rect 7006 22448 7012 22460
rect 7064 22488 7070 22500
rect 7285 22491 7343 22497
rect 7285 22488 7297 22491
rect 7064 22460 7297 22488
rect 7064 22448 7070 22460
rect 7285 22457 7297 22460
rect 7331 22488 7343 22491
rect 7374 22488 7380 22500
rect 7331 22460 7380 22488
rect 7331 22457 7343 22460
rect 7285 22451 7343 22457
rect 7374 22448 7380 22460
rect 7432 22448 7438 22500
rect 7926 22448 7932 22500
rect 7984 22488 7990 22500
rect 8938 22497 8944 22500
rect 8205 22491 8263 22497
rect 8205 22488 8217 22491
rect 7984 22460 8217 22488
rect 7984 22448 7990 22460
rect 8205 22457 8217 22460
rect 8251 22488 8263 22491
rect 8932 22488 8944 22497
rect 8251 22460 8944 22488
rect 8251 22457 8263 22460
rect 8205 22451 8263 22457
rect 8932 22451 8944 22460
rect 8938 22448 8944 22451
rect 8996 22448 9002 22500
rect 9950 22448 9956 22500
rect 10008 22448 10014 22500
rect 10778 22448 10784 22500
rect 10836 22488 10842 22500
rect 14200 22488 14228 22596
rect 14277 22559 14335 22565
rect 14277 22525 14289 22559
rect 14323 22525 14335 22559
rect 14384 22556 14412 22596
rect 18046 22584 18052 22636
rect 18104 22624 18110 22636
rect 18506 22624 18512 22636
rect 18104 22596 18512 22624
rect 18104 22584 18110 22596
rect 18506 22584 18512 22596
rect 18564 22584 18570 22636
rect 18690 22624 18696 22636
rect 18603 22596 18696 22624
rect 18690 22584 18696 22596
rect 18748 22624 18754 22636
rect 19426 22624 19432 22636
rect 18748 22596 19432 22624
rect 18748 22584 18754 22596
rect 19426 22584 19432 22596
rect 19484 22584 19490 22636
rect 20257 22627 20315 22633
rect 20257 22593 20269 22627
rect 20303 22624 20315 22627
rect 20438 22624 20444 22636
rect 20303 22596 20444 22624
rect 20303 22593 20315 22596
rect 20257 22587 20315 22593
rect 20438 22584 20444 22596
rect 20496 22584 20502 22636
rect 16298 22556 16304 22568
rect 14384 22528 16304 22556
rect 14277 22519 14335 22525
rect 10836 22460 14228 22488
rect 10836 22448 10842 22460
rect 3326 22420 3332 22432
rect 2884 22392 3332 22420
rect 2685 22383 2743 22389
rect 3326 22380 3332 22392
rect 3384 22380 3390 22432
rect 3786 22380 3792 22432
rect 3844 22420 3850 22432
rect 5258 22420 5264 22432
rect 3844 22392 5264 22420
rect 3844 22380 3850 22392
rect 5258 22380 5264 22392
rect 5316 22380 5322 22432
rect 5626 22420 5632 22432
rect 5587 22392 5632 22420
rect 5626 22380 5632 22392
rect 5684 22380 5690 22432
rect 6270 22380 6276 22432
rect 6328 22420 6334 22432
rect 6546 22420 6552 22432
rect 6328 22392 6552 22420
rect 6328 22380 6334 22392
rect 6546 22380 6552 22392
rect 6604 22380 6610 22432
rect 10042 22420 10048 22432
rect 10003 22392 10048 22420
rect 10042 22380 10048 22392
rect 10100 22380 10106 22432
rect 11882 22420 11888 22432
rect 11843 22392 11888 22420
rect 11882 22380 11888 22392
rect 11940 22380 11946 22432
rect 13446 22420 13452 22432
rect 13407 22392 13452 22420
rect 13446 22380 13452 22392
rect 13504 22380 13510 22432
rect 13538 22380 13544 22432
rect 13596 22420 13602 22432
rect 13722 22420 13728 22432
rect 13596 22392 13728 22420
rect 13596 22380 13602 22392
rect 13722 22380 13728 22392
rect 13780 22380 13786 22432
rect 14182 22420 14188 22432
rect 14095 22392 14188 22420
rect 14182 22380 14188 22392
rect 14240 22420 14246 22432
rect 14292 22420 14320 22519
rect 16298 22516 16304 22528
rect 16356 22556 16362 22568
rect 16853 22559 16911 22565
rect 16853 22556 16865 22559
rect 16356 22528 16865 22556
rect 16356 22516 16362 22528
rect 16853 22525 16865 22528
rect 16899 22556 16911 22559
rect 17405 22559 17463 22565
rect 17405 22556 17417 22559
rect 16899 22528 17417 22556
rect 16899 22525 16911 22528
rect 16853 22519 16911 22525
rect 17405 22525 17417 22528
rect 17451 22525 17463 22559
rect 17405 22519 17463 22525
rect 17862 22516 17868 22568
rect 17920 22556 17926 22568
rect 18417 22559 18475 22565
rect 18417 22556 18429 22559
rect 17920 22528 18429 22556
rect 17920 22516 17926 22528
rect 18417 22525 18429 22528
rect 18463 22556 18475 22559
rect 18966 22556 18972 22568
rect 18463 22528 18972 22556
rect 18463 22525 18475 22528
rect 18417 22519 18475 22525
rect 18966 22516 18972 22528
rect 19024 22516 19030 22568
rect 19242 22516 19248 22568
rect 19300 22556 19306 22568
rect 19794 22556 19800 22568
rect 19300 22528 19800 22556
rect 19300 22516 19306 22528
rect 19794 22516 19800 22528
rect 19852 22516 19858 22568
rect 20070 22556 20076 22568
rect 20031 22528 20076 22556
rect 20070 22516 20076 22528
rect 20128 22516 20134 22568
rect 20548 22556 20576 22664
rect 20714 22652 20720 22664
rect 20772 22652 20778 22704
rect 22557 22695 22615 22701
rect 22557 22661 22569 22695
rect 22603 22692 22615 22695
rect 22738 22692 22744 22704
rect 22603 22664 22744 22692
rect 22603 22661 22615 22664
rect 22557 22655 22615 22661
rect 22738 22652 22744 22664
rect 22796 22652 22802 22704
rect 21450 22584 21456 22636
rect 21508 22624 21514 22636
rect 21729 22627 21787 22633
rect 21729 22624 21741 22627
rect 21508 22596 21741 22624
rect 21508 22584 21514 22596
rect 21729 22593 21741 22596
rect 21775 22593 21787 22627
rect 21729 22587 21787 22593
rect 20714 22556 20720 22568
rect 20548 22528 20720 22556
rect 20714 22516 20720 22528
rect 20772 22516 20778 22568
rect 20990 22516 20996 22568
rect 21048 22556 21054 22568
rect 21545 22559 21603 22565
rect 21545 22556 21557 22559
rect 21048 22528 21557 22556
rect 21048 22516 21054 22528
rect 21545 22525 21557 22528
rect 21591 22525 21603 22559
rect 21545 22519 21603 22525
rect 21637 22559 21695 22565
rect 21637 22525 21649 22559
rect 21683 22556 21695 22559
rect 21818 22556 21824 22568
rect 21683 22528 21824 22556
rect 21683 22525 21695 22528
rect 21637 22519 21695 22525
rect 14544 22491 14602 22497
rect 14544 22457 14556 22491
rect 14590 22488 14602 22491
rect 14642 22488 14648 22500
rect 14590 22460 14648 22488
rect 14590 22457 14602 22460
rect 14544 22451 14602 22457
rect 14642 22448 14648 22460
rect 14700 22448 14706 22500
rect 16482 22448 16488 22500
rect 16540 22488 16546 22500
rect 16669 22491 16727 22497
rect 16669 22488 16681 22491
rect 16540 22460 16681 22488
rect 16540 22448 16546 22460
rect 16669 22457 16681 22460
rect 16715 22488 16727 22491
rect 18138 22488 18144 22500
rect 16715 22460 18144 22488
rect 16715 22457 16727 22460
rect 16669 22451 16727 22457
rect 18138 22448 18144 22460
rect 18196 22448 18202 22500
rect 19153 22491 19211 22497
rect 19153 22457 19165 22491
rect 19199 22488 19211 22491
rect 19981 22491 20039 22497
rect 19981 22488 19993 22491
rect 19199 22460 19993 22488
rect 19199 22457 19211 22460
rect 19153 22451 19211 22457
rect 19981 22457 19993 22460
rect 20027 22488 20039 22491
rect 21652 22488 21680 22519
rect 21818 22516 21824 22528
rect 21876 22516 21882 22568
rect 23658 22556 23664 22568
rect 23619 22528 23664 22556
rect 23658 22516 23664 22528
rect 23716 22556 23722 22568
rect 24213 22559 24271 22565
rect 24213 22556 24225 22559
rect 23716 22528 24225 22556
rect 23716 22516 23722 22528
rect 24213 22525 24225 22528
rect 24259 22525 24271 22559
rect 24213 22519 24271 22525
rect 24670 22488 24676 22500
rect 20027 22460 21680 22488
rect 24631 22460 24676 22488
rect 20027 22457 20039 22460
rect 19981 22451 20039 22457
rect 24670 22448 24676 22460
rect 24728 22448 24734 22500
rect 15286 22420 15292 22432
rect 14240 22392 15292 22420
rect 14240 22380 14246 22392
rect 15286 22380 15292 22392
rect 15344 22380 15350 22432
rect 18046 22420 18052 22432
rect 18007 22392 18052 22420
rect 18046 22380 18052 22392
rect 18104 22380 18110 22432
rect 18230 22380 18236 22432
rect 18288 22420 18294 22432
rect 20990 22420 20996 22432
rect 18288 22392 20996 22420
rect 18288 22380 18294 22392
rect 20990 22380 20996 22392
rect 21048 22380 21054 22432
rect 21177 22423 21235 22429
rect 21177 22389 21189 22423
rect 21223 22420 21235 22423
rect 21358 22420 21364 22432
rect 21223 22392 21364 22420
rect 21223 22389 21235 22392
rect 21177 22383 21235 22389
rect 21358 22380 21364 22392
rect 21416 22380 21422 22432
rect 23198 22420 23204 22432
rect 23159 22392 23204 22420
rect 23198 22380 23204 22392
rect 23256 22380 23262 22432
rect 24762 22420 24768 22432
rect 24723 22392 24768 22420
rect 24762 22380 24768 22392
rect 24820 22380 24826 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1854 22176 1860 22228
rect 1912 22216 1918 22228
rect 1912 22188 2452 22216
rect 1912 22176 1918 22188
rect 1765 22151 1823 22157
rect 1765 22148 1777 22151
rect 1044 22120 1777 22148
rect 1765 22117 1777 22120
rect 1811 22148 1823 22151
rect 2225 22151 2283 22157
rect 2225 22148 2237 22151
rect 1811 22120 2237 22148
rect 1811 22117 1823 22120
rect 1765 22111 1823 22117
rect 2225 22117 2237 22120
rect 2271 22117 2283 22151
rect 2225 22111 2283 22117
rect 1026 22040 1032 22092
rect 1084 22080 1090 22092
rect 1486 22080 1492 22092
rect 1084 22052 1492 22080
rect 1084 22040 1090 22052
rect 1486 22040 1492 22052
rect 1544 22040 1550 22092
rect 1118 21972 1124 22024
rect 1176 22012 1182 22024
rect 2424 22021 2452 22188
rect 4062 22176 4068 22228
rect 4120 22216 4126 22228
rect 4338 22216 4344 22228
rect 4120 22188 4344 22216
rect 4120 22176 4126 22188
rect 4338 22176 4344 22188
rect 4396 22216 4402 22228
rect 4801 22219 4859 22225
rect 4801 22216 4813 22219
rect 4396 22188 4813 22216
rect 4396 22176 4402 22188
rect 4801 22185 4813 22188
rect 4847 22185 4859 22219
rect 5442 22216 5448 22228
rect 5403 22188 5448 22216
rect 4801 22179 4859 22185
rect 5442 22176 5448 22188
rect 5500 22176 5506 22228
rect 6178 22176 6184 22228
rect 6236 22216 6242 22228
rect 6825 22219 6883 22225
rect 6825 22216 6837 22219
rect 6236 22188 6837 22216
rect 6236 22176 6242 22188
rect 6825 22185 6837 22188
rect 6871 22185 6883 22219
rect 6825 22179 6883 22185
rect 8021 22219 8079 22225
rect 8021 22185 8033 22219
rect 8067 22216 8079 22219
rect 8202 22216 8208 22228
rect 8067 22188 8208 22216
rect 8067 22185 8079 22188
rect 8021 22179 8079 22185
rect 8202 22176 8208 22188
rect 8260 22176 8266 22228
rect 9858 22216 9864 22228
rect 9819 22188 9864 22216
rect 9858 22176 9864 22188
rect 9916 22176 9922 22228
rect 10321 22219 10379 22225
rect 10321 22185 10333 22219
rect 10367 22216 10379 22219
rect 10686 22216 10692 22228
rect 10367 22188 10692 22216
rect 10367 22185 10379 22188
rect 10321 22179 10379 22185
rect 10686 22176 10692 22188
rect 10744 22176 10750 22228
rect 13538 22216 13544 22228
rect 13499 22188 13544 22216
rect 13538 22176 13544 22188
rect 13596 22176 13602 22228
rect 13740 22188 14044 22216
rect 2958 22108 2964 22160
rect 3016 22148 3022 22160
rect 3016 22120 3648 22148
rect 3016 22108 3022 22120
rect 3234 22040 3240 22092
rect 3292 22040 3298 22092
rect 2317 22015 2375 22021
rect 2317 22012 2329 22015
rect 1176 21984 2329 22012
rect 1176 21972 1182 21984
rect 2317 21981 2329 21984
rect 2363 21981 2375 22015
rect 2317 21975 2375 21981
rect 2409 22015 2467 22021
rect 2409 21981 2421 22015
rect 2455 22012 2467 22015
rect 2774 22012 2780 22024
rect 2455 21984 2780 22012
rect 2455 21981 2467 21984
rect 2409 21975 2467 21981
rect 2774 21972 2780 21984
rect 2832 21972 2838 22024
rect 1857 21947 1915 21953
rect 1857 21913 1869 21947
rect 1903 21944 1915 21947
rect 1946 21944 1952 21956
rect 1903 21916 1952 21944
rect 1903 21913 1915 21916
rect 1857 21907 1915 21913
rect 1946 21904 1952 21916
rect 2004 21904 2010 21956
rect 3252 21888 3280 22040
rect 3620 22024 3648 22120
rect 4706 22108 4712 22160
rect 4764 22148 4770 22160
rect 5460 22148 5488 22176
rect 4764 22120 5488 22148
rect 4764 22108 4770 22120
rect 5626 22108 5632 22160
rect 5684 22148 5690 22160
rect 8386 22148 8392 22160
rect 5684 22120 6592 22148
rect 8347 22120 8392 22148
rect 5684 22108 5690 22120
rect 4341 22083 4399 22089
rect 4341 22049 4353 22083
rect 4387 22080 4399 22083
rect 4522 22080 4528 22092
rect 4387 22052 4528 22080
rect 4387 22049 4399 22052
rect 4341 22043 4399 22049
rect 4522 22040 4528 22052
rect 4580 22040 4586 22092
rect 6362 22080 6368 22092
rect 6323 22052 6368 22080
rect 6362 22040 6368 22052
rect 6420 22040 6426 22092
rect 3602 21972 3608 22024
rect 3660 21972 3666 22024
rect 4154 21972 4160 22024
rect 4212 22012 4218 22024
rect 4890 22012 4896 22024
rect 4212 21984 4896 22012
rect 4212 21972 4218 21984
rect 4890 21972 4896 21984
rect 4948 21972 4954 22024
rect 4982 21972 4988 22024
rect 5040 22012 5046 22024
rect 6564 22012 6592 22120
rect 8386 22108 8392 22120
rect 8444 22108 8450 22160
rect 10042 22108 10048 22160
rect 10100 22148 10106 22160
rect 10100 22120 11008 22148
rect 10100 22108 10106 22120
rect 9398 22080 9404 22092
rect 9359 22052 9404 22080
rect 9398 22040 9404 22052
rect 9456 22040 9462 22092
rect 9674 22080 9680 22092
rect 9635 22052 9680 22080
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 10980 22080 11008 22120
rect 12710 22108 12716 22160
rect 12768 22148 12774 22160
rect 13740 22148 13768 22188
rect 13906 22148 13912 22160
rect 12768 22120 13768 22148
rect 13867 22120 13912 22148
rect 12768 22108 12774 22120
rect 13906 22108 13912 22120
rect 13964 22108 13970 22160
rect 11330 22089 11336 22092
rect 11324 22080 11336 22089
rect 10980 22052 11336 22080
rect 11324 22043 11336 22052
rect 11330 22040 11336 22043
rect 11388 22040 11394 22092
rect 14016 22080 14044 22188
rect 16114 22176 16120 22228
rect 16172 22216 16178 22228
rect 16298 22216 16304 22228
rect 16172 22188 16304 22216
rect 16172 22176 16178 22188
rect 16298 22176 16304 22188
rect 16356 22176 16362 22228
rect 16758 22176 16764 22228
rect 16816 22216 16822 22228
rect 16942 22216 16948 22228
rect 16816 22188 16948 22216
rect 16816 22176 16822 22188
rect 16942 22176 16948 22188
rect 17000 22176 17006 22228
rect 17770 22176 17776 22228
rect 17828 22216 17834 22228
rect 18509 22219 18567 22225
rect 18509 22216 18521 22219
rect 17828 22188 18521 22216
rect 17828 22176 17834 22188
rect 18509 22185 18521 22188
rect 18555 22185 18567 22219
rect 18509 22179 18567 22185
rect 19337 22219 19395 22225
rect 19337 22185 19349 22219
rect 19383 22216 19395 22219
rect 20070 22216 20076 22228
rect 19383 22188 20076 22216
rect 19383 22185 19395 22188
rect 19337 22179 19395 22185
rect 20070 22176 20076 22188
rect 20128 22176 20134 22228
rect 20254 22216 20260 22228
rect 20215 22188 20260 22216
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 20901 22219 20959 22225
rect 20901 22185 20913 22219
rect 20947 22216 20959 22219
rect 21266 22216 21272 22228
rect 20947 22188 21272 22216
rect 20947 22185 20959 22188
rect 20901 22179 20959 22185
rect 21266 22176 21272 22188
rect 21324 22176 21330 22228
rect 22002 22216 22008 22228
rect 21376 22188 22008 22216
rect 16482 22148 16488 22160
rect 15304 22120 16488 22148
rect 15304 22092 15332 22120
rect 16482 22108 16488 22120
rect 16540 22108 16546 22160
rect 18049 22151 18107 22157
rect 18049 22117 18061 22151
rect 18095 22148 18107 22151
rect 18690 22148 18696 22160
rect 18095 22120 18696 22148
rect 18095 22117 18107 22120
rect 18049 22111 18107 22117
rect 18524 22092 18552 22120
rect 18690 22108 18696 22120
rect 18748 22108 18754 22160
rect 20346 22108 20352 22160
rect 20404 22148 20410 22160
rect 20441 22151 20499 22157
rect 20441 22148 20453 22151
rect 20404 22120 20453 22148
rect 20404 22108 20410 22120
rect 20441 22117 20453 22120
rect 20487 22117 20499 22151
rect 20441 22111 20499 22117
rect 14921 22083 14979 22089
rect 14921 22080 14933 22083
rect 14016 22052 14933 22080
rect 14921 22049 14933 22052
rect 14967 22049 14979 22083
rect 15286 22080 15292 22092
rect 15199 22052 15292 22080
rect 14921 22043 14979 22049
rect 15286 22040 15292 22052
rect 15344 22040 15350 22092
rect 15556 22083 15614 22089
rect 15556 22049 15568 22083
rect 15602 22080 15614 22083
rect 15838 22080 15844 22092
rect 15602 22052 15844 22080
rect 15602 22049 15614 22052
rect 15556 22043 15614 22049
rect 15838 22040 15844 22052
rect 15896 22040 15902 22092
rect 15930 22040 15936 22092
rect 15988 22080 15994 22092
rect 15988 22052 16528 22080
rect 15988 22040 15994 22052
rect 6638 22012 6644 22024
rect 5040 21984 5085 22012
rect 6564 21984 6644 22012
rect 5040 21972 5046 21984
rect 6638 21972 6644 21984
rect 6696 21972 6702 22024
rect 6730 21972 6736 22024
rect 6788 22012 6794 22024
rect 6917 22015 6975 22021
rect 6917 22012 6929 22015
rect 6788 21984 6929 22012
rect 6788 21972 6794 21984
rect 6917 21981 6929 21984
rect 6963 21981 6975 22015
rect 7098 22012 7104 22024
rect 7059 21984 7104 22012
rect 6917 21975 6975 21981
rect 7098 21972 7104 21984
rect 7156 21972 7162 22024
rect 8478 22012 8484 22024
rect 8439 21984 8484 22012
rect 8478 21972 8484 21984
rect 8536 21972 8542 22024
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 21981 8631 22015
rect 8573 21975 8631 21981
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 22012 9183 22015
rect 9582 22012 9588 22024
rect 9171 21984 9588 22012
rect 9171 21981 9183 21984
rect 9125 21975 9183 21981
rect 6454 21944 6460 21956
rect 6415 21916 6460 21944
rect 6454 21904 6460 21916
rect 6512 21904 6518 21956
rect 8294 21904 8300 21956
rect 8352 21944 8358 21956
rect 8588 21944 8616 21975
rect 9582 21972 9588 21984
rect 9640 21972 9646 22024
rect 11054 22012 11060 22024
rect 11015 21984 11060 22012
rect 11054 21972 11060 21984
rect 11112 21972 11118 22024
rect 13998 22012 14004 22024
rect 13959 21984 14004 22012
rect 13998 21972 14004 21984
rect 14056 21972 14062 22024
rect 14093 22015 14151 22021
rect 14093 21981 14105 22015
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 8352 21916 8616 21944
rect 12437 21947 12495 21953
rect 8352 21904 8358 21916
rect 12437 21913 12449 21947
rect 12483 21944 12495 21947
rect 12526 21944 12532 21956
rect 12483 21916 12532 21944
rect 12483 21913 12495 21916
rect 12437 21907 12495 21913
rect 12526 21904 12532 21916
rect 12584 21944 12590 21956
rect 12802 21944 12808 21956
rect 12584 21916 12808 21944
rect 12584 21904 12590 21916
rect 12802 21904 12808 21916
rect 12860 21944 12866 21956
rect 14108 21944 14136 21975
rect 16500 21956 16528 22052
rect 16942 22040 16948 22092
rect 17000 22080 17006 22092
rect 17221 22083 17279 22089
rect 17221 22080 17233 22083
rect 17000 22052 17233 22080
rect 17000 22040 17006 22052
rect 17221 22049 17233 22052
rect 17267 22049 17279 22083
rect 17221 22043 17279 22049
rect 17494 22040 17500 22092
rect 17552 22040 17558 22092
rect 17681 22083 17739 22089
rect 17681 22049 17693 22083
rect 17727 22080 17739 22083
rect 17862 22080 17868 22092
rect 17727 22052 17868 22080
rect 17727 22049 17739 22052
rect 17681 22043 17739 22049
rect 17862 22040 17868 22052
rect 17920 22040 17926 22092
rect 18506 22040 18512 22092
rect 18564 22040 18570 22092
rect 18874 22040 18880 22092
rect 18932 22080 18938 22092
rect 19702 22080 19708 22092
rect 18932 22052 19288 22080
rect 19663 22052 19708 22080
rect 18932 22040 18938 22052
rect 17126 21972 17132 22024
rect 17184 22012 17190 22024
rect 17512 22012 17540 22040
rect 18598 22012 18604 22024
rect 17184 21984 17540 22012
rect 18559 21984 18604 22012
rect 17184 21972 17190 21984
rect 18598 21972 18604 21984
rect 18656 21972 18662 22024
rect 18690 21972 18696 22024
rect 18748 22012 18754 22024
rect 18748 21984 18793 22012
rect 18748 21972 18754 21984
rect 19150 21972 19156 22024
rect 19208 21972 19214 22024
rect 19260 22012 19288 22052
rect 19702 22040 19708 22052
rect 19760 22040 19766 22092
rect 20162 22040 20168 22092
rect 20220 22080 20226 22092
rect 20714 22080 20720 22092
rect 20220 22052 20720 22080
rect 20220 22040 20226 22052
rect 20714 22040 20720 22052
rect 20772 22040 20778 22092
rect 20254 22012 20260 22024
rect 19260 21984 20260 22012
rect 20254 21972 20260 21984
rect 20312 21972 20318 22024
rect 20346 21972 20352 22024
rect 20404 22012 20410 22024
rect 21376 22012 21404 22188
rect 22002 22176 22008 22188
rect 22060 22176 22066 22228
rect 22462 22216 22468 22228
rect 22423 22188 22468 22216
rect 22462 22176 22468 22188
rect 22520 22176 22526 22228
rect 22649 22219 22707 22225
rect 22649 22185 22661 22219
rect 22695 22185 22707 22219
rect 23014 22216 23020 22228
rect 22975 22188 23020 22216
rect 22649 22179 22707 22185
rect 21453 22151 21511 22157
rect 21453 22117 21465 22151
rect 21499 22148 21511 22151
rect 22097 22151 22155 22157
rect 22097 22148 22109 22151
rect 21499 22120 22109 22148
rect 21499 22117 21511 22120
rect 21453 22111 21511 22117
rect 22097 22117 22109 22120
rect 22143 22148 22155 22151
rect 22664 22148 22692 22179
rect 23014 22176 23020 22188
rect 23072 22176 23078 22228
rect 22143 22120 22692 22148
rect 24581 22151 24639 22157
rect 22143 22117 22155 22120
rect 22097 22111 22155 22117
rect 24581 22117 24593 22151
rect 24627 22148 24639 22151
rect 24627 22120 24808 22148
rect 24627 22117 24639 22120
rect 24581 22111 24639 22117
rect 22830 22040 22836 22092
rect 22888 22080 22894 22092
rect 24026 22080 24032 22092
rect 22888 22052 24032 22080
rect 22888 22040 22894 22052
rect 24026 22040 24032 22052
rect 24084 22040 24090 22092
rect 24780 22080 24808 22120
rect 24854 22080 24860 22092
rect 24780 22052 24860 22080
rect 24854 22040 24860 22052
rect 24912 22080 24918 22092
rect 25222 22080 25228 22092
rect 24912 22052 25228 22080
rect 24912 22040 24918 22052
rect 25222 22040 25228 22052
rect 25280 22040 25286 22092
rect 21545 22015 21603 22021
rect 21545 22012 21557 22015
rect 20404 21984 21557 22012
rect 20404 21972 20410 21984
rect 21545 21981 21557 21984
rect 21591 21981 21603 22015
rect 21726 22012 21732 22024
rect 21687 21984 21732 22012
rect 21545 21975 21603 21981
rect 21726 21972 21732 21984
rect 21784 21972 21790 22024
rect 22738 21972 22744 22024
rect 22796 22012 22802 22024
rect 23109 22015 23167 22021
rect 23109 22012 23121 22015
rect 22796 21984 23121 22012
rect 22796 21972 22802 21984
rect 23109 21981 23121 21984
rect 23155 21981 23167 22015
rect 23290 22012 23296 22024
rect 23251 21984 23296 22012
rect 23109 21975 23167 21981
rect 23290 21972 23296 21984
rect 23348 21972 23354 22024
rect 24118 22012 24124 22024
rect 23584 21984 24124 22012
rect 12860 21916 14136 21944
rect 12860 21904 12866 21916
rect 16482 21904 16488 21956
rect 16540 21904 16546 21956
rect 17494 21904 17500 21956
rect 17552 21944 17558 21956
rect 17678 21944 17684 21956
rect 17552 21916 17684 21944
rect 17552 21904 17558 21916
rect 17678 21904 17684 21916
rect 17736 21904 17742 21956
rect 18141 21947 18199 21953
rect 18141 21913 18153 21947
rect 18187 21944 18199 21947
rect 19168 21944 19196 21972
rect 19337 21947 19395 21953
rect 19337 21944 19349 21947
rect 18187 21916 19196 21944
rect 19260 21916 19349 21944
rect 18187 21913 18199 21916
rect 18141 21907 18199 21913
rect 19260 21888 19288 21916
rect 19337 21913 19349 21916
rect 19383 21913 19395 21947
rect 19337 21907 19395 21913
rect 19613 21947 19671 21953
rect 19613 21913 19625 21947
rect 19659 21944 19671 21947
rect 19794 21944 19800 21956
rect 19659 21916 19800 21944
rect 19659 21913 19671 21916
rect 19613 21907 19671 21913
rect 19794 21904 19800 21916
rect 19852 21904 19858 21956
rect 20070 21904 20076 21956
rect 20128 21944 20134 21956
rect 23584 21944 23612 21984
rect 24118 21972 24124 21984
rect 24176 21972 24182 22024
rect 24210 21972 24216 22024
rect 24268 22012 24274 22024
rect 24673 22015 24731 22021
rect 24673 22012 24685 22015
rect 24268 21984 24685 22012
rect 24268 21972 24274 21984
rect 24673 21981 24685 21984
rect 24719 21981 24731 22015
rect 24673 21975 24731 21981
rect 24765 22015 24823 22021
rect 24765 21981 24777 22015
rect 24811 21981 24823 22015
rect 24765 21975 24823 21981
rect 20128 21916 23612 21944
rect 20128 21904 20134 21916
rect 23934 21904 23940 21956
rect 23992 21944 23998 21956
rect 24780 21944 24808 21975
rect 23992 21916 24808 21944
rect 23992 21904 23998 21916
rect 2961 21879 3019 21885
rect 2961 21845 2973 21879
rect 3007 21876 3019 21879
rect 3234 21876 3240 21888
rect 3007 21848 3240 21876
rect 3007 21845 3019 21848
rect 2961 21839 3019 21845
rect 3234 21836 3240 21848
rect 3292 21836 3298 21888
rect 3510 21876 3516 21888
rect 3471 21848 3516 21876
rect 3510 21836 3516 21848
rect 3568 21836 3574 21888
rect 3786 21876 3792 21888
rect 3747 21848 3792 21876
rect 3786 21836 3792 21848
rect 3844 21876 3850 21888
rect 4433 21879 4491 21885
rect 4433 21876 4445 21879
rect 3844 21848 4445 21876
rect 3844 21836 3850 21848
rect 4433 21845 4445 21848
rect 4479 21845 4491 21879
rect 4433 21839 4491 21845
rect 5997 21879 6055 21885
rect 5997 21845 6009 21879
rect 6043 21876 6055 21879
rect 6086 21876 6092 21888
rect 6043 21848 6092 21876
rect 6043 21845 6055 21848
rect 5997 21839 6055 21845
rect 6086 21836 6092 21848
rect 6144 21836 6150 21888
rect 6362 21836 6368 21888
rect 6420 21876 6426 21888
rect 7282 21876 7288 21888
rect 6420 21848 7288 21876
rect 6420 21836 6426 21848
rect 7282 21836 7288 21848
rect 7340 21836 7346 21888
rect 7558 21836 7564 21888
rect 7616 21876 7622 21888
rect 7653 21879 7711 21885
rect 7653 21876 7665 21879
rect 7616 21848 7665 21876
rect 7616 21836 7622 21848
rect 7653 21845 7665 21848
rect 7699 21845 7711 21879
rect 7653 21839 7711 21845
rect 10134 21836 10140 21888
rect 10192 21876 10198 21888
rect 10597 21879 10655 21885
rect 10597 21876 10609 21879
rect 10192 21848 10609 21876
rect 10192 21836 10198 21848
rect 10597 21845 10609 21848
rect 10643 21845 10655 21879
rect 10597 21839 10655 21845
rect 13262 21836 13268 21888
rect 13320 21876 13326 21888
rect 13357 21879 13415 21885
rect 13357 21876 13369 21879
rect 13320 21848 13369 21876
rect 13320 21836 13326 21848
rect 13357 21845 13369 21848
rect 13403 21876 13415 21879
rect 14182 21876 14188 21888
rect 13403 21848 14188 21876
rect 13403 21845 13415 21848
rect 13357 21839 13415 21845
rect 14182 21836 14188 21848
rect 14240 21836 14246 21888
rect 14642 21876 14648 21888
rect 14555 21848 14648 21876
rect 14642 21836 14648 21848
rect 14700 21876 14706 21888
rect 16669 21879 16727 21885
rect 16669 21876 16681 21879
rect 14700 21848 16681 21876
rect 14700 21836 14706 21848
rect 16669 21845 16681 21848
rect 16715 21845 16727 21879
rect 19242 21876 19248 21888
rect 19203 21848 19248 21876
rect 16669 21839 16727 21845
rect 19242 21836 19248 21848
rect 19300 21836 19306 21888
rect 19886 21876 19892 21888
rect 19847 21848 19892 21876
rect 19886 21836 19892 21848
rect 19944 21836 19950 21888
rect 20441 21879 20499 21885
rect 20441 21845 20453 21879
rect 20487 21876 20499 21879
rect 20530 21876 20536 21888
rect 20487 21848 20536 21876
rect 20487 21845 20499 21848
rect 20441 21839 20499 21845
rect 20530 21836 20536 21848
rect 20588 21836 20594 21888
rect 20714 21876 20720 21888
rect 20675 21848 20720 21876
rect 20714 21836 20720 21848
rect 20772 21876 20778 21888
rect 20901 21879 20959 21885
rect 20901 21876 20913 21879
rect 20772 21848 20913 21876
rect 20772 21836 20778 21848
rect 20901 21845 20913 21848
rect 20947 21845 20959 21879
rect 20901 21839 20959 21845
rect 21085 21879 21143 21885
rect 21085 21845 21097 21879
rect 21131 21876 21143 21879
rect 22002 21876 22008 21888
rect 21131 21848 22008 21876
rect 21131 21845 21143 21848
rect 21085 21839 21143 21845
rect 22002 21836 22008 21848
rect 22060 21836 22066 21888
rect 23750 21876 23756 21888
rect 23711 21848 23756 21876
rect 23750 21836 23756 21848
rect 23808 21836 23814 21888
rect 24026 21876 24032 21888
rect 23987 21848 24032 21876
rect 24026 21836 24032 21848
rect 24084 21836 24090 21888
rect 24118 21836 24124 21888
rect 24176 21876 24182 21888
rect 24213 21879 24271 21885
rect 24213 21876 24225 21879
rect 24176 21848 24225 21876
rect 24176 21836 24182 21848
rect 24213 21845 24225 21848
rect 24259 21845 24271 21879
rect 24213 21839 24271 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1302 21632 1308 21684
rect 1360 21672 1366 21684
rect 1673 21675 1731 21681
rect 1673 21672 1685 21675
rect 1360 21644 1685 21672
rect 1360 21632 1366 21644
rect 1673 21641 1685 21644
rect 1719 21641 1731 21675
rect 1854 21672 1860 21684
rect 1815 21644 1860 21672
rect 1673 21635 1731 21641
rect 1688 21536 1716 21635
rect 1854 21632 1860 21644
rect 1912 21632 1918 21684
rect 4890 21632 4896 21684
rect 4948 21672 4954 21684
rect 4985 21675 5043 21681
rect 4985 21672 4997 21675
rect 4948 21644 4997 21672
rect 4948 21632 4954 21644
rect 4985 21641 4997 21644
rect 5031 21641 5043 21675
rect 4985 21635 5043 21641
rect 5074 21632 5080 21684
rect 5132 21672 5138 21684
rect 5132 21644 8616 21672
rect 5132 21632 5138 21644
rect 3237 21607 3295 21613
rect 3237 21604 3249 21607
rect 2332 21576 3249 21604
rect 2332 21545 2360 21576
rect 3237 21573 3249 21576
rect 3283 21573 3295 21607
rect 3418 21604 3424 21616
rect 3379 21576 3424 21604
rect 3237 21567 3295 21573
rect 2317 21539 2375 21545
rect 2317 21536 2329 21539
rect 1688 21508 2329 21536
rect 2317 21505 2329 21508
rect 2363 21505 2375 21539
rect 2317 21499 2375 21505
rect 2501 21539 2559 21545
rect 2501 21505 2513 21539
rect 2547 21536 2559 21539
rect 2774 21536 2780 21548
rect 2547 21508 2780 21536
rect 2547 21505 2559 21508
rect 2501 21499 2559 21505
rect 2774 21496 2780 21508
rect 2832 21496 2838 21548
rect 658 21428 664 21480
rect 716 21468 722 21480
rect 2225 21471 2283 21477
rect 2225 21468 2237 21471
rect 716 21440 2237 21468
rect 716 21428 722 21440
rect 2225 21437 2237 21440
rect 2271 21468 2283 21471
rect 2869 21471 2927 21477
rect 2869 21468 2881 21471
rect 2271 21440 2881 21468
rect 2271 21437 2283 21440
rect 2225 21431 2283 21437
rect 2869 21437 2881 21440
rect 2915 21437 2927 21471
rect 3252 21468 3280 21567
rect 3418 21564 3424 21576
rect 3476 21564 3482 21616
rect 3878 21564 3884 21616
rect 3936 21604 3942 21616
rect 6822 21604 6828 21616
rect 3936 21576 6828 21604
rect 3936 21564 3942 21576
rect 6822 21564 6828 21576
rect 6880 21564 6886 21616
rect 8588 21604 8616 21644
rect 8938 21632 8944 21684
rect 8996 21672 9002 21684
rect 9033 21675 9091 21681
rect 9033 21672 9045 21675
rect 8996 21644 9045 21672
rect 8996 21632 9002 21644
rect 9033 21641 9045 21644
rect 9079 21641 9091 21675
rect 9033 21635 9091 21641
rect 10137 21675 10195 21681
rect 10137 21641 10149 21675
rect 10183 21672 10195 21675
rect 11054 21672 11060 21684
rect 10183 21644 11060 21672
rect 10183 21641 10195 21644
rect 10137 21635 10195 21641
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 11330 21632 11336 21684
rect 11388 21672 11394 21684
rect 11517 21675 11575 21681
rect 11517 21672 11529 21675
rect 11388 21644 11529 21672
rect 11388 21632 11394 21644
rect 11517 21641 11529 21644
rect 11563 21641 11575 21675
rect 11517 21635 11575 21641
rect 11882 21632 11888 21684
rect 11940 21672 11946 21684
rect 12618 21672 12624 21684
rect 11940 21644 12624 21672
rect 11940 21632 11946 21644
rect 12618 21632 12624 21644
rect 12676 21632 12682 21684
rect 12802 21672 12808 21684
rect 12763 21644 12808 21672
rect 12802 21632 12808 21644
rect 12860 21632 12866 21684
rect 13173 21675 13231 21681
rect 13173 21641 13185 21675
rect 13219 21672 13231 21675
rect 13998 21672 14004 21684
rect 13219 21644 14004 21672
rect 13219 21641 13231 21644
rect 13173 21635 13231 21641
rect 9214 21604 9220 21616
rect 8588 21576 9220 21604
rect 9214 21564 9220 21576
rect 9272 21564 9278 21616
rect 9674 21564 9680 21616
rect 9732 21604 9738 21616
rect 9769 21607 9827 21613
rect 9769 21604 9781 21607
rect 9732 21576 9781 21604
rect 9732 21564 9738 21576
rect 9769 21573 9781 21576
rect 9815 21604 9827 21607
rect 13188 21604 13216 21635
rect 13998 21632 14004 21644
rect 14056 21632 14062 21684
rect 15286 21672 15292 21684
rect 15247 21644 15292 21672
rect 15286 21632 15292 21644
rect 15344 21632 15350 21684
rect 16758 21632 16764 21684
rect 16816 21672 16822 21684
rect 17034 21672 17040 21684
rect 16816 21644 17040 21672
rect 16816 21632 16822 21644
rect 17034 21632 17040 21644
rect 17092 21632 17098 21684
rect 17497 21675 17555 21681
rect 17497 21641 17509 21675
rect 17543 21672 17555 21675
rect 18046 21672 18052 21684
rect 17543 21644 18052 21672
rect 17543 21641 17555 21644
rect 17497 21635 17555 21641
rect 18046 21632 18052 21644
rect 18104 21672 18110 21684
rect 18598 21672 18604 21684
rect 18104 21644 18604 21672
rect 18104 21632 18110 21644
rect 18598 21632 18604 21644
rect 18656 21632 18662 21684
rect 19702 21632 19708 21684
rect 19760 21672 19766 21684
rect 20533 21675 20591 21681
rect 20533 21672 20545 21675
rect 19760 21644 20545 21672
rect 19760 21632 19766 21644
rect 20533 21641 20545 21644
rect 20579 21641 20591 21675
rect 21082 21672 21088 21684
rect 21043 21644 21088 21672
rect 20533 21635 20591 21641
rect 21082 21632 21088 21644
rect 21140 21632 21146 21684
rect 23014 21672 23020 21684
rect 22975 21644 23020 21672
rect 23014 21632 23020 21644
rect 23072 21632 23078 21684
rect 24854 21632 24860 21684
rect 24912 21672 24918 21684
rect 25041 21675 25099 21681
rect 25041 21672 25053 21675
rect 24912 21644 25053 21672
rect 24912 21632 24918 21644
rect 25041 21641 25053 21644
rect 25087 21641 25099 21675
rect 25406 21672 25412 21684
rect 25367 21644 25412 21672
rect 25041 21635 25099 21641
rect 25406 21632 25412 21644
rect 25464 21632 25470 21684
rect 9815 21576 13216 21604
rect 9815 21573 9827 21576
rect 9769 21567 9827 21573
rect 21450 21564 21456 21616
rect 21508 21604 21514 21616
rect 23290 21604 23296 21616
rect 21508 21576 23296 21604
rect 21508 21564 21514 21576
rect 23290 21564 23296 21576
rect 23348 21604 23354 21616
rect 23385 21607 23443 21613
rect 23385 21604 23397 21607
rect 23348 21576 23397 21604
rect 23348 21564 23354 21576
rect 23385 21573 23397 21576
rect 23431 21573 23443 21607
rect 23385 21567 23443 21573
rect 23750 21564 23756 21616
rect 23808 21604 23814 21616
rect 23808 21576 24348 21604
rect 23808 21564 23814 21576
rect 3510 21496 3516 21548
rect 3568 21536 3574 21548
rect 3973 21539 4031 21545
rect 3973 21536 3985 21539
rect 3568 21508 3985 21536
rect 3568 21496 3574 21508
rect 3973 21505 3985 21508
rect 4019 21505 4031 21539
rect 3973 21499 4031 21505
rect 4525 21539 4583 21545
rect 4525 21505 4537 21539
rect 4571 21536 4583 21539
rect 5534 21536 5540 21548
rect 4571 21508 5540 21536
rect 4571 21505 4583 21508
rect 4525 21499 4583 21505
rect 3881 21471 3939 21477
rect 3881 21468 3893 21471
rect 3252 21440 3893 21468
rect 2869 21431 2927 21437
rect 3881 21437 3893 21440
rect 3927 21437 3939 21471
rect 3988 21468 4016 21499
rect 5534 21496 5540 21508
rect 5592 21496 5598 21548
rect 9858 21496 9864 21548
rect 9916 21536 9922 21548
rect 10689 21539 10747 21545
rect 10689 21536 10701 21539
rect 9916 21508 10701 21536
rect 9916 21496 9922 21508
rect 10689 21505 10701 21508
rect 10735 21536 10747 21539
rect 11885 21539 11943 21545
rect 11885 21536 11897 21539
rect 10735 21508 11897 21536
rect 10735 21505 10747 21508
rect 10689 21499 10747 21505
rect 11885 21505 11897 21508
rect 11931 21505 11943 21539
rect 13262 21536 13268 21548
rect 13223 21508 13268 21536
rect 11885 21499 11943 21505
rect 13262 21496 13268 21508
rect 13320 21496 13326 21548
rect 16301 21539 16359 21545
rect 16301 21505 16313 21539
rect 16347 21536 16359 21539
rect 17037 21539 17095 21545
rect 17037 21536 17049 21539
rect 16347 21508 17049 21536
rect 16347 21505 16359 21508
rect 16301 21499 16359 21505
rect 17037 21505 17049 21508
rect 17083 21536 17095 21539
rect 17586 21536 17592 21548
rect 17083 21508 17592 21536
rect 17083 21505 17095 21508
rect 17037 21499 17095 21505
rect 17586 21496 17592 21508
rect 17644 21496 17650 21548
rect 18138 21496 18144 21548
rect 18196 21536 18202 21548
rect 18598 21536 18604 21548
rect 18196 21508 18604 21536
rect 18196 21496 18202 21508
rect 18598 21496 18604 21508
rect 18656 21496 18662 21548
rect 19794 21496 19800 21548
rect 19852 21536 19858 21548
rect 20438 21536 20444 21548
rect 19852 21508 20444 21536
rect 19852 21496 19858 21508
rect 20438 21496 20444 21508
rect 20496 21536 20502 21548
rect 20898 21536 20904 21548
rect 20496 21508 20904 21536
rect 20496 21496 20502 21508
rect 20898 21496 20904 21508
rect 20956 21536 20962 21548
rect 21729 21539 21787 21545
rect 21729 21536 21741 21539
rect 20956 21508 21741 21536
rect 20956 21496 20962 21508
rect 21729 21505 21741 21508
rect 21775 21536 21787 21539
rect 22370 21536 22376 21548
rect 21775 21508 22376 21536
rect 21775 21505 21787 21508
rect 21729 21499 21787 21505
rect 22370 21496 22376 21508
rect 22428 21496 22434 21548
rect 24026 21496 24032 21548
rect 24084 21536 24090 21548
rect 24320 21545 24348 21576
rect 24121 21539 24179 21545
rect 24121 21536 24133 21539
rect 24084 21508 24133 21536
rect 24084 21496 24090 21508
rect 24121 21505 24133 21508
rect 24167 21505 24179 21539
rect 24121 21499 24179 21505
rect 24305 21539 24363 21545
rect 24305 21505 24317 21539
rect 24351 21536 24363 21539
rect 24394 21536 24400 21548
rect 24351 21508 24400 21536
rect 24351 21505 24363 21508
rect 24305 21499 24363 21505
rect 24394 21496 24400 21508
rect 24452 21496 24458 21548
rect 6089 21471 6147 21477
rect 6089 21468 6101 21471
rect 3988 21440 6101 21468
rect 3881 21431 3939 21437
rect 6089 21437 6101 21440
rect 6135 21468 6147 21471
rect 7098 21468 7104 21480
rect 6135 21440 7104 21468
rect 6135 21437 6147 21440
rect 6089 21431 6147 21437
rect 3896 21400 3924 21431
rect 7098 21428 7104 21440
rect 7156 21428 7162 21480
rect 7558 21428 7564 21480
rect 7616 21468 7622 21480
rect 7653 21471 7711 21477
rect 7653 21468 7665 21471
rect 7616 21440 7665 21468
rect 7616 21428 7622 21440
rect 7653 21437 7665 21440
rect 7699 21437 7711 21471
rect 7653 21431 7711 21437
rect 9674 21428 9680 21480
rect 9732 21468 9738 21480
rect 11146 21468 11152 21480
rect 9732 21440 11152 21468
rect 9732 21428 9738 21440
rect 11146 21428 11152 21440
rect 11204 21468 11210 21480
rect 11241 21471 11299 21477
rect 11241 21468 11253 21471
rect 11204 21440 11253 21468
rect 11204 21428 11210 21440
rect 11241 21437 11253 21440
rect 11287 21468 11299 21471
rect 13280 21468 13308 21496
rect 16390 21468 16396 21480
rect 11287 21440 13308 21468
rect 13464 21440 16396 21468
rect 11287 21437 11299 21440
rect 11241 21431 11299 21437
rect 4801 21403 4859 21409
rect 4801 21400 4813 21403
rect 3896 21372 4813 21400
rect 4801 21369 4813 21372
rect 4847 21400 4859 21403
rect 5353 21403 5411 21409
rect 5353 21400 5365 21403
rect 4847 21372 5365 21400
rect 4847 21369 4859 21372
rect 4801 21363 4859 21369
rect 5353 21369 5365 21372
rect 5399 21369 5411 21403
rect 5353 21363 5411 21369
rect 6178 21360 6184 21412
rect 6236 21400 6242 21412
rect 7009 21403 7067 21409
rect 7009 21400 7021 21403
rect 6236 21372 7021 21400
rect 6236 21360 6242 21372
rect 7009 21369 7021 21372
rect 7055 21369 7067 21403
rect 7116 21400 7144 21428
rect 7898 21403 7956 21409
rect 7898 21400 7910 21403
rect 7116 21372 7910 21400
rect 7009 21363 7067 21369
rect 7898 21369 7910 21372
rect 7944 21400 7956 21403
rect 8294 21400 8300 21412
rect 7944 21372 8300 21400
rect 7944 21369 7956 21372
rect 7898 21363 7956 21369
rect 8294 21360 8300 21372
rect 8352 21360 8358 21412
rect 10597 21403 10655 21409
rect 10597 21369 10609 21403
rect 10643 21400 10655 21403
rect 10686 21400 10692 21412
rect 10643 21372 10692 21400
rect 10643 21369 10655 21372
rect 10597 21363 10655 21369
rect 10686 21360 10692 21372
rect 10744 21360 10750 21412
rect 11790 21360 11796 21412
rect 11848 21400 11854 21412
rect 13464 21400 13492 21440
rect 16390 21428 16396 21440
rect 16448 21468 16454 21480
rect 16761 21471 16819 21477
rect 16761 21468 16773 21471
rect 16448 21440 16773 21468
rect 16448 21428 16454 21440
rect 16761 21437 16773 21440
rect 16807 21437 16819 21471
rect 16761 21431 16819 21437
rect 17865 21471 17923 21477
rect 17865 21437 17877 21471
rect 17911 21468 17923 21471
rect 18690 21468 18696 21480
rect 17911 21440 18696 21468
rect 17911 21437 17923 21440
rect 17865 21431 17923 21437
rect 18690 21428 18696 21440
rect 18748 21428 18754 21480
rect 21174 21428 21180 21480
rect 21232 21468 21238 21480
rect 21453 21471 21511 21477
rect 21453 21468 21465 21471
rect 21232 21440 21465 21468
rect 21232 21428 21238 21440
rect 21453 21437 21465 21440
rect 21499 21468 21511 21471
rect 23014 21468 23020 21480
rect 21499 21440 23020 21468
rect 21499 21437 21511 21440
rect 21453 21431 21511 21437
rect 23014 21428 23020 21440
rect 23072 21428 23078 21480
rect 25225 21471 25283 21477
rect 25225 21437 25237 21471
rect 25271 21468 25283 21471
rect 25271 21440 25820 21468
rect 25271 21437 25283 21440
rect 25225 21431 25283 21437
rect 11848 21372 13492 21400
rect 13532 21403 13590 21409
rect 11848 21360 11854 21372
rect 13532 21369 13544 21403
rect 13578 21400 13590 21403
rect 13998 21400 14004 21412
rect 13578 21372 14004 21400
rect 13578 21369 13590 21372
rect 13532 21363 13590 21369
rect 13998 21360 14004 21372
rect 14056 21400 14062 21412
rect 14458 21400 14464 21412
rect 14056 21372 14464 21400
rect 14056 21360 14062 21372
rect 14458 21360 14464 21372
rect 14516 21360 14522 21412
rect 16666 21400 16672 21412
rect 14559 21372 16672 21400
rect 2038 21292 2044 21344
rect 2096 21332 2102 21344
rect 2590 21332 2596 21344
rect 2096 21304 2596 21332
rect 2096 21292 2102 21304
rect 2590 21292 2596 21304
rect 2648 21292 2654 21344
rect 3510 21292 3516 21344
rect 3568 21332 3574 21344
rect 3789 21335 3847 21341
rect 3789 21332 3801 21335
rect 3568 21304 3801 21332
rect 3568 21292 3574 21304
rect 3789 21301 3801 21304
rect 3835 21301 3847 21335
rect 3789 21295 3847 21301
rect 5442 21292 5448 21344
rect 5500 21332 5506 21344
rect 6549 21335 6607 21341
rect 5500 21304 5545 21332
rect 5500 21292 5506 21304
rect 6549 21301 6561 21335
rect 6595 21332 6607 21335
rect 6730 21332 6736 21344
rect 6595 21304 6736 21332
rect 6595 21301 6607 21304
rect 6549 21295 6607 21301
rect 6730 21292 6736 21304
rect 6788 21292 6794 21344
rect 7561 21335 7619 21341
rect 7561 21301 7573 21335
rect 7607 21332 7619 21335
rect 8386 21332 8392 21344
rect 7607 21304 8392 21332
rect 7607 21301 7619 21304
rect 7561 21295 7619 21301
rect 8386 21292 8392 21304
rect 8444 21292 8450 21344
rect 10134 21292 10140 21344
rect 10192 21332 10198 21344
rect 10505 21335 10563 21341
rect 10505 21332 10517 21335
rect 10192 21304 10517 21332
rect 10192 21292 10198 21304
rect 10505 21301 10517 21304
rect 10551 21301 10563 21335
rect 10505 21295 10563 21301
rect 10870 21292 10876 21344
rect 10928 21332 10934 21344
rect 14559 21332 14587 21372
rect 16666 21360 16672 21372
rect 16724 21360 16730 21412
rect 18506 21360 18512 21412
rect 18564 21400 18570 21412
rect 18846 21403 18904 21409
rect 18846 21400 18858 21403
rect 18564 21372 18858 21400
rect 18564 21360 18570 21372
rect 18846 21369 18858 21372
rect 18892 21369 18904 21403
rect 18846 21363 18904 21369
rect 21082 21360 21088 21412
rect 21140 21400 21146 21412
rect 21910 21400 21916 21412
rect 21140 21372 21916 21400
rect 21140 21360 21146 21372
rect 21910 21360 21916 21372
rect 21968 21360 21974 21412
rect 23934 21360 23940 21412
rect 23992 21400 23998 21412
rect 24029 21403 24087 21409
rect 24029 21400 24041 21403
rect 23992 21372 24041 21400
rect 23992 21360 23998 21372
rect 24029 21369 24041 21372
rect 24075 21369 24087 21403
rect 24029 21363 24087 21369
rect 25792 21344 25820 21440
rect 10928 21304 14587 21332
rect 14645 21335 14703 21341
rect 10928 21292 10934 21304
rect 14645 21301 14657 21335
rect 14691 21332 14703 21335
rect 14734 21332 14740 21344
rect 14691 21304 14740 21332
rect 14691 21301 14703 21304
rect 14645 21295 14703 21301
rect 14734 21292 14740 21304
rect 14792 21332 14798 21344
rect 15657 21335 15715 21341
rect 15657 21332 15669 21335
rect 14792 21304 15669 21332
rect 14792 21292 14798 21304
rect 15657 21301 15669 21304
rect 15703 21332 15715 21335
rect 15838 21332 15844 21344
rect 15703 21304 15844 21332
rect 15703 21301 15715 21304
rect 15657 21295 15715 21301
rect 15838 21292 15844 21304
rect 15896 21292 15902 21344
rect 16390 21332 16396 21344
rect 16351 21304 16396 21332
rect 16390 21292 16396 21304
rect 16448 21292 16454 21344
rect 16853 21335 16911 21341
rect 16853 21301 16865 21335
rect 16899 21332 16911 21335
rect 17034 21332 17040 21344
rect 16899 21304 17040 21332
rect 16899 21301 16911 21304
rect 16853 21295 16911 21301
rect 17034 21292 17040 21304
rect 17092 21332 17098 21344
rect 17862 21332 17868 21344
rect 17092 21304 17868 21332
rect 17092 21292 17098 21304
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 18417 21335 18475 21341
rect 18417 21301 18429 21335
rect 18463 21332 18475 21335
rect 18598 21332 18604 21344
rect 18463 21304 18604 21332
rect 18463 21301 18475 21304
rect 18417 21295 18475 21301
rect 18598 21292 18604 21304
rect 18656 21292 18662 21344
rect 18690 21292 18696 21344
rect 18748 21332 18754 21344
rect 19334 21332 19340 21344
rect 18748 21304 19340 21332
rect 18748 21292 18754 21304
rect 19334 21292 19340 21304
rect 19392 21332 19398 21344
rect 19981 21335 20039 21341
rect 19981 21332 19993 21335
rect 19392 21304 19993 21332
rect 19392 21292 19398 21304
rect 19981 21301 19993 21304
rect 20027 21301 20039 21335
rect 19981 21295 20039 21301
rect 20622 21292 20628 21344
rect 20680 21332 20686 21344
rect 20901 21335 20959 21341
rect 20901 21332 20913 21335
rect 20680 21304 20913 21332
rect 20680 21292 20686 21304
rect 20901 21301 20913 21304
rect 20947 21332 20959 21335
rect 21545 21335 21603 21341
rect 21545 21332 21557 21335
rect 20947 21304 21557 21332
rect 20947 21301 20959 21304
rect 20901 21295 20959 21301
rect 21545 21301 21557 21304
rect 21591 21301 21603 21335
rect 21545 21295 21603 21301
rect 21726 21292 21732 21344
rect 21784 21332 21790 21344
rect 22097 21335 22155 21341
rect 22097 21332 22109 21335
rect 21784 21304 22109 21332
rect 21784 21292 21790 21304
rect 22097 21301 22109 21304
rect 22143 21332 22155 21335
rect 22462 21332 22468 21344
rect 22143 21304 22468 21332
rect 22143 21301 22155 21304
rect 22097 21295 22155 21301
rect 22462 21292 22468 21304
rect 22520 21292 22526 21344
rect 22738 21332 22744 21344
rect 22699 21304 22744 21332
rect 22738 21292 22744 21304
rect 22796 21292 22802 21344
rect 23661 21335 23719 21341
rect 23661 21301 23673 21335
rect 23707 21332 23719 21335
rect 23750 21332 23756 21344
rect 23707 21304 23756 21332
rect 23707 21301 23719 21304
rect 23661 21295 23719 21301
rect 23750 21292 23756 21304
rect 23808 21292 23814 21344
rect 24578 21292 24584 21344
rect 24636 21332 24642 21344
rect 24673 21335 24731 21341
rect 24673 21332 24685 21335
rect 24636 21304 24685 21332
rect 24636 21292 24642 21304
rect 24673 21301 24685 21304
rect 24719 21301 24731 21335
rect 25774 21332 25780 21344
rect 25735 21304 25780 21332
rect 24673 21295 24731 21301
rect 25774 21292 25780 21304
rect 25832 21292 25838 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1118 21088 1124 21140
rect 1176 21128 1182 21140
rect 1765 21131 1823 21137
rect 1765 21128 1777 21131
rect 1176 21100 1777 21128
rect 1176 21088 1182 21100
rect 1765 21097 1777 21100
rect 1811 21097 1823 21131
rect 1765 21091 1823 21097
rect 1949 21131 2007 21137
rect 1949 21097 1961 21131
rect 1995 21128 2007 21131
rect 2314 21128 2320 21140
rect 1995 21100 2320 21128
rect 1995 21097 2007 21100
rect 1949 21091 2007 21097
rect 1780 21060 1808 21091
rect 2314 21088 2320 21100
rect 2372 21088 2378 21140
rect 2409 21131 2467 21137
rect 2409 21097 2421 21131
rect 2455 21128 2467 21131
rect 3142 21128 3148 21140
rect 2455 21100 3148 21128
rect 2455 21097 2467 21100
rect 2409 21091 2467 21097
rect 3142 21088 3148 21100
rect 3200 21088 3206 21140
rect 4062 21128 4068 21140
rect 4023 21100 4068 21128
rect 4062 21088 4068 21100
rect 4120 21088 4126 21140
rect 5442 21128 5448 21140
rect 5403 21100 5448 21128
rect 5442 21088 5448 21100
rect 5500 21128 5506 21140
rect 5629 21131 5687 21137
rect 5629 21128 5641 21131
rect 5500 21100 5641 21128
rect 5500 21088 5506 21100
rect 5629 21097 5641 21100
rect 5675 21097 5687 21131
rect 7098 21128 7104 21140
rect 7059 21100 7104 21128
rect 5629 21091 5687 21097
rect 7098 21088 7104 21100
rect 7156 21088 7162 21140
rect 8294 21128 8300 21140
rect 8255 21100 8300 21128
rect 8294 21088 8300 21100
rect 8352 21128 8358 21140
rect 9030 21128 9036 21140
rect 8352 21100 8423 21128
rect 8991 21100 9036 21128
rect 8352 21088 8358 21100
rect 3326 21060 3332 21072
rect 1780 21032 3332 21060
rect 3326 21020 3332 21032
rect 3384 21060 3390 21072
rect 4525 21063 4583 21069
rect 4525 21060 4537 21063
rect 3384 21032 4537 21060
rect 3384 21020 3390 21032
rect 4525 21029 4537 21032
rect 4571 21029 4583 21063
rect 4525 21023 4583 21029
rect 6086 21020 6092 21072
rect 6144 21060 6150 21072
rect 7653 21063 7711 21069
rect 7653 21060 7665 21063
rect 6144 21032 7665 21060
rect 6144 21020 6150 21032
rect 7653 21029 7665 21032
rect 7699 21060 7711 21063
rect 8202 21060 8208 21072
rect 7699 21032 8208 21060
rect 7699 21029 7711 21032
rect 7653 21023 7711 21029
rect 8202 21020 8208 21032
rect 8260 21020 8266 21072
rect 8395 21060 8423 21100
rect 9030 21088 9036 21100
rect 9088 21088 9094 21140
rect 11790 21128 11796 21140
rect 11751 21100 11796 21128
rect 11790 21088 11796 21100
rect 11848 21088 11854 21140
rect 12250 21128 12256 21140
rect 12211 21100 12256 21128
rect 12250 21088 12256 21100
rect 12308 21088 12314 21140
rect 13630 21128 13636 21140
rect 13591 21100 13636 21128
rect 13630 21088 13636 21100
rect 13688 21088 13694 21140
rect 14274 21128 14280 21140
rect 14235 21100 14280 21128
rect 14274 21088 14280 21100
rect 14332 21088 14338 21140
rect 14550 21088 14556 21140
rect 14608 21128 14614 21140
rect 15746 21128 15752 21140
rect 14608 21100 15752 21128
rect 14608 21088 14614 21100
rect 15746 21088 15752 21100
rect 15804 21088 15810 21140
rect 16853 21131 16911 21137
rect 16853 21097 16865 21131
rect 16899 21128 16911 21131
rect 17402 21128 17408 21140
rect 16899 21100 17408 21128
rect 16899 21097 16911 21100
rect 16853 21091 16911 21097
rect 17402 21088 17408 21100
rect 17460 21088 17466 21140
rect 17589 21131 17647 21137
rect 17589 21097 17601 21131
rect 17635 21128 17647 21131
rect 18049 21131 18107 21137
rect 18049 21128 18061 21131
rect 17635 21100 18061 21128
rect 17635 21097 17647 21100
rect 17589 21091 17647 21097
rect 18049 21097 18061 21100
rect 18095 21128 18107 21131
rect 19245 21131 19303 21137
rect 19245 21128 19257 21131
rect 18095 21100 19257 21128
rect 18095 21097 18107 21100
rect 18049 21091 18107 21097
rect 19245 21097 19257 21100
rect 19291 21097 19303 21131
rect 20346 21128 20352 21140
rect 20307 21100 20352 21128
rect 19245 21091 19303 21097
rect 20346 21088 20352 21100
rect 20404 21088 20410 21140
rect 20717 21131 20775 21137
rect 20717 21097 20729 21131
rect 20763 21128 20775 21131
rect 20898 21128 20904 21140
rect 20763 21100 20904 21128
rect 20763 21097 20775 21100
rect 20717 21091 20775 21097
rect 20898 21088 20904 21100
rect 20956 21088 20962 21140
rect 21174 21128 21180 21140
rect 21135 21100 21180 21128
rect 21174 21088 21180 21100
rect 21232 21088 21238 21140
rect 24581 21131 24639 21137
rect 24581 21097 24593 21131
rect 24627 21128 24639 21131
rect 24762 21128 24768 21140
rect 24627 21100 24768 21128
rect 24627 21097 24639 21100
rect 24581 21091 24639 21097
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 8395 21032 11192 21060
rect 1486 20952 1492 21004
rect 1544 20992 1550 21004
rect 2317 20995 2375 21001
rect 2317 20992 2329 20995
rect 1544 20964 2329 20992
rect 1544 20952 1550 20964
rect 2317 20961 2329 20964
rect 2363 20961 2375 20995
rect 2774 20992 2780 21004
rect 2317 20955 2375 20961
rect 2608 20964 2780 20992
rect 2332 20856 2360 20955
rect 2608 20933 2636 20964
rect 2774 20952 2780 20964
rect 2832 20992 2838 21004
rect 2961 20995 3019 21001
rect 2961 20992 2973 20995
rect 2832 20964 2973 20992
rect 2832 20952 2838 20964
rect 2961 20961 2973 20964
rect 3007 20961 3019 20995
rect 2961 20955 3019 20961
rect 4154 20952 4160 21004
rect 4212 20992 4218 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4212 20964 4445 20992
rect 4212 20952 4218 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 5994 20992 6000 21004
rect 4433 20955 4491 20961
rect 5552 20964 6000 20992
rect 2593 20927 2651 20933
rect 2593 20893 2605 20927
rect 2639 20893 2651 20927
rect 2593 20887 2651 20893
rect 3881 20927 3939 20933
rect 3881 20893 3893 20927
rect 3927 20924 3939 20927
rect 4709 20927 4767 20933
rect 4709 20924 4721 20927
rect 3927 20896 4721 20924
rect 3927 20893 3939 20896
rect 3881 20887 3939 20893
rect 4709 20893 4721 20896
rect 4755 20924 4767 20927
rect 5442 20924 5448 20936
rect 4755 20896 5448 20924
rect 4755 20893 4767 20896
rect 4709 20887 4767 20893
rect 5442 20884 5448 20896
rect 5500 20884 5506 20936
rect 2866 20856 2872 20868
rect 2332 20828 2872 20856
rect 2866 20816 2872 20828
rect 2924 20816 2930 20868
rect 3142 20816 3148 20868
rect 3200 20856 3206 20868
rect 5552 20856 5580 20964
rect 5994 20952 6000 20964
rect 6052 20952 6058 21004
rect 7561 20995 7619 21001
rect 7561 20961 7573 20995
rect 7607 20992 7619 20995
rect 7926 20992 7932 21004
rect 7607 20964 7932 20992
rect 7607 20961 7619 20964
rect 7561 20955 7619 20961
rect 7926 20952 7932 20964
rect 7984 20952 7990 21004
rect 9674 20952 9680 21004
rect 9732 20992 9738 21004
rect 9769 20995 9827 21001
rect 9769 20992 9781 20995
rect 9732 20964 9781 20992
rect 9732 20952 9738 20964
rect 9769 20961 9781 20964
rect 9815 20961 9827 20995
rect 9769 20955 9827 20961
rect 9858 20952 9864 21004
rect 9916 20992 9922 21004
rect 10025 20995 10083 21001
rect 10025 20992 10037 20995
rect 9916 20964 10037 20992
rect 9916 20952 9922 20964
rect 10025 20961 10037 20964
rect 10071 20961 10083 20995
rect 10025 20955 10083 20961
rect 6086 20924 6092 20936
rect 6047 20896 6092 20924
rect 6086 20884 6092 20896
rect 6144 20884 6150 20936
rect 6273 20927 6331 20933
rect 6273 20893 6285 20927
rect 6319 20924 6331 20927
rect 6454 20924 6460 20936
rect 6319 20896 6460 20924
rect 6319 20893 6331 20896
rect 6273 20887 6331 20893
rect 6454 20884 6460 20896
rect 6512 20884 6518 20936
rect 7745 20927 7803 20933
rect 7745 20893 7757 20927
rect 7791 20893 7803 20927
rect 7745 20887 7803 20893
rect 11164 20924 11192 21032
rect 11422 21020 11428 21072
rect 11480 21060 11486 21072
rect 13446 21060 13452 21072
rect 11480 21032 13452 21060
rect 11480 21020 11486 21032
rect 13446 21020 13452 21032
rect 13504 21020 13510 21072
rect 15102 21060 15108 21072
rect 15063 21032 15108 21060
rect 15102 21020 15108 21032
rect 15160 21020 15166 21072
rect 16485 21063 16543 21069
rect 16485 21029 16497 21063
rect 16531 21060 16543 21063
rect 16942 21060 16948 21072
rect 16531 21032 16948 21060
rect 16531 21029 16543 21032
rect 16485 21023 16543 21029
rect 16942 21020 16948 21032
rect 17000 21020 17006 21072
rect 18138 21060 18144 21072
rect 18099 21032 18144 21060
rect 18138 21020 18144 21032
rect 18196 21020 18202 21072
rect 18690 21020 18696 21072
rect 18748 21060 18754 21072
rect 19061 21063 19119 21069
rect 19061 21060 19073 21063
rect 18748 21032 19073 21060
rect 18748 21020 18754 21032
rect 19061 21029 19073 21032
rect 19107 21029 19119 21063
rect 19061 21023 19119 21029
rect 20806 21020 20812 21072
rect 20864 21060 20870 21072
rect 21542 21060 21548 21072
rect 20864 21032 21548 21060
rect 20864 21020 20870 21032
rect 21542 21020 21548 21032
rect 21600 21020 21606 21072
rect 22922 21020 22928 21072
rect 22980 21060 22986 21072
rect 24670 21060 24676 21072
rect 22980 21032 24676 21060
rect 22980 21020 22986 21032
rect 24670 21020 24676 21032
rect 24728 21020 24734 21072
rect 12161 20995 12219 21001
rect 12161 20961 12173 20995
rect 12207 20992 12219 20995
rect 12618 20992 12624 21004
rect 12207 20964 12624 20992
rect 12207 20961 12219 20964
rect 12161 20955 12219 20961
rect 12618 20952 12624 20964
rect 12676 20952 12682 21004
rect 12710 20952 12716 21004
rect 12768 20992 12774 21004
rect 14093 20995 14151 21001
rect 12768 20964 12813 20992
rect 12768 20952 12774 20964
rect 14093 20961 14105 20995
rect 14139 20992 14151 20995
rect 14274 20992 14280 21004
rect 14139 20964 14280 20992
rect 14139 20961 14151 20964
rect 14093 20955 14151 20961
rect 14274 20952 14280 20964
rect 14332 20952 14338 21004
rect 15286 20952 15292 21004
rect 15344 20992 15350 21004
rect 15657 20995 15715 21001
rect 15657 20992 15669 20995
rect 15344 20964 15669 20992
rect 15344 20952 15350 20964
rect 15657 20961 15669 20964
rect 15703 20961 15715 20995
rect 18506 20992 18512 21004
rect 15657 20955 15715 20961
rect 18340 20964 18512 20992
rect 12894 20924 12900 20936
rect 11164 20896 12900 20924
rect 3200 20828 5580 20856
rect 3200 20816 3206 20828
rect 7282 20816 7288 20868
rect 7340 20856 7346 20868
rect 7760 20856 7788 20887
rect 7340 20828 7788 20856
rect 7340 20816 7346 20828
rect 8478 20816 8484 20868
rect 8536 20856 8542 20868
rect 8665 20859 8723 20865
rect 8665 20856 8677 20859
rect 8536 20828 8677 20856
rect 8536 20816 8542 20828
rect 8665 20825 8677 20828
rect 8711 20856 8723 20859
rect 9582 20856 9588 20868
rect 8711 20828 9588 20856
rect 8711 20825 8723 20828
rect 8665 20819 8723 20825
rect 9582 20816 9588 20828
rect 9640 20816 9646 20868
rect 11164 20865 11192 20896
rect 12894 20884 12900 20896
rect 12952 20884 12958 20936
rect 15838 20924 15844 20936
rect 15799 20896 15844 20924
rect 15838 20884 15844 20896
rect 15896 20884 15902 20936
rect 17862 20884 17868 20936
rect 17920 20924 17926 20936
rect 18340 20933 18368 20964
rect 18506 20952 18512 20964
rect 18564 20992 18570 21004
rect 18785 20995 18843 21001
rect 18785 20992 18797 20995
rect 18564 20964 18797 20992
rect 18564 20952 18570 20964
rect 18785 20961 18797 20964
rect 18831 20961 18843 20995
rect 18785 20955 18843 20961
rect 19613 20995 19671 21001
rect 19613 20961 19625 20995
rect 19659 20992 19671 20995
rect 19978 20992 19984 21004
rect 19659 20964 19984 20992
rect 19659 20961 19671 20964
rect 19613 20955 19671 20961
rect 19978 20952 19984 20964
rect 20036 20952 20042 21004
rect 21450 20952 21456 21004
rect 21508 20992 21514 21004
rect 21985 20995 22043 21001
rect 21985 20992 21997 20995
rect 21508 20964 21997 20992
rect 21508 20952 21514 20964
rect 21985 20961 21997 20964
rect 22031 20961 22043 20995
rect 21985 20955 22043 20961
rect 23934 20952 23940 21004
rect 23992 20992 23998 21004
rect 25225 20995 25283 21001
rect 25225 20992 25237 20995
rect 23992 20964 25237 20992
rect 23992 20952 23998 20964
rect 25225 20961 25237 20964
rect 25271 20961 25283 20995
rect 25225 20955 25283 20961
rect 18325 20927 18383 20933
rect 18325 20924 18337 20927
rect 17920 20896 18337 20924
rect 17920 20884 17926 20896
rect 18325 20893 18337 20896
rect 18371 20893 18383 20927
rect 18325 20887 18383 20893
rect 19150 20884 19156 20936
rect 19208 20924 19214 20936
rect 19705 20927 19763 20933
rect 19705 20924 19717 20927
rect 19208 20896 19717 20924
rect 19208 20884 19214 20896
rect 19705 20893 19717 20896
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 19797 20927 19855 20933
rect 19797 20893 19809 20927
rect 19843 20893 19855 20927
rect 19797 20887 19855 20893
rect 11149 20859 11207 20865
rect 11149 20825 11161 20859
rect 11195 20825 11207 20859
rect 11149 20819 11207 20825
rect 12066 20816 12072 20868
rect 12124 20856 12130 20868
rect 12250 20856 12256 20868
rect 12124 20828 12256 20856
rect 12124 20816 12130 20828
rect 12250 20816 12256 20828
rect 12308 20816 12314 20868
rect 14458 20816 14464 20868
rect 14516 20856 14522 20868
rect 14737 20859 14795 20865
rect 14737 20856 14749 20859
rect 14516 20828 14749 20856
rect 14516 20816 14522 20828
rect 14737 20825 14749 20828
rect 14783 20856 14795 20859
rect 15289 20859 15347 20865
rect 15289 20856 15301 20859
rect 14783 20828 15301 20856
rect 14783 20825 14795 20828
rect 14737 20819 14795 20825
rect 15289 20825 15301 20828
rect 15335 20825 15347 20859
rect 15289 20819 15347 20825
rect 17221 20859 17279 20865
rect 17221 20825 17233 20859
rect 17267 20856 17279 20859
rect 17681 20859 17739 20865
rect 17681 20856 17693 20859
rect 17267 20828 17693 20856
rect 17267 20825 17279 20828
rect 17221 20819 17279 20825
rect 17681 20825 17693 20828
rect 17727 20856 17739 20859
rect 17770 20856 17776 20868
rect 17727 20828 17776 20856
rect 17727 20825 17739 20828
rect 17681 20819 17739 20825
rect 17770 20816 17776 20828
rect 17828 20816 17834 20868
rect 18506 20816 18512 20868
rect 18564 20856 18570 20868
rect 19242 20856 19248 20868
rect 18564 20828 19248 20856
rect 18564 20816 18570 20828
rect 19242 20816 19248 20828
rect 19300 20856 19306 20868
rect 19812 20856 19840 20887
rect 20254 20884 20260 20936
rect 20312 20924 20318 20936
rect 20622 20924 20628 20936
rect 20312 20896 20628 20924
rect 20312 20884 20318 20896
rect 20622 20884 20628 20896
rect 20680 20884 20686 20936
rect 20898 20884 20904 20936
rect 20956 20924 20962 20936
rect 21729 20927 21787 20933
rect 21729 20924 21741 20927
rect 20956 20896 21741 20924
rect 20956 20884 20962 20896
rect 21729 20893 21741 20896
rect 21775 20893 21787 20927
rect 24765 20927 24823 20933
rect 24765 20924 24777 20927
rect 21729 20887 21787 20893
rect 23676 20896 24777 20924
rect 19300 20828 19840 20856
rect 19300 20816 19306 20828
rect 23676 20800 23704 20896
rect 24765 20893 24777 20896
rect 24811 20893 24823 20927
rect 24765 20887 24823 20893
rect 24394 20816 24400 20868
rect 24452 20856 24458 20868
rect 24452 20828 24808 20856
rect 24452 20816 24458 20828
rect 24780 20800 24808 20828
rect 3510 20788 3516 20800
rect 3471 20760 3516 20788
rect 3510 20748 3516 20760
rect 3568 20748 3574 20800
rect 4982 20748 4988 20800
rect 5040 20788 5046 20800
rect 5077 20791 5135 20797
rect 5077 20788 5089 20791
rect 5040 20760 5089 20788
rect 5040 20748 5046 20760
rect 5077 20757 5089 20760
rect 5123 20757 5135 20791
rect 6730 20788 6736 20800
rect 6691 20760 6736 20788
rect 5077 20751 5135 20757
rect 6730 20748 6736 20760
rect 6788 20748 6794 20800
rect 6914 20748 6920 20800
rect 6972 20788 6978 20800
rect 7193 20791 7251 20797
rect 7193 20788 7205 20791
rect 6972 20760 7205 20788
rect 6972 20748 6978 20760
rect 7193 20757 7205 20760
rect 7239 20757 7251 20791
rect 9398 20788 9404 20800
rect 9359 20760 9404 20788
rect 7193 20751 7251 20757
rect 9398 20748 9404 20760
rect 9456 20748 9462 20800
rect 13998 20788 14004 20800
rect 13959 20760 14004 20788
rect 13998 20748 14004 20760
rect 14056 20748 14062 20800
rect 21358 20748 21364 20800
rect 21416 20788 21422 20800
rect 21910 20788 21916 20800
rect 21416 20760 21916 20788
rect 21416 20748 21422 20760
rect 21910 20748 21916 20760
rect 21968 20748 21974 20800
rect 22462 20748 22468 20800
rect 22520 20788 22526 20800
rect 23109 20791 23167 20797
rect 23109 20788 23121 20791
rect 22520 20760 23121 20788
rect 22520 20748 22526 20760
rect 23109 20757 23121 20760
rect 23155 20788 23167 20791
rect 23658 20788 23664 20800
rect 23155 20760 23664 20788
rect 23155 20757 23167 20760
rect 23109 20751 23167 20757
rect 23658 20748 23664 20760
rect 23716 20748 23722 20800
rect 24026 20788 24032 20800
rect 23987 20760 24032 20788
rect 24026 20748 24032 20760
rect 24084 20748 24090 20800
rect 24118 20748 24124 20800
rect 24176 20788 24182 20800
rect 24213 20791 24271 20797
rect 24213 20788 24225 20791
rect 24176 20760 24225 20788
rect 24176 20748 24182 20760
rect 24213 20757 24225 20760
rect 24259 20757 24271 20791
rect 24213 20751 24271 20757
rect 24762 20748 24768 20800
rect 24820 20748 24826 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1210 20544 1216 20596
rect 1268 20584 1274 20596
rect 1765 20587 1823 20593
rect 1765 20584 1777 20587
rect 1268 20556 1777 20584
rect 1268 20544 1274 20556
rect 1765 20553 1777 20556
rect 1811 20553 1823 20587
rect 1765 20547 1823 20553
rect 1949 20587 2007 20593
rect 1949 20553 1961 20587
rect 1995 20584 2007 20587
rect 2130 20584 2136 20596
rect 1995 20556 2136 20584
rect 1995 20553 2007 20556
rect 1949 20547 2007 20553
rect 1780 20448 1808 20547
rect 2130 20544 2136 20556
rect 2188 20544 2194 20596
rect 3053 20587 3111 20593
rect 3053 20553 3065 20587
rect 3099 20584 3111 20587
rect 3142 20584 3148 20596
rect 3099 20556 3148 20584
rect 3099 20553 3111 20556
rect 3053 20547 3111 20553
rect 3142 20544 3148 20556
rect 3200 20544 3206 20596
rect 5994 20544 6000 20596
rect 6052 20584 6058 20596
rect 6181 20587 6239 20593
rect 6181 20584 6193 20587
rect 6052 20556 6193 20584
rect 6052 20544 6058 20556
rect 6181 20553 6193 20556
rect 6227 20553 6239 20587
rect 6181 20547 6239 20553
rect 6454 20544 6460 20596
rect 6512 20584 6518 20596
rect 6549 20587 6607 20593
rect 6549 20584 6561 20587
rect 6512 20556 6561 20584
rect 6512 20544 6518 20556
rect 6549 20553 6561 20556
rect 6595 20553 6607 20587
rect 6549 20547 6607 20553
rect 2866 20476 2872 20528
rect 2924 20516 2930 20528
rect 3329 20519 3387 20525
rect 3329 20516 3341 20519
rect 2924 20488 3341 20516
rect 2924 20476 2930 20488
rect 3329 20485 3341 20488
rect 3375 20516 3387 20519
rect 3694 20516 3700 20528
rect 3375 20488 3700 20516
rect 3375 20485 3387 20488
rect 3329 20479 3387 20485
rect 3694 20476 3700 20488
rect 3752 20476 3758 20528
rect 2406 20448 2412 20460
rect 1780 20420 2412 20448
rect 2406 20408 2412 20420
rect 2464 20408 2470 20460
rect 2498 20408 2504 20460
rect 2556 20448 2562 20460
rect 2593 20451 2651 20457
rect 2593 20448 2605 20451
rect 2556 20420 2605 20448
rect 2556 20408 2562 20420
rect 2593 20417 2605 20420
rect 2639 20448 2651 20451
rect 2774 20448 2780 20460
rect 2639 20420 2780 20448
rect 2639 20417 2651 20420
rect 2593 20411 2651 20417
rect 2774 20408 2780 20420
rect 2832 20408 2838 20460
rect 5258 20408 5264 20460
rect 5316 20448 5322 20460
rect 5994 20448 6000 20460
rect 5316 20420 6000 20448
rect 5316 20408 5322 20420
rect 5994 20408 6000 20420
rect 6052 20408 6058 20460
rect 6564 20448 6592 20547
rect 6822 20544 6828 20596
rect 6880 20584 6886 20596
rect 6880 20556 8708 20584
rect 6880 20544 6886 20556
rect 8680 20516 8708 20556
rect 9582 20544 9588 20596
rect 9640 20584 9646 20596
rect 10229 20587 10287 20593
rect 10229 20584 10241 20587
rect 9640 20556 10241 20584
rect 9640 20544 9646 20556
rect 10229 20553 10241 20556
rect 10275 20553 10287 20587
rect 10229 20547 10287 20553
rect 12437 20587 12495 20593
rect 12437 20553 12449 20587
rect 12483 20584 12495 20587
rect 12618 20584 12624 20596
rect 12483 20556 12624 20584
rect 12483 20553 12495 20556
rect 12437 20547 12495 20553
rect 12618 20544 12624 20556
rect 12676 20544 12682 20596
rect 12894 20544 12900 20596
rect 12952 20584 12958 20596
rect 13449 20587 13507 20593
rect 13449 20584 13461 20587
rect 12952 20556 13461 20584
rect 12952 20544 12958 20556
rect 13449 20553 13461 20556
rect 13495 20553 13507 20587
rect 13449 20547 13507 20553
rect 14001 20587 14059 20593
rect 14001 20553 14013 20587
rect 14047 20584 14059 20587
rect 14090 20584 14096 20596
rect 14047 20556 14096 20584
rect 14047 20553 14059 20556
rect 14001 20547 14059 20553
rect 14090 20544 14096 20556
rect 14148 20544 14154 20596
rect 15746 20584 15752 20596
rect 15707 20556 15752 20584
rect 15746 20544 15752 20556
rect 15804 20544 15810 20596
rect 17773 20587 17831 20593
rect 17773 20553 17785 20587
rect 17819 20584 17831 20587
rect 17862 20584 17868 20596
rect 17819 20556 17868 20584
rect 17819 20553 17831 20556
rect 17773 20547 17831 20553
rect 17862 20544 17868 20556
rect 17920 20544 17926 20596
rect 18506 20584 18512 20596
rect 18467 20556 18512 20584
rect 18506 20544 18512 20556
rect 18564 20544 18570 20596
rect 21085 20587 21143 20593
rect 21085 20553 21097 20587
rect 21131 20584 21143 20587
rect 21450 20584 21456 20596
rect 21131 20556 21456 20584
rect 21131 20553 21143 20556
rect 21085 20547 21143 20553
rect 21450 20544 21456 20556
rect 21508 20584 21514 20596
rect 22186 20584 22192 20596
rect 21508 20556 22192 20584
rect 21508 20544 21514 20556
rect 22186 20544 22192 20556
rect 22244 20544 22250 20596
rect 22646 20544 22652 20596
rect 22704 20584 22710 20596
rect 22922 20584 22928 20596
rect 22704 20556 22928 20584
rect 22704 20544 22710 20556
rect 22922 20544 22928 20556
rect 22980 20544 22986 20596
rect 12069 20519 12127 20525
rect 12069 20516 12081 20519
rect 8680 20488 12081 20516
rect 12069 20485 12081 20488
rect 12115 20516 12127 20519
rect 12161 20519 12219 20525
rect 12161 20516 12173 20519
rect 12115 20488 12173 20516
rect 12115 20485 12127 20488
rect 12069 20479 12127 20485
rect 12161 20485 12173 20488
rect 12207 20485 12219 20519
rect 12161 20479 12219 20485
rect 13909 20519 13967 20525
rect 13909 20485 13921 20519
rect 13955 20516 13967 20519
rect 16390 20516 16396 20528
rect 13955 20488 14688 20516
rect 16351 20488 16396 20516
rect 13955 20485 13967 20488
rect 13909 20479 13967 20485
rect 14660 20460 14688 20488
rect 16390 20476 16396 20488
rect 16448 20476 16454 20528
rect 7098 20448 7104 20460
rect 6564 20420 7104 20448
rect 7098 20408 7104 20420
rect 7156 20448 7162 20460
rect 7156 20420 7880 20448
rect 7156 20408 7162 20420
rect 7852 20392 7880 20420
rect 9858 20408 9864 20460
rect 9916 20448 9922 20460
rect 10781 20451 10839 20457
rect 10781 20448 10793 20451
rect 9916 20420 10793 20448
rect 9916 20408 9922 20420
rect 10781 20417 10793 20420
rect 10827 20448 10839 20451
rect 11241 20451 11299 20457
rect 11241 20448 11253 20451
rect 10827 20420 11253 20448
rect 10827 20417 10839 20420
rect 10781 20411 10839 20417
rect 11241 20417 11253 20420
rect 11287 20448 11299 20451
rect 11793 20451 11851 20457
rect 11793 20448 11805 20451
rect 11287 20420 11805 20448
rect 11287 20417 11299 20420
rect 11241 20411 11299 20417
rect 11793 20417 11805 20420
rect 11839 20448 11851 20451
rect 12989 20451 13047 20457
rect 12989 20448 13001 20451
rect 11839 20420 13001 20448
rect 11839 20417 11851 20420
rect 11793 20411 11851 20417
rect 12989 20417 13001 20420
rect 13035 20417 13047 20451
rect 14458 20448 14464 20460
rect 14419 20420 14464 20448
rect 12989 20411 13047 20417
rect 14458 20408 14464 20420
rect 14516 20408 14522 20460
rect 14642 20448 14648 20460
rect 14603 20420 14648 20448
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 16942 20448 16948 20460
rect 16903 20420 16948 20448
rect 16942 20408 16948 20420
rect 17000 20408 17006 20460
rect 18598 20408 18604 20460
rect 18656 20448 18662 20460
rect 18969 20451 19027 20457
rect 18969 20448 18981 20451
rect 18656 20420 18981 20448
rect 18656 20408 18662 20420
rect 18969 20417 18981 20420
rect 19015 20448 19027 20451
rect 19061 20451 19119 20457
rect 19061 20448 19073 20451
rect 19015 20420 19073 20448
rect 19015 20417 19027 20420
rect 18969 20411 19027 20417
rect 19061 20417 19073 20420
rect 19107 20417 19119 20451
rect 19061 20411 19119 20417
rect 21542 20408 21548 20460
rect 21600 20448 21606 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21600 20420 22017 20448
rect 21600 20408 21606 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22189 20451 22247 20457
rect 22189 20417 22201 20451
rect 22235 20448 22247 20451
rect 22370 20448 22376 20460
rect 22235 20420 22376 20448
rect 22235 20417 22247 20420
rect 22189 20411 22247 20417
rect 22370 20408 22376 20420
rect 22428 20448 22434 20460
rect 22925 20451 22983 20457
rect 22925 20448 22937 20451
rect 22428 20420 22937 20448
rect 22428 20408 22434 20420
rect 22925 20417 22937 20420
rect 22971 20417 22983 20451
rect 22925 20411 22983 20417
rect 3326 20340 3332 20392
rect 3384 20380 3390 20392
rect 3697 20383 3755 20389
rect 3697 20380 3709 20383
rect 3384 20352 3709 20380
rect 3384 20340 3390 20352
rect 3697 20349 3709 20352
rect 3743 20349 3755 20383
rect 3697 20343 3755 20349
rect 3881 20383 3939 20389
rect 3881 20349 3893 20383
rect 3927 20380 3939 20383
rect 4706 20380 4712 20392
rect 3927 20352 4712 20380
rect 3927 20349 3939 20352
rect 3881 20343 3939 20349
rect 4706 20340 4712 20352
rect 4764 20340 4770 20392
rect 5810 20380 5816 20392
rect 5771 20352 5816 20380
rect 5810 20340 5816 20352
rect 5868 20380 5874 20392
rect 6086 20380 6092 20392
rect 5868 20352 6092 20380
rect 5868 20340 5874 20352
rect 6086 20340 6092 20352
rect 6144 20340 6150 20392
rect 7745 20383 7803 20389
rect 7745 20349 7757 20383
rect 7791 20349 7803 20383
rect 7745 20343 7803 20349
rect 3510 20272 3516 20324
rect 3568 20312 3574 20324
rect 4126 20315 4184 20321
rect 4126 20312 4138 20315
rect 3568 20284 4138 20312
rect 3568 20272 3574 20284
rect 4126 20281 4138 20284
rect 4172 20312 4184 20315
rect 4982 20312 4988 20324
rect 4172 20284 4988 20312
rect 4172 20281 4184 20284
rect 4126 20275 4184 20281
rect 4982 20272 4988 20284
rect 5040 20272 5046 20324
rect 7558 20272 7564 20324
rect 7616 20312 7622 20324
rect 7653 20315 7711 20321
rect 7653 20312 7665 20315
rect 7616 20284 7665 20312
rect 7616 20272 7622 20284
rect 7653 20281 7665 20284
rect 7699 20312 7711 20315
rect 7760 20312 7788 20343
rect 7834 20340 7840 20392
rect 7892 20380 7898 20392
rect 8001 20383 8059 20389
rect 8001 20380 8013 20383
rect 7892 20352 8013 20380
rect 7892 20340 7898 20352
rect 8001 20349 8013 20352
rect 8047 20349 8059 20383
rect 8001 20343 8059 20349
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 10689 20383 10747 20389
rect 10689 20380 10701 20383
rect 9732 20352 9777 20380
rect 10060 20352 10701 20380
rect 9732 20340 9738 20352
rect 9692 20312 9720 20340
rect 7699 20284 9720 20312
rect 7699 20281 7711 20284
rect 7653 20275 7711 20281
rect 10060 20256 10088 20352
rect 10689 20349 10701 20352
rect 10735 20380 10747 20383
rect 11606 20380 11612 20392
rect 10735 20352 11612 20380
rect 10735 20349 10747 20352
rect 10689 20343 10747 20349
rect 11606 20340 11612 20352
rect 11664 20340 11670 20392
rect 13814 20380 13820 20392
rect 11900 20352 13820 20380
rect 10597 20315 10655 20321
rect 10597 20281 10609 20315
rect 10643 20312 10655 20315
rect 10778 20312 10784 20324
rect 10643 20284 10784 20312
rect 10643 20281 10655 20284
rect 10597 20275 10655 20281
rect 10778 20272 10784 20284
rect 10836 20312 10842 20324
rect 11900 20312 11928 20352
rect 13814 20340 13820 20352
rect 13872 20340 13878 20392
rect 19334 20389 19340 20392
rect 19328 20380 19340 20389
rect 19295 20352 19340 20380
rect 19328 20343 19340 20352
rect 19334 20340 19340 20343
rect 19392 20340 19398 20392
rect 22649 20383 22707 20389
rect 22649 20349 22661 20383
rect 22695 20380 22707 20383
rect 23014 20380 23020 20392
rect 22695 20352 23020 20380
rect 22695 20349 22707 20352
rect 22649 20343 22707 20349
rect 23014 20340 23020 20352
rect 23072 20380 23078 20392
rect 23477 20383 23535 20389
rect 23477 20380 23489 20383
rect 23072 20352 23489 20380
rect 23072 20340 23078 20352
rect 23477 20349 23489 20352
rect 23523 20380 23535 20383
rect 23661 20383 23719 20389
rect 23661 20380 23673 20383
rect 23523 20352 23673 20380
rect 23523 20349 23535 20352
rect 23477 20343 23535 20349
rect 23661 20349 23673 20352
rect 23707 20349 23719 20383
rect 25958 20380 25964 20392
rect 25919 20352 25964 20380
rect 23661 20343 23719 20349
rect 25958 20340 25964 20352
rect 26016 20340 26022 20392
rect 10836 20284 11928 20312
rect 10836 20272 10842 20284
rect 11974 20272 11980 20324
rect 12032 20312 12038 20324
rect 12069 20315 12127 20321
rect 12069 20312 12081 20315
rect 12032 20284 12081 20312
rect 12032 20272 12038 20284
rect 12069 20281 12081 20284
rect 12115 20312 12127 20315
rect 12805 20315 12863 20321
rect 12805 20312 12817 20315
rect 12115 20284 12817 20312
rect 12115 20281 12127 20284
rect 12069 20275 12127 20281
rect 12805 20281 12817 20284
rect 12851 20281 12863 20315
rect 12805 20275 12863 20281
rect 13722 20272 13728 20324
rect 13780 20312 13786 20324
rect 14734 20312 14740 20324
rect 13780 20284 14740 20312
rect 13780 20272 13786 20284
rect 14734 20272 14740 20284
rect 14792 20312 14798 20324
rect 15289 20315 15347 20321
rect 15289 20312 15301 20315
rect 14792 20284 15301 20312
rect 14792 20272 14798 20284
rect 15289 20281 15301 20284
rect 15335 20281 15347 20315
rect 15289 20275 15347 20281
rect 16482 20272 16488 20324
rect 16540 20312 16546 20324
rect 16761 20315 16819 20321
rect 16761 20312 16773 20315
rect 16540 20284 16773 20312
rect 16540 20272 16546 20284
rect 16761 20281 16773 20284
rect 16807 20312 16819 20315
rect 18049 20315 18107 20321
rect 18049 20312 18061 20315
rect 16807 20284 18061 20312
rect 16807 20281 16819 20284
rect 16761 20275 16819 20281
rect 18049 20281 18061 20284
rect 18095 20281 18107 20315
rect 18049 20275 18107 20281
rect 20714 20272 20720 20324
rect 20772 20312 20778 20324
rect 21453 20315 21511 20321
rect 21453 20312 21465 20315
rect 20772 20284 21465 20312
rect 20772 20272 20778 20284
rect 21453 20281 21465 20284
rect 21499 20312 21511 20315
rect 21913 20315 21971 20321
rect 21913 20312 21925 20315
rect 21499 20284 21925 20312
rect 21499 20281 21511 20284
rect 21453 20275 21511 20281
rect 21913 20281 21925 20284
rect 21959 20281 21971 20315
rect 23906 20315 23964 20321
rect 23906 20312 23918 20315
rect 21913 20275 21971 20281
rect 23676 20284 23918 20312
rect 23676 20256 23704 20284
rect 23906 20281 23918 20284
rect 23952 20312 23964 20315
rect 25593 20315 25651 20321
rect 25593 20312 25605 20315
rect 23952 20284 25605 20312
rect 23952 20281 23964 20284
rect 23906 20275 23964 20281
rect 25593 20281 25605 20284
rect 25639 20281 25651 20315
rect 25593 20275 25651 20281
rect 2314 20244 2320 20256
rect 2227 20216 2320 20244
rect 2314 20204 2320 20216
rect 2372 20244 2378 20256
rect 4338 20244 4344 20256
rect 2372 20216 4344 20244
rect 2372 20204 2378 20216
rect 4338 20204 4344 20216
rect 4396 20204 4402 20256
rect 5258 20244 5264 20256
rect 5219 20216 5264 20244
rect 5258 20204 5264 20216
rect 5316 20204 5322 20256
rect 7190 20244 7196 20256
rect 7151 20216 7196 20244
rect 7190 20204 7196 20216
rect 7248 20204 7254 20256
rect 8754 20204 8760 20256
rect 8812 20244 8818 20256
rect 9125 20247 9183 20253
rect 9125 20244 9137 20247
rect 8812 20216 9137 20244
rect 8812 20204 8818 20216
rect 9125 20213 9137 20216
rect 9171 20213 9183 20247
rect 10042 20244 10048 20256
rect 10003 20216 10048 20244
rect 9125 20207 9183 20213
rect 10042 20204 10048 20216
rect 10100 20204 10106 20256
rect 12894 20244 12900 20256
rect 12855 20216 12900 20244
rect 12894 20204 12900 20216
rect 12952 20204 12958 20256
rect 14274 20204 14280 20256
rect 14332 20244 14338 20256
rect 14369 20247 14427 20253
rect 14369 20244 14381 20247
rect 14332 20216 14381 20244
rect 14332 20204 14338 20216
rect 14369 20213 14381 20216
rect 14415 20213 14427 20247
rect 16206 20244 16212 20256
rect 16167 20216 16212 20244
rect 14369 20207 14427 20213
rect 16206 20204 16212 20216
rect 16264 20244 16270 20256
rect 16853 20247 16911 20253
rect 16853 20244 16865 20247
rect 16264 20216 16865 20244
rect 16264 20204 16270 20216
rect 16853 20213 16865 20216
rect 16899 20244 16911 20247
rect 17310 20244 17316 20256
rect 16899 20216 17316 20244
rect 16899 20213 16911 20216
rect 16853 20207 16911 20213
rect 17310 20204 17316 20216
rect 17368 20204 17374 20256
rect 18322 20204 18328 20256
rect 18380 20244 18386 20256
rect 19334 20244 19340 20256
rect 18380 20216 19340 20244
rect 18380 20204 18386 20216
rect 19334 20204 19340 20216
rect 19392 20204 19398 20256
rect 20438 20244 20444 20256
rect 20399 20216 20444 20244
rect 20438 20204 20444 20216
rect 20496 20204 20502 20256
rect 21542 20244 21548 20256
rect 21503 20216 21548 20244
rect 21542 20204 21548 20216
rect 21600 20204 21606 20256
rect 23658 20204 23664 20256
rect 23716 20204 23722 20256
rect 24026 20204 24032 20256
rect 24084 20244 24090 20256
rect 25041 20247 25099 20253
rect 25041 20244 25053 20247
rect 24084 20216 25053 20244
rect 24084 20204 24090 20216
rect 25041 20213 25053 20216
rect 25087 20213 25099 20247
rect 25041 20207 25099 20213
rect 25774 20204 25780 20256
rect 25832 20244 25838 20256
rect 25958 20244 25964 20256
rect 25832 20216 25964 20244
rect 25832 20204 25838 20216
rect 25958 20204 25964 20216
rect 26016 20204 26022 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 934 20000 940 20052
rect 992 20040 998 20052
rect 2041 20043 2099 20049
rect 2041 20040 2053 20043
rect 992 20012 2053 20040
rect 992 20000 998 20012
rect 2041 20009 2053 20012
rect 2087 20040 2099 20043
rect 2314 20040 2320 20052
rect 2087 20012 2320 20040
rect 2087 20009 2099 20012
rect 2041 20003 2099 20009
rect 2314 20000 2320 20012
rect 2372 20000 2378 20052
rect 4982 20000 4988 20052
rect 5040 20040 5046 20052
rect 6825 20043 6883 20049
rect 6825 20040 6837 20043
rect 5040 20012 6837 20040
rect 5040 20000 5046 20012
rect 6825 20009 6837 20012
rect 6871 20040 6883 20043
rect 7190 20040 7196 20052
rect 6871 20012 7196 20040
rect 6871 20009 6883 20012
rect 6825 20003 6883 20009
rect 7190 20000 7196 20012
rect 7248 20000 7254 20052
rect 7834 20040 7840 20052
rect 7795 20012 7840 20040
rect 7834 20000 7840 20012
rect 7892 20000 7898 20052
rect 8294 20040 8300 20052
rect 8255 20012 8300 20040
rect 8294 20000 8300 20012
rect 8352 20000 8358 20052
rect 9674 20040 9680 20052
rect 9635 20012 9680 20040
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 10134 20000 10140 20052
rect 10192 20040 10198 20052
rect 10321 20043 10379 20049
rect 10321 20040 10333 20043
rect 10192 20012 10333 20040
rect 10192 20000 10198 20012
rect 10321 20009 10333 20012
rect 10367 20040 10379 20043
rect 10778 20040 10784 20052
rect 10367 20012 10784 20040
rect 10367 20009 10379 20012
rect 10321 20003 10379 20009
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 11054 20000 11060 20052
rect 11112 20000 11118 20052
rect 11149 20043 11207 20049
rect 11149 20009 11161 20043
rect 11195 20040 11207 20043
rect 11514 20040 11520 20052
rect 11195 20012 11520 20040
rect 11195 20009 11207 20012
rect 11149 20003 11207 20009
rect 11514 20000 11520 20012
rect 11572 20000 11578 20052
rect 12529 20043 12587 20049
rect 12529 20009 12541 20043
rect 12575 20040 12587 20043
rect 12894 20040 12900 20052
rect 12575 20012 12900 20040
rect 12575 20009 12587 20012
rect 12529 20003 12587 20009
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 15102 20040 15108 20052
rect 15063 20012 15108 20040
rect 15102 20000 15108 20012
rect 15160 20000 15166 20052
rect 15654 20000 15660 20052
rect 15712 20040 15718 20052
rect 15749 20043 15807 20049
rect 15749 20040 15761 20043
rect 15712 20012 15761 20040
rect 15712 20000 15718 20012
rect 15749 20009 15761 20012
rect 15795 20009 15807 20043
rect 16482 20040 16488 20052
rect 16443 20012 16488 20040
rect 15749 20003 15807 20009
rect 16482 20000 16488 20012
rect 16540 20000 16546 20052
rect 16850 20000 16856 20052
rect 16908 20040 16914 20052
rect 17402 20040 17408 20052
rect 16908 20012 17408 20040
rect 16908 20000 16914 20012
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 18138 20040 18144 20052
rect 18099 20012 18144 20040
rect 18138 20000 18144 20012
rect 18196 20000 18202 20052
rect 18966 20000 18972 20052
rect 19024 20040 19030 20052
rect 19024 20012 19104 20040
rect 19024 20000 19030 20012
rect 2866 19972 2872 19984
rect 2827 19944 2872 19972
rect 2866 19932 2872 19944
rect 2924 19932 2930 19984
rect 3510 19972 3516 19984
rect 3471 19944 3516 19972
rect 3510 19932 3516 19944
rect 3568 19932 3574 19984
rect 3881 19975 3939 19981
rect 3881 19941 3893 19975
rect 3927 19972 3939 19975
rect 4154 19972 4160 19984
rect 3927 19944 4160 19972
rect 3927 19941 3939 19944
rect 3881 19935 3939 19941
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19904 2835 19907
rect 3786 19904 3792 19916
rect 2823 19876 3792 19904
rect 2823 19873 2835 19876
rect 2777 19867 2835 19873
rect 3786 19864 3792 19876
rect 3844 19864 3850 19916
rect 1397 19839 1455 19845
rect 1397 19805 1409 19839
rect 1443 19805 1455 19839
rect 3050 19836 3056 19848
rect 3011 19808 3056 19836
rect 1397 19799 1455 19805
rect 1412 19768 1440 19799
rect 3050 19796 3056 19808
rect 3108 19796 3114 19848
rect 3896 19768 3924 19935
rect 4154 19932 4160 19944
rect 4212 19932 4218 19984
rect 11072 19972 11100 20000
rect 12069 19975 12127 19981
rect 12069 19972 12081 19975
rect 11072 19944 12081 19972
rect 12069 19941 12081 19944
rect 12115 19941 12127 19975
rect 12069 19935 12127 19941
rect 17126 19932 17132 19984
rect 17184 19972 17190 19984
rect 17497 19975 17555 19981
rect 17497 19972 17509 19975
rect 17184 19944 17509 19972
rect 17184 19932 17190 19944
rect 17497 19941 17509 19944
rect 17543 19972 17555 19975
rect 17770 19972 17776 19984
rect 17543 19944 17776 19972
rect 17543 19941 17555 19944
rect 17497 19935 17555 19941
rect 17770 19932 17776 19944
rect 17828 19932 17834 19984
rect 19076 19981 19104 20012
rect 19426 20000 19432 20052
rect 19484 20040 19490 20052
rect 19613 20043 19671 20049
rect 19613 20040 19625 20043
rect 19484 20012 19625 20040
rect 19484 20000 19490 20012
rect 19613 20009 19625 20012
rect 19659 20009 19671 20043
rect 19613 20003 19671 20009
rect 22094 20000 22100 20052
rect 22152 20040 22158 20052
rect 23201 20043 23259 20049
rect 23201 20040 23213 20043
rect 22152 20012 23213 20040
rect 22152 20000 22158 20012
rect 23201 20009 23213 20012
rect 23247 20040 23259 20043
rect 23845 20043 23903 20049
rect 23845 20040 23857 20043
rect 23247 20012 23857 20040
rect 23247 20009 23259 20012
rect 23201 20003 23259 20009
rect 23845 20009 23857 20012
rect 23891 20009 23903 20043
rect 23845 20003 23903 20009
rect 24489 20043 24547 20049
rect 24489 20009 24501 20043
rect 24535 20040 24547 20043
rect 24670 20040 24676 20052
rect 24535 20012 24676 20040
rect 24535 20009 24547 20012
rect 24489 20003 24547 20009
rect 24670 20000 24676 20012
rect 24728 20000 24734 20052
rect 24854 20040 24860 20052
rect 24815 20012 24860 20040
rect 24854 20000 24860 20012
rect 24912 20000 24918 20052
rect 25130 20040 25136 20052
rect 25091 20012 25136 20040
rect 25130 20000 25136 20012
rect 25188 20000 25194 20052
rect 19061 19975 19119 19981
rect 19061 19941 19073 19975
rect 19107 19972 19119 19975
rect 19242 19972 19248 19984
rect 19107 19944 19248 19972
rect 19107 19941 19119 19944
rect 19061 19935 19119 19941
rect 19242 19932 19248 19944
rect 19300 19932 19306 19984
rect 21168 19975 21226 19981
rect 21168 19941 21180 19975
rect 21214 19972 21226 19975
rect 21266 19972 21272 19984
rect 21214 19944 21272 19972
rect 21214 19941 21226 19944
rect 21168 19935 21226 19941
rect 21266 19932 21272 19944
rect 21324 19932 21330 19984
rect 23106 19932 23112 19984
rect 23164 19972 23170 19984
rect 24578 19972 24584 19984
rect 23164 19944 24584 19972
rect 23164 19932 23170 19944
rect 24578 19932 24584 19944
rect 24636 19932 24642 19984
rect 4062 19904 4068 19916
rect 4023 19876 4068 19904
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 4706 19904 4712 19916
rect 4619 19876 4712 19904
rect 4706 19864 4712 19876
rect 4764 19904 4770 19916
rect 4982 19904 4988 19916
rect 4764 19876 4988 19904
rect 4764 19864 4770 19876
rect 4982 19864 4988 19876
rect 5040 19904 5046 19916
rect 5445 19907 5503 19913
rect 5445 19904 5457 19907
rect 5040 19876 5457 19904
rect 5040 19864 5046 19876
rect 5445 19873 5457 19876
rect 5491 19873 5503 19907
rect 5445 19867 5503 19873
rect 5534 19864 5540 19916
rect 5592 19904 5598 19916
rect 5712 19907 5770 19913
rect 5712 19904 5724 19907
rect 5592 19876 5724 19904
rect 5592 19864 5598 19876
rect 5712 19873 5724 19876
rect 5758 19904 5770 19907
rect 6730 19904 6736 19916
rect 5758 19876 6736 19904
rect 5758 19873 5770 19876
rect 5712 19867 5770 19873
rect 6730 19864 6736 19876
rect 6788 19864 6794 19916
rect 7469 19907 7527 19913
rect 7469 19873 7481 19907
rect 7515 19904 7527 19907
rect 8018 19904 8024 19916
rect 7515 19876 8024 19904
rect 7515 19873 7527 19876
rect 7469 19867 7527 19873
rect 8018 19864 8024 19876
rect 8076 19904 8082 19916
rect 8389 19907 8447 19913
rect 8389 19904 8401 19907
rect 8076 19876 8401 19904
rect 8076 19864 8082 19876
rect 8389 19873 8401 19876
rect 8435 19873 8447 19907
rect 8389 19867 8447 19873
rect 11057 19907 11115 19913
rect 11057 19873 11069 19907
rect 11103 19904 11115 19907
rect 11882 19904 11888 19916
rect 11103 19876 11888 19904
rect 11103 19873 11115 19876
rect 11057 19867 11115 19873
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 12802 19864 12808 19916
rect 12860 19904 12866 19916
rect 12969 19907 13027 19913
rect 12969 19904 12981 19907
rect 12860 19876 12981 19904
rect 12860 19864 12866 19876
rect 12969 19873 12981 19876
rect 13015 19873 13027 19907
rect 12969 19867 13027 19873
rect 15657 19907 15715 19913
rect 15657 19873 15669 19907
rect 15703 19904 15715 19907
rect 16482 19904 16488 19916
rect 15703 19876 16488 19904
rect 15703 19873 15715 19876
rect 15657 19867 15715 19873
rect 16482 19864 16488 19876
rect 16540 19864 16546 19916
rect 16942 19864 16948 19916
rect 17000 19904 17006 19916
rect 17000 19876 17632 19904
rect 17000 19864 17006 19876
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19836 8631 19839
rect 8754 19836 8760 19848
rect 8619 19808 8760 19836
rect 8619 19805 8631 19808
rect 8573 19799 8631 19805
rect 8754 19796 8760 19808
rect 8812 19796 8818 19848
rect 11238 19836 11244 19848
rect 11199 19808 11244 19836
rect 11238 19796 11244 19808
rect 11296 19796 11302 19848
rect 11698 19836 11704 19848
rect 11659 19808 11704 19836
rect 11698 19796 11704 19808
rect 11756 19796 11762 19848
rect 12710 19836 12716 19848
rect 12671 19808 12716 19836
rect 12710 19796 12716 19808
rect 12768 19796 12774 19848
rect 15746 19796 15752 19848
rect 15804 19836 15810 19848
rect 17604 19845 17632 19876
rect 18506 19864 18512 19916
rect 18564 19904 18570 19916
rect 24688 19913 24716 20000
rect 18969 19907 19027 19913
rect 18969 19904 18981 19907
rect 18564 19876 18981 19904
rect 18564 19864 18570 19876
rect 18969 19873 18981 19876
rect 19015 19873 19027 19907
rect 18969 19867 19027 19873
rect 19429 19907 19487 19913
rect 19429 19873 19441 19907
rect 19475 19904 19487 19907
rect 23753 19907 23811 19913
rect 19475 19876 21956 19904
rect 19475 19873 19487 19876
rect 19429 19867 19487 19873
rect 15841 19839 15899 19845
rect 15841 19836 15853 19839
rect 15804 19808 15853 19836
rect 15804 19796 15810 19808
rect 15841 19805 15853 19808
rect 15887 19805 15899 19839
rect 15841 19799 15899 19805
rect 17589 19839 17647 19845
rect 17589 19805 17601 19839
rect 17635 19805 17647 19839
rect 17589 19799 17647 19805
rect 18417 19839 18475 19845
rect 18417 19805 18429 19839
rect 18463 19836 18475 19839
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 18463 19808 19257 19836
rect 18463 19805 18475 19808
rect 18417 19799 18475 19805
rect 19245 19805 19257 19808
rect 19291 19836 19303 19839
rect 20898 19836 20904 19848
rect 19291 19808 20392 19836
rect 20859 19808 20904 19836
rect 19291 19805 19303 19808
rect 19245 19799 19303 19805
rect 1412 19740 3924 19768
rect 4154 19728 4160 19780
rect 4212 19768 4218 19780
rect 5077 19771 5135 19777
rect 5077 19768 5089 19771
rect 4212 19740 5089 19768
rect 4212 19728 4218 19740
rect 5077 19737 5089 19740
rect 5123 19768 5135 19771
rect 5442 19768 5448 19780
rect 5123 19740 5448 19768
rect 5123 19737 5135 19740
rect 5077 19731 5135 19737
rect 5442 19728 5448 19740
rect 5500 19728 5506 19780
rect 7926 19768 7932 19780
rect 7887 19740 7932 19768
rect 7926 19728 7932 19740
rect 7984 19728 7990 19780
rect 9125 19771 9183 19777
rect 9125 19737 9137 19771
rect 9171 19768 9183 19771
rect 9582 19768 9588 19780
rect 9171 19740 9588 19768
rect 9171 19737 9183 19740
rect 9125 19731 9183 19737
rect 9582 19728 9588 19740
rect 9640 19768 9646 19780
rect 10689 19771 10747 19777
rect 10689 19768 10701 19771
rect 9640 19740 10701 19768
rect 9640 19728 9646 19740
rect 10689 19737 10701 19740
rect 10735 19737 10747 19771
rect 10689 19731 10747 19737
rect 10778 19728 10784 19780
rect 10836 19768 10842 19780
rect 11146 19768 11152 19780
rect 10836 19740 11152 19768
rect 10836 19728 10842 19740
rect 11146 19728 11152 19740
rect 11204 19728 11210 19780
rect 13814 19728 13820 19780
rect 13872 19768 13878 19780
rect 14274 19768 14280 19780
rect 13872 19740 14280 19768
rect 13872 19728 13878 19740
rect 14274 19728 14280 19740
rect 14332 19768 14338 19780
rect 14645 19771 14703 19777
rect 14645 19768 14657 19771
rect 14332 19740 14657 19768
rect 14332 19728 14338 19740
rect 14645 19737 14657 19740
rect 14691 19737 14703 19771
rect 17034 19768 17040 19780
rect 16995 19740 17040 19768
rect 14645 19731 14703 19737
rect 17034 19728 17040 19740
rect 17092 19728 17098 19780
rect 19334 19728 19340 19780
rect 19392 19768 19398 19780
rect 19429 19771 19487 19777
rect 19429 19768 19441 19771
rect 19392 19740 19441 19768
rect 19392 19728 19398 19740
rect 19429 19737 19441 19740
rect 19475 19737 19487 19771
rect 19429 19731 19487 19737
rect 1486 19660 1492 19712
rect 1544 19700 1550 19712
rect 2409 19703 2467 19709
rect 2409 19700 2421 19703
rect 1544 19672 2421 19700
rect 1544 19660 1550 19672
rect 2409 19669 2421 19672
rect 2455 19669 2467 19703
rect 4246 19700 4252 19712
rect 4207 19672 4252 19700
rect 2409 19663 2467 19669
rect 4246 19660 4252 19672
rect 4304 19660 4310 19712
rect 4338 19660 4344 19712
rect 4396 19700 4402 19712
rect 4706 19700 4712 19712
rect 4396 19672 4712 19700
rect 4396 19660 4402 19672
rect 4706 19660 4712 19672
rect 4764 19700 4770 19712
rect 7466 19700 7472 19712
rect 4764 19672 7472 19700
rect 4764 19660 4770 19672
rect 7466 19660 7472 19672
rect 7524 19660 7530 19712
rect 9490 19700 9496 19712
rect 9451 19672 9496 19700
rect 9490 19660 9496 19672
rect 9548 19700 9554 19712
rect 9858 19700 9864 19712
rect 9548 19672 9864 19700
rect 9548 19660 9554 19672
rect 9858 19660 9864 19672
rect 9916 19660 9922 19712
rect 13998 19660 14004 19712
rect 14056 19700 14062 19712
rect 14093 19703 14151 19709
rect 14093 19700 14105 19703
rect 14056 19672 14105 19700
rect 14056 19660 14062 19672
rect 14093 19669 14105 19672
rect 14139 19700 14151 19703
rect 14550 19700 14556 19712
rect 14139 19672 14556 19700
rect 14139 19669 14151 19672
rect 14093 19663 14151 19669
rect 14550 19660 14556 19672
rect 14608 19660 14614 19712
rect 15289 19703 15347 19709
rect 15289 19669 15301 19703
rect 15335 19700 15347 19703
rect 15378 19700 15384 19712
rect 15335 19672 15384 19700
rect 15335 19669 15347 19672
rect 15289 19663 15347 19669
rect 15378 19660 15384 19672
rect 15436 19660 15442 19712
rect 16942 19700 16948 19712
rect 16903 19672 16948 19700
rect 16942 19660 16948 19672
rect 17000 19660 17006 19712
rect 18598 19700 18604 19712
rect 18559 19672 18604 19700
rect 18598 19660 18604 19672
rect 18656 19660 18662 19712
rect 20364 19709 20392 19808
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 20714 19768 20720 19780
rect 20675 19740 20720 19768
rect 20714 19728 20720 19740
rect 20772 19728 20778 19780
rect 21928 19768 21956 19876
rect 23753 19873 23765 19907
rect 23799 19873 23811 19907
rect 24673 19907 24731 19913
rect 24673 19904 24685 19907
rect 24583 19876 24685 19904
rect 23753 19867 23811 19873
rect 24673 19873 24685 19876
rect 24719 19904 24731 19907
rect 24937 19907 24995 19913
rect 24937 19904 24949 19907
rect 24719 19876 24949 19904
rect 24719 19873 24731 19876
rect 24673 19867 24731 19873
rect 24937 19873 24949 19876
rect 24983 19873 24995 19907
rect 24937 19867 24995 19873
rect 22002 19796 22008 19848
rect 22060 19836 22066 19848
rect 22833 19839 22891 19845
rect 22833 19836 22845 19839
rect 22060 19808 22845 19836
rect 22060 19796 22066 19808
rect 22833 19805 22845 19808
rect 22879 19836 22891 19839
rect 23768 19836 23796 19867
rect 24026 19836 24032 19848
rect 22879 19808 23796 19836
rect 23987 19808 24032 19836
rect 22879 19805 22891 19808
rect 22833 19799 22891 19805
rect 24026 19796 24032 19808
rect 24084 19796 24090 19848
rect 26326 19768 26332 19780
rect 21928 19740 26332 19768
rect 26326 19728 26332 19740
rect 26384 19728 26390 19780
rect 20349 19703 20407 19709
rect 20349 19669 20361 19703
rect 20395 19700 20407 19703
rect 20438 19700 20444 19712
rect 20395 19672 20444 19700
rect 20395 19669 20407 19672
rect 20349 19663 20407 19669
rect 20438 19660 20444 19672
rect 20496 19660 20502 19712
rect 22186 19660 22192 19712
rect 22244 19700 22250 19712
rect 22281 19703 22339 19709
rect 22281 19700 22293 19703
rect 22244 19672 22293 19700
rect 22244 19660 22250 19672
rect 22281 19669 22293 19672
rect 22327 19669 22339 19703
rect 22281 19663 22339 19669
rect 23106 19660 23112 19712
rect 23164 19700 23170 19712
rect 23385 19703 23443 19709
rect 23385 19700 23397 19703
rect 23164 19672 23397 19700
rect 23164 19660 23170 19672
rect 23385 19669 23397 19672
rect 23431 19669 23443 19703
rect 23385 19663 23443 19669
rect 24673 19703 24731 19709
rect 24673 19669 24685 19703
rect 24719 19700 24731 19703
rect 24946 19700 24952 19712
rect 24719 19672 24952 19700
rect 24719 19669 24731 19672
rect 24673 19663 24731 19669
rect 24946 19660 24952 19672
rect 25004 19660 25010 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1762 19456 1768 19508
rect 1820 19496 1826 19508
rect 2130 19496 2136 19508
rect 1820 19468 2136 19496
rect 1820 19456 1826 19468
rect 2130 19456 2136 19468
rect 2188 19456 2194 19508
rect 7558 19456 7564 19508
rect 7616 19496 7622 19508
rect 7837 19499 7895 19505
rect 7837 19496 7849 19499
rect 7616 19468 7849 19496
rect 7616 19456 7622 19468
rect 7837 19465 7849 19468
rect 7883 19465 7895 19499
rect 7837 19459 7895 19465
rect 3050 19320 3056 19372
rect 3108 19360 3114 19372
rect 3789 19363 3847 19369
rect 3789 19360 3801 19363
rect 3108 19332 3801 19360
rect 3108 19320 3114 19332
rect 3789 19329 3801 19332
rect 3835 19360 3847 19363
rect 7852 19360 7880 19459
rect 8294 19456 8300 19508
rect 8352 19496 8358 19508
rect 9401 19499 9459 19505
rect 8352 19468 8975 19496
rect 8352 19456 8358 19468
rect 8947 19428 8975 19468
rect 9401 19465 9413 19499
rect 9447 19496 9459 19499
rect 9490 19496 9496 19508
rect 9447 19468 9496 19496
rect 9447 19465 9459 19468
rect 9401 19459 9459 19465
rect 9490 19456 9496 19468
rect 9548 19456 9554 19508
rect 12710 19496 12716 19508
rect 12671 19468 12716 19496
rect 12710 19456 12716 19468
rect 12768 19456 12774 19508
rect 16574 19496 16580 19508
rect 13648 19468 16580 19496
rect 8947 19400 9076 19428
rect 8021 19363 8079 19369
rect 8021 19360 8033 19363
rect 3835 19332 4384 19360
rect 3835 19329 3847 19332
rect 3789 19323 3847 19329
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19261 1823 19295
rect 1765 19255 1823 19261
rect 4065 19295 4123 19301
rect 4065 19261 4077 19295
rect 4111 19292 4123 19295
rect 4249 19295 4307 19301
rect 4249 19292 4261 19295
rect 4111 19264 4261 19292
rect 4111 19261 4123 19264
rect 4065 19255 4123 19261
rect 4249 19261 4261 19264
rect 4295 19261 4307 19295
rect 4356 19292 4384 19332
rect 6748 19332 8033 19360
rect 4522 19301 4528 19304
rect 4516 19292 4528 19301
rect 4356 19264 4528 19292
rect 4249 19255 4307 19261
rect 4516 19255 4528 19264
rect 4580 19292 4586 19304
rect 5258 19292 5264 19304
rect 4580 19264 5264 19292
rect 1673 19159 1731 19165
rect 1673 19125 1685 19159
rect 1719 19156 1731 19159
rect 1780 19156 1808 19255
rect 2032 19227 2090 19233
rect 2032 19193 2044 19227
rect 2078 19224 2090 19227
rect 2498 19224 2504 19236
rect 2078 19196 2504 19224
rect 2078 19193 2090 19196
rect 2032 19187 2090 19193
rect 2498 19184 2504 19196
rect 2556 19224 2562 19236
rect 3234 19224 3240 19236
rect 2556 19196 3240 19224
rect 2556 19184 2562 19196
rect 3234 19184 3240 19196
rect 3292 19224 3298 19236
rect 4154 19224 4160 19236
rect 3292 19196 4160 19224
rect 3292 19184 3298 19196
rect 4154 19184 4160 19196
rect 4212 19184 4218 19236
rect 4264 19224 4292 19255
rect 4522 19252 4528 19255
rect 4580 19252 4586 19264
rect 5258 19252 5264 19264
rect 5316 19252 5322 19304
rect 6748 19292 6776 19332
rect 8021 19329 8033 19332
rect 8067 19329 8079 19363
rect 9048 19360 9076 19400
rect 11514 19388 11520 19440
rect 11572 19428 11578 19440
rect 12161 19431 12219 19437
rect 12161 19428 12173 19431
rect 11572 19400 12173 19428
rect 11572 19388 11578 19400
rect 12161 19397 12173 19400
rect 12207 19397 12219 19431
rect 13648 19428 13676 19468
rect 16574 19456 16580 19468
rect 16632 19456 16638 19508
rect 16850 19496 16856 19508
rect 16811 19468 16856 19496
rect 16850 19456 16856 19468
rect 16908 19456 16914 19508
rect 17402 19496 17408 19508
rect 17363 19468 17408 19496
rect 17402 19456 17408 19468
rect 17460 19456 17466 19508
rect 20254 19456 20260 19508
rect 20312 19496 20318 19508
rect 21450 19496 21456 19508
rect 20312 19468 21456 19496
rect 20312 19456 20318 19468
rect 21450 19456 21456 19468
rect 21508 19456 21514 19508
rect 24946 19496 24952 19508
rect 24907 19468 24952 19496
rect 24946 19456 24952 19468
rect 25004 19456 25010 19508
rect 15102 19428 15108 19440
rect 12161 19391 12219 19397
rect 13188 19400 13676 19428
rect 15063 19400 15108 19428
rect 9048 19332 9628 19360
rect 8021 19323 8079 19329
rect 6472 19264 6776 19292
rect 6825 19295 6883 19301
rect 4982 19224 4988 19236
rect 4264 19196 4988 19224
rect 4982 19184 4988 19196
rect 5040 19184 5046 19236
rect 6472 19168 6500 19264
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 9600 19292 9628 19332
rect 11238 19320 11244 19372
rect 11296 19360 11302 19372
rect 11333 19363 11391 19369
rect 11333 19360 11345 19363
rect 11296 19332 11345 19360
rect 11296 19320 11302 19332
rect 11333 19329 11345 19332
rect 11379 19329 11391 19363
rect 11882 19360 11888 19372
rect 11795 19332 11888 19360
rect 11333 19323 11391 19329
rect 11882 19320 11888 19332
rect 11940 19360 11946 19372
rect 13188 19360 13216 19400
rect 15102 19388 15108 19400
rect 15160 19388 15166 19440
rect 20070 19428 20076 19440
rect 19444 19400 20076 19428
rect 11940 19332 13216 19360
rect 11940 19320 11946 19332
rect 13262 19320 13268 19372
rect 13320 19360 13326 19372
rect 13722 19360 13728 19372
rect 13320 19332 13728 19360
rect 13320 19320 13326 19332
rect 13722 19320 13728 19332
rect 13780 19320 13786 19372
rect 14550 19320 14556 19372
rect 14608 19360 14614 19372
rect 15657 19363 15715 19369
rect 15657 19360 15669 19363
rect 14608 19332 15669 19360
rect 14608 19320 14614 19332
rect 15657 19329 15669 19332
rect 15703 19360 15715 19363
rect 15746 19360 15752 19372
rect 15703 19332 15752 19360
rect 15703 19329 15715 19332
rect 15657 19323 15715 19329
rect 15746 19320 15752 19332
rect 15804 19320 15810 19372
rect 18966 19320 18972 19372
rect 19024 19360 19030 19372
rect 19245 19363 19303 19369
rect 19245 19360 19257 19363
rect 19024 19332 19257 19360
rect 19024 19320 19030 19332
rect 19245 19329 19257 19332
rect 19291 19329 19303 19363
rect 19245 19323 19303 19329
rect 6871 19264 7512 19292
rect 9600 19264 10640 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 7484 19168 7512 19264
rect 7926 19184 7932 19236
rect 7984 19224 7990 19236
rect 8266 19227 8324 19233
rect 8266 19224 8278 19227
rect 7984 19196 8278 19224
rect 7984 19184 7990 19196
rect 8266 19193 8278 19196
rect 8312 19193 8324 19227
rect 8266 19187 8324 19193
rect 1946 19156 1952 19168
rect 1719 19128 1952 19156
rect 1719 19125 1731 19128
rect 1673 19119 1731 19125
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 3145 19159 3203 19165
rect 3145 19125 3157 19159
rect 3191 19156 3203 19159
rect 3602 19156 3608 19168
rect 3191 19128 3608 19156
rect 3191 19125 3203 19128
rect 3145 19119 3203 19125
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 5626 19156 5632 19168
rect 5587 19128 5632 19156
rect 5626 19116 5632 19128
rect 5684 19116 5690 19168
rect 6273 19159 6331 19165
rect 6273 19125 6285 19159
rect 6319 19156 6331 19159
rect 6454 19156 6460 19168
rect 6319 19128 6460 19156
rect 6319 19125 6331 19128
rect 6273 19119 6331 19125
rect 6454 19116 6460 19128
rect 6512 19116 6518 19168
rect 6641 19159 6699 19165
rect 6641 19125 6653 19159
rect 6687 19156 6699 19159
rect 6730 19156 6736 19168
rect 6687 19128 6736 19156
rect 6687 19125 6699 19128
rect 6641 19119 6699 19125
rect 6730 19116 6736 19128
rect 6788 19116 6794 19168
rect 6914 19116 6920 19168
rect 6972 19156 6978 19168
rect 7009 19159 7067 19165
rect 7009 19156 7021 19159
rect 6972 19128 7021 19156
rect 6972 19116 6978 19128
rect 7009 19125 7021 19128
rect 7055 19125 7067 19159
rect 7466 19156 7472 19168
rect 7427 19128 7472 19156
rect 7009 19119 7067 19125
rect 7466 19116 7472 19128
rect 7524 19116 7530 19168
rect 10042 19116 10048 19168
rect 10100 19156 10106 19168
rect 10229 19159 10287 19165
rect 10229 19156 10241 19159
rect 10100 19128 10241 19156
rect 10100 19116 10106 19128
rect 10229 19125 10241 19128
rect 10275 19125 10287 19159
rect 10612 19156 10640 19264
rect 10778 19252 10784 19304
rect 10836 19292 10842 19304
rect 12710 19292 12716 19304
rect 10836 19264 12716 19292
rect 10836 19252 10842 19264
rect 12710 19252 12716 19264
rect 12768 19292 12774 19304
rect 14090 19292 14096 19304
rect 12768 19264 14096 19292
rect 12768 19252 12774 19264
rect 14090 19252 14096 19264
rect 14148 19252 14154 19304
rect 14277 19295 14335 19301
rect 14277 19261 14289 19295
rect 14323 19292 14335 19295
rect 15562 19292 15568 19304
rect 14323 19264 15568 19292
rect 14323 19261 14335 19264
rect 14277 19255 14335 19261
rect 15562 19252 15568 19264
rect 15620 19252 15626 19304
rect 16942 19292 16948 19304
rect 16903 19264 16948 19292
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 17954 19252 17960 19304
rect 18012 19292 18018 19304
rect 19058 19292 19064 19304
rect 18012 19264 19064 19292
rect 18012 19252 18018 19264
rect 19058 19252 19064 19264
rect 19116 19252 19122 19304
rect 19444 19292 19472 19400
rect 20070 19388 20076 19400
rect 20128 19388 20134 19440
rect 20714 19388 20720 19440
rect 20772 19428 20778 19440
rect 23106 19428 23112 19440
rect 20772 19400 23112 19428
rect 20772 19388 20778 19400
rect 20438 19320 20444 19372
rect 20496 19360 20502 19372
rect 20901 19363 20959 19369
rect 20901 19360 20913 19363
rect 20496 19332 20913 19360
rect 20496 19320 20502 19332
rect 20901 19329 20913 19332
rect 20947 19360 20959 19363
rect 21174 19360 21180 19372
rect 20947 19332 21180 19360
rect 20947 19329 20959 19332
rect 20901 19323 20959 19329
rect 21174 19320 21180 19332
rect 21232 19320 21238 19372
rect 22480 19369 22508 19400
rect 23106 19388 23112 19400
rect 23164 19388 23170 19440
rect 23477 19431 23535 19437
rect 23477 19397 23489 19431
rect 23523 19428 23535 19431
rect 24026 19428 24032 19440
rect 23523 19400 24032 19428
rect 23523 19397 23535 19400
rect 23477 19391 23535 19397
rect 22465 19363 22523 19369
rect 22465 19329 22477 19363
rect 22511 19329 22523 19363
rect 22646 19360 22652 19372
rect 22607 19332 22652 19360
rect 22465 19323 22523 19329
rect 22646 19320 22652 19332
rect 22704 19320 22710 19372
rect 19260 19264 19472 19292
rect 10689 19227 10747 19233
rect 10689 19193 10701 19227
rect 10735 19224 10747 19227
rect 11149 19227 11207 19233
rect 11149 19224 11161 19227
rect 10735 19196 11161 19224
rect 10735 19193 10747 19196
rect 10689 19187 10747 19193
rect 11149 19193 11161 19196
rect 11195 19224 11207 19227
rect 12250 19224 12256 19236
rect 11195 19196 12256 19224
rect 11195 19193 11207 19196
rect 11149 19187 11207 19193
rect 12250 19184 12256 19196
rect 12308 19224 12314 19236
rect 12618 19224 12624 19236
rect 12308 19196 12624 19224
rect 12308 19184 12314 19196
rect 12618 19184 12624 19196
rect 12676 19184 12682 19236
rect 13814 19224 13820 19236
rect 13188 19196 13820 19224
rect 10781 19159 10839 19165
rect 10781 19156 10793 19159
rect 10612 19128 10793 19156
rect 10229 19119 10287 19125
rect 10781 19125 10793 19128
rect 10827 19125 10839 19159
rect 10781 19119 10839 19125
rect 11054 19116 11060 19168
rect 11112 19156 11118 19168
rect 13188 19165 13216 19196
rect 13814 19184 13820 19196
rect 13872 19184 13878 19236
rect 15473 19227 15531 19233
rect 15473 19193 15485 19227
rect 15519 19224 15531 19227
rect 15838 19224 15844 19236
rect 15519 19196 15844 19224
rect 15519 19193 15531 19196
rect 15473 19187 15531 19193
rect 15838 19184 15844 19196
rect 15896 19184 15902 19236
rect 18598 19184 18604 19236
rect 18656 19224 18662 19236
rect 19153 19227 19211 19233
rect 19153 19224 19165 19227
rect 18656 19196 19165 19224
rect 18656 19184 18662 19196
rect 19153 19193 19165 19196
rect 19199 19193 19211 19227
rect 19153 19187 19211 19193
rect 19260 19168 19288 19264
rect 19518 19252 19524 19304
rect 19576 19292 19582 19304
rect 20073 19295 20131 19301
rect 20073 19292 20085 19295
rect 19576 19264 20085 19292
rect 19576 19252 19582 19264
rect 20073 19261 20085 19264
rect 20119 19292 20131 19295
rect 20717 19295 20775 19301
rect 20717 19292 20729 19295
rect 20119 19264 20729 19292
rect 20119 19261 20131 19264
rect 20073 19255 20131 19261
rect 20717 19261 20729 19264
rect 20763 19261 20775 19295
rect 20717 19255 20775 19261
rect 20990 19252 20996 19304
rect 21048 19292 21054 19304
rect 22094 19292 22100 19304
rect 21048 19264 22100 19292
rect 21048 19252 21054 19264
rect 22094 19252 22100 19264
rect 22152 19252 22158 19304
rect 23106 19292 23112 19304
rect 23019 19264 23112 19292
rect 23106 19252 23112 19264
rect 23164 19292 23170 19304
rect 23492 19292 23520 19391
rect 24026 19388 24032 19400
rect 24084 19428 24090 19440
rect 24084 19400 24256 19428
rect 24084 19388 24090 19400
rect 24228 19369 24256 19400
rect 25130 19388 25136 19440
rect 25188 19428 25194 19440
rect 25188 19400 25636 19428
rect 25188 19388 25194 19400
rect 25608 19372 25636 19400
rect 24213 19363 24271 19369
rect 24213 19329 24225 19363
rect 24259 19329 24271 19363
rect 24213 19323 24271 19329
rect 25590 19320 25596 19372
rect 25648 19320 25654 19372
rect 23164 19264 23520 19292
rect 24029 19295 24087 19301
rect 23164 19252 23170 19264
rect 24029 19261 24041 19295
rect 24075 19292 24087 19295
rect 24118 19292 24124 19304
rect 24075 19264 24124 19292
rect 24075 19261 24087 19264
rect 24029 19255 24087 19261
rect 24118 19252 24124 19264
rect 24176 19252 24182 19304
rect 25130 19252 25136 19304
rect 25188 19292 25194 19304
rect 25225 19295 25283 19301
rect 25225 19292 25237 19295
rect 25188 19264 25237 19292
rect 25188 19252 25194 19264
rect 25225 19261 25237 19264
rect 25271 19292 25283 19295
rect 25777 19295 25835 19301
rect 25777 19292 25789 19295
rect 25271 19264 25789 19292
rect 25271 19261 25283 19264
rect 25225 19255 25283 19261
rect 25777 19261 25789 19264
rect 25823 19261 25835 19295
rect 25777 19255 25835 19261
rect 19334 19184 19340 19236
rect 19392 19224 19398 19236
rect 19705 19227 19763 19233
rect 19705 19224 19717 19227
rect 19392 19196 19717 19224
rect 19392 19184 19398 19196
rect 19705 19193 19717 19196
rect 19751 19193 19763 19227
rect 19705 19187 19763 19193
rect 21266 19184 21272 19236
rect 21324 19224 21330 19236
rect 21637 19227 21695 19233
rect 21637 19224 21649 19227
rect 21324 19196 21649 19224
rect 21324 19184 21330 19196
rect 21637 19193 21649 19196
rect 21683 19193 21695 19227
rect 22370 19224 22376 19236
rect 22283 19196 22376 19224
rect 21637 19187 21695 19193
rect 22370 19184 22376 19196
rect 22428 19224 22434 19236
rect 22428 19196 23704 19224
rect 22428 19184 22434 19196
rect 11241 19159 11299 19165
rect 11241 19156 11253 19159
rect 11112 19128 11253 19156
rect 11112 19116 11118 19128
rect 11241 19125 11253 19128
rect 11287 19125 11299 19159
rect 11241 19119 11299 19125
rect 13173 19159 13231 19165
rect 13173 19125 13185 19159
rect 13219 19125 13231 19159
rect 13538 19156 13544 19168
rect 13499 19128 13544 19156
rect 13173 19119 13231 19125
rect 13538 19116 13544 19128
rect 13596 19116 13602 19168
rect 13630 19116 13636 19168
rect 13688 19156 13694 19168
rect 14550 19156 14556 19168
rect 13688 19128 13733 19156
rect 14511 19128 14556 19156
rect 13688 19116 13694 19128
rect 14550 19116 14556 19128
rect 14608 19156 14614 19168
rect 14921 19159 14979 19165
rect 14921 19156 14933 19159
rect 14608 19128 14933 19156
rect 14608 19116 14614 19128
rect 14921 19125 14933 19128
rect 14967 19125 14979 19159
rect 16206 19156 16212 19168
rect 16167 19128 16212 19156
rect 14921 19119 14979 19125
rect 16206 19116 16212 19128
rect 16264 19156 16270 19168
rect 16482 19156 16488 19168
rect 16264 19128 16488 19156
rect 16264 19116 16270 19128
rect 16482 19116 16488 19128
rect 16540 19116 16546 19168
rect 17126 19156 17132 19168
rect 17087 19128 17132 19156
rect 17126 19116 17132 19128
rect 17184 19116 17190 19168
rect 17770 19156 17776 19168
rect 17731 19128 17776 19156
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 18506 19156 18512 19168
rect 18467 19128 18512 19156
rect 18506 19116 18512 19128
rect 18564 19116 18570 19168
rect 18690 19156 18696 19168
rect 18651 19128 18696 19156
rect 18690 19116 18696 19128
rect 18748 19116 18754 19168
rect 19242 19116 19248 19168
rect 19300 19116 19306 19168
rect 20254 19156 20260 19168
rect 20215 19128 20260 19156
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 20438 19116 20444 19168
rect 20496 19156 20502 19168
rect 20625 19159 20683 19165
rect 20625 19156 20637 19159
rect 20496 19128 20637 19156
rect 20496 19116 20502 19128
rect 20625 19125 20637 19128
rect 20671 19125 20683 19159
rect 20625 19119 20683 19125
rect 20898 19116 20904 19168
rect 20956 19156 20962 19168
rect 21361 19159 21419 19165
rect 21361 19156 21373 19159
rect 20956 19128 21373 19156
rect 20956 19116 20962 19128
rect 21361 19125 21373 19128
rect 21407 19156 21419 19159
rect 21542 19156 21548 19168
rect 21407 19128 21548 19156
rect 21407 19125 21419 19128
rect 21361 19119 21419 19125
rect 21542 19116 21548 19128
rect 21600 19116 21606 19168
rect 21726 19116 21732 19168
rect 21784 19156 21790 19168
rect 23676 19165 23704 19196
rect 22005 19159 22063 19165
rect 22005 19156 22017 19159
rect 21784 19128 22017 19156
rect 21784 19116 21790 19128
rect 22005 19125 22017 19128
rect 22051 19125 22063 19159
rect 22005 19119 22063 19125
rect 23661 19159 23719 19165
rect 23661 19125 23673 19159
rect 23707 19125 23719 19159
rect 23661 19119 23719 19125
rect 24121 19159 24179 19165
rect 24121 19125 24133 19159
rect 24167 19156 24179 19159
rect 24210 19156 24216 19168
rect 24167 19128 24216 19156
rect 24167 19125 24179 19128
rect 24121 19119 24179 19125
rect 24210 19116 24216 19128
rect 24268 19116 24274 19168
rect 25409 19159 25467 19165
rect 25409 19125 25421 19159
rect 25455 19156 25467 19159
rect 25682 19156 25688 19168
rect 25455 19128 25688 19156
rect 25455 19125 25467 19128
rect 25409 19119 25467 19125
rect 25682 19116 25688 19128
rect 25740 19116 25746 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18921 1639 18955
rect 1581 18915 1639 18921
rect 1596 18884 1624 18915
rect 2774 18912 2780 18964
rect 2832 18952 2838 18964
rect 2832 18924 2877 18952
rect 2832 18912 2838 18924
rect 4522 18912 4528 18964
rect 4580 18952 4586 18964
rect 4617 18955 4675 18961
rect 4617 18952 4629 18955
rect 4580 18924 4629 18952
rect 4580 18912 4586 18924
rect 4617 18921 4629 18924
rect 4663 18921 4675 18955
rect 4617 18915 4675 18921
rect 5442 18912 5448 18964
rect 5500 18952 5506 18964
rect 6733 18955 6791 18961
rect 6733 18952 6745 18955
rect 5500 18924 6745 18952
rect 5500 18912 5506 18924
rect 6733 18921 6745 18924
rect 6779 18921 6791 18955
rect 8018 18952 8024 18964
rect 7979 18924 8024 18952
rect 6733 18915 6791 18921
rect 8018 18912 8024 18924
rect 8076 18912 8082 18964
rect 10042 18912 10048 18964
rect 10100 18952 10106 18964
rect 11054 18952 11060 18964
rect 10100 18924 11060 18952
rect 10100 18912 10106 18924
rect 11054 18912 11060 18924
rect 11112 18912 11118 18964
rect 12161 18955 12219 18961
rect 12161 18921 12173 18955
rect 12207 18921 12219 18955
rect 12802 18952 12808 18964
rect 12763 18924 12808 18952
rect 12161 18915 12219 18921
rect 2498 18884 2504 18896
rect 1596 18856 2504 18884
rect 2498 18844 2504 18856
rect 2556 18844 2562 18896
rect 2590 18844 2596 18896
rect 2648 18884 2654 18896
rect 2869 18887 2927 18893
rect 2869 18884 2881 18887
rect 2648 18856 2881 18884
rect 2648 18844 2654 18856
rect 2869 18853 2881 18856
rect 2915 18884 2927 18887
rect 3326 18884 3332 18896
rect 2915 18856 3332 18884
rect 2915 18853 2927 18856
rect 2869 18847 2927 18853
rect 3326 18844 3332 18856
rect 3384 18844 3390 18896
rect 5626 18893 5632 18896
rect 5620 18884 5632 18893
rect 4356 18856 5632 18884
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 1578 18816 1584 18828
rect 1443 18788 1584 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 1578 18776 1584 18788
rect 1636 18816 1642 18828
rect 2406 18816 2412 18828
rect 1636 18788 2412 18816
rect 1636 18776 1642 18788
rect 2406 18776 2412 18788
rect 2464 18776 2470 18828
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18816 4123 18819
rect 4154 18816 4160 18828
rect 4111 18788 4160 18816
rect 4111 18785 4123 18788
rect 4065 18779 4123 18785
rect 4154 18776 4160 18788
rect 4212 18776 4218 18828
rect 3053 18751 3111 18757
rect 3053 18717 3065 18751
rect 3099 18748 3111 18751
rect 4356 18748 4384 18856
rect 5620 18847 5632 18856
rect 5626 18844 5632 18847
rect 5684 18844 5690 18896
rect 7650 18844 7656 18896
rect 7708 18884 7714 18896
rect 9401 18887 9459 18893
rect 9401 18884 9413 18887
rect 7708 18856 9413 18884
rect 7708 18844 7714 18856
rect 9401 18853 9413 18856
rect 9447 18853 9459 18887
rect 11238 18884 11244 18896
rect 9401 18847 9459 18853
rect 10612 18856 11244 18884
rect 4982 18776 4988 18828
rect 5040 18816 5046 18828
rect 5353 18819 5411 18825
rect 5353 18816 5365 18819
rect 5040 18788 5365 18816
rect 5040 18776 5046 18788
rect 5353 18785 5365 18788
rect 5399 18816 5411 18819
rect 6454 18816 6460 18828
rect 5399 18788 6460 18816
rect 5399 18785 5411 18788
rect 5353 18779 5411 18785
rect 6454 18776 6460 18788
rect 6512 18776 6518 18828
rect 7558 18776 7564 18828
rect 7616 18816 7622 18828
rect 8389 18819 8447 18825
rect 8389 18816 8401 18819
rect 7616 18788 8401 18816
rect 7616 18776 7622 18788
rect 8389 18785 8401 18788
rect 8435 18785 8447 18819
rect 8389 18779 8447 18785
rect 8481 18819 8539 18825
rect 8481 18785 8493 18819
rect 8527 18816 8539 18819
rect 8846 18816 8852 18828
rect 8527 18788 8852 18816
rect 8527 18785 8539 18788
rect 8481 18779 8539 18785
rect 8846 18776 8852 18788
rect 8904 18776 8910 18828
rect 9674 18816 9680 18828
rect 9635 18788 9680 18816
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 10612 18757 10640 18856
rect 11238 18844 11244 18856
rect 11296 18884 11302 18896
rect 12176 18884 12204 18915
rect 12802 18912 12808 18924
rect 12860 18912 12866 18964
rect 13262 18952 13268 18964
rect 13223 18924 13268 18952
rect 13262 18912 13268 18924
rect 13320 18912 13326 18964
rect 13630 18912 13636 18964
rect 13688 18952 13694 18964
rect 14829 18955 14887 18961
rect 14829 18952 14841 18955
rect 13688 18924 14841 18952
rect 13688 18912 13694 18924
rect 14829 18921 14841 18924
rect 14875 18952 14887 18955
rect 15102 18952 15108 18964
rect 14875 18924 15108 18952
rect 14875 18921 14887 18924
rect 14829 18915 14887 18921
rect 15102 18912 15108 18924
rect 15160 18912 15166 18964
rect 15470 18952 15476 18964
rect 15431 18924 15476 18952
rect 15470 18912 15476 18924
rect 15528 18912 15534 18964
rect 15654 18912 15660 18964
rect 15712 18952 15718 18964
rect 16117 18955 16175 18961
rect 16117 18952 16129 18955
rect 15712 18924 16129 18952
rect 15712 18912 15718 18924
rect 16117 18921 16129 18924
rect 16163 18921 16175 18955
rect 16117 18915 16175 18921
rect 17678 18912 17684 18964
rect 17736 18952 17742 18964
rect 17773 18955 17831 18961
rect 17773 18952 17785 18955
rect 17736 18924 17785 18952
rect 17736 18912 17742 18924
rect 17773 18921 17785 18924
rect 17819 18921 17831 18955
rect 17773 18915 17831 18921
rect 19981 18955 20039 18961
rect 19981 18921 19993 18955
rect 20027 18952 20039 18955
rect 20070 18952 20076 18964
rect 20027 18924 20076 18952
rect 20027 18921 20039 18924
rect 19981 18915 20039 18921
rect 20070 18912 20076 18924
rect 20128 18912 20134 18964
rect 20901 18955 20959 18961
rect 20901 18921 20913 18955
rect 20947 18952 20959 18955
rect 22002 18952 22008 18964
rect 20947 18924 22008 18952
rect 20947 18921 20959 18924
rect 20901 18915 20959 18921
rect 22002 18912 22008 18924
rect 22060 18912 22066 18964
rect 22097 18955 22155 18961
rect 22097 18921 22109 18955
rect 22143 18952 22155 18955
rect 22646 18952 22652 18964
rect 22143 18924 22652 18952
rect 22143 18921 22155 18924
rect 22097 18915 22155 18921
rect 22646 18912 22652 18924
rect 22704 18952 22710 18964
rect 23845 18955 23903 18961
rect 23845 18952 23857 18955
rect 22704 18924 23857 18952
rect 22704 18912 22710 18924
rect 23845 18921 23857 18924
rect 23891 18921 23903 18955
rect 23845 18915 23903 18921
rect 24118 18912 24124 18964
rect 24176 18952 24182 18964
rect 24765 18955 24823 18961
rect 24765 18952 24777 18955
rect 24176 18924 24777 18952
rect 24176 18912 24182 18924
rect 24765 18921 24777 18924
rect 24811 18921 24823 18955
rect 24765 18915 24823 18921
rect 25133 18955 25191 18961
rect 25133 18921 25145 18955
rect 25179 18952 25191 18955
rect 25222 18952 25228 18964
rect 25179 18924 25228 18952
rect 25179 18921 25191 18924
rect 25133 18915 25191 18921
rect 25222 18912 25228 18924
rect 25280 18912 25286 18964
rect 11296 18856 12204 18884
rect 11296 18844 11302 18856
rect 13354 18844 13360 18896
rect 13412 18884 13418 18896
rect 13817 18887 13875 18893
rect 13817 18884 13829 18887
rect 13412 18856 13829 18884
rect 13412 18844 13418 18856
rect 13817 18853 13829 18856
rect 13863 18853 13875 18887
rect 15838 18884 15844 18896
rect 15799 18856 15844 18884
rect 13817 18847 13875 18853
rect 15838 18844 15844 18856
rect 15896 18844 15902 18896
rect 20717 18887 20775 18893
rect 20717 18853 20729 18887
rect 20763 18884 20775 18887
rect 21361 18887 21419 18893
rect 21361 18884 21373 18887
rect 20763 18856 21373 18884
rect 20763 18853 20775 18856
rect 20717 18847 20775 18853
rect 21361 18853 21373 18856
rect 21407 18884 21419 18887
rect 21910 18884 21916 18896
rect 21407 18856 21916 18884
rect 21407 18853 21419 18856
rect 21361 18847 21419 18853
rect 21910 18844 21916 18856
rect 21968 18844 21974 18896
rect 22554 18844 22560 18896
rect 22612 18884 22618 18896
rect 22732 18887 22790 18893
rect 22732 18884 22744 18887
rect 22612 18856 22744 18884
rect 22612 18844 22618 18856
rect 22732 18853 22744 18856
rect 22778 18884 22790 18887
rect 23106 18884 23112 18896
rect 22778 18856 23112 18884
rect 22778 18853 22790 18856
rect 22732 18847 22790 18853
rect 23106 18844 23112 18856
rect 23164 18844 23170 18896
rect 10778 18816 10784 18828
rect 10739 18788 10784 18816
rect 10778 18776 10784 18788
rect 10836 18776 10842 18828
rect 11048 18819 11106 18825
rect 11048 18785 11060 18819
rect 11094 18816 11106 18819
rect 11330 18816 11336 18828
rect 11094 18788 11336 18816
rect 11094 18785 11106 18788
rect 11048 18779 11106 18785
rect 11330 18776 11336 18788
rect 11388 18776 11394 18828
rect 13170 18776 13176 18828
rect 13228 18816 13234 18828
rect 13446 18816 13452 18828
rect 13228 18788 13452 18816
rect 13228 18776 13234 18788
rect 13446 18776 13452 18788
rect 13504 18776 13510 18828
rect 13722 18816 13728 18828
rect 13683 18788 13728 18816
rect 13722 18776 13728 18788
rect 13780 18776 13786 18828
rect 15289 18819 15347 18825
rect 15289 18785 15301 18819
rect 15335 18816 15347 18819
rect 15378 18816 15384 18828
rect 15335 18788 15384 18816
rect 15335 18785 15347 18788
rect 15289 18779 15347 18785
rect 15378 18776 15384 18788
rect 15436 18776 15442 18828
rect 16660 18819 16718 18825
rect 16660 18785 16672 18819
rect 16706 18816 16718 18819
rect 17402 18816 17408 18828
rect 16706 18788 17408 18816
rect 16706 18785 16718 18788
rect 16660 18779 16718 18785
rect 17402 18776 17408 18788
rect 17460 18776 17466 18828
rect 19058 18776 19064 18828
rect 19116 18816 19122 18828
rect 19245 18819 19303 18825
rect 19245 18816 19257 18819
rect 19116 18788 19257 18816
rect 19116 18776 19122 18788
rect 19245 18785 19257 18788
rect 19291 18785 19303 18819
rect 19245 18779 19303 18785
rect 19337 18819 19395 18825
rect 19337 18785 19349 18819
rect 19383 18816 19395 18819
rect 20254 18816 20260 18828
rect 19383 18788 20260 18816
rect 19383 18785 19395 18788
rect 19337 18779 19395 18785
rect 20254 18776 20260 18788
rect 20312 18776 20318 18828
rect 20990 18776 20996 18828
rect 21048 18816 21054 18828
rect 21269 18819 21327 18825
rect 21269 18816 21281 18819
rect 21048 18788 21281 18816
rect 21048 18776 21054 18788
rect 21269 18785 21281 18788
rect 21315 18785 21327 18819
rect 21269 18779 21327 18785
rect 22465 18819 22523 18825
rect 22465 18785 22477 18819
rect 22511 18816 22523 18819
rect 23014 18816 23020 18828
rect 22511 18788 23020 18816
rect 22511 18785 22523 18788
rect 22465 18779 22523 18785
rect 3099 18720 4384 18748
rect 8573 18751 8631 18757
rect 3099 18717 3111 18720
rect 3053 18711 3111 18717
rect 8573 18717 8585 18751
rect 8619 18748 8631 18751
rect 10229 18751 10287 18757
rect 10229 18748 10241 18751
rect 8619 18720 10241 18748
rect 8619 18717 8631 18720
rect 8573 18711 8631 18717
rect 10229 18717 10241 18720
rect 10275 18748 10287 18751
rect 10597 18751 10655 18757
rect 10597 18748 10609 18751
rect 10275 18720 10609 18748
rect 10275 18717 10287 18720
rect 10229 18711 10287 18717
rect 10597 18717 10609 18720
rect 10643 18717 10655 18751
rect 10597 18711 10655 18717
rect 13909 18751 13967 18757
rect 13909 18717 13921 18751
rect 13955 18748 13967 18751
rect 14550 18748 14556 18760
rect 13955 18720 14556 18748
rect 13955 18717 13967 18720
rect 13909 18711 13967 18717
rect 2498 18640 2504 18692
rect 2556 18680 2562 18692
rect 3068 18680 3096 18711
rect 2556 18652 3096 18680
rect 2556 18640 2562 18652
rect 7098 18640 7104 18692
rect 7156 18680 7162 18692
rect 8588 18680 8616 18711
rect 7156 18652 8616 18680
rect 7156 18640 7162 18652
rect 8662 18640 8668 18692
rect 8720 18680 8726 18692
rect 9861 18683 9919 18689
rect 9861 18680 9873 18683
rect 8720 18652 9873 18680
rect 8720 18640 8726 18652
rect 9861 18649 9873 18652
rect 9907 18649 9919 18683
rect 9861 18643 9919 18649
rect 13446 18640 13452 18692
rect 13504 18680 13510 18692
rect 13924 18680 13952 18711
rect 14550 18708 14556 18720
rect 14608 18708 14614 18760
rect 15838 18708 15844 18760
rect 15896 18748 15902 18760
rect 16393 18751 16451 18757
rect 16393 18748 16405 18751
rect 15896 18720 16405 18748
rect 15896 18708 15902 18720
rect 16393 18717 16405 18720
rect 16439 18717 16451 18751
rect 16393 18711 16451 18717
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18748 18475 18751
rect 19426 18748 19432 18760
rect 18463 18720 19432 18748
rect 18463 18717 18475 18720
rect 18417 18711 18475 18717
rect 19426 18708 19432 18720
rect 19484 18708 19490 18760
rect 21450 18708 21456 18760
rect 21508 18748 21514 18760
rect 21508 18720 21553 18748
rect 21508 18708 21514 18720
rect 13504 18652 13952 18680
rect 13504 18640 13510 18652
rect 20070 18640 20076 18692
rect 20128 18680 20134 18692
rect 20622 18680 20628 18692
rect 20128 18652 20628 18680
rect 20128 18640 20134 18652
rect 20622 18640 20628 18652
rect 20680 18640 20686 18692
rect 1946 18612 1952 18624
rect 1907 18584 1952 18612
rect 1946 18572 1952 18584
rect 2004 18572 2010 18624
rect 2409 18615 2467 18621
rect 2409 18581 2421 18615
rect 2455 18612 2467 18615
rect 3050 18612 3056 18624
rect 2455 18584 3056 18612
rect 2455 18581 2467 18584
rect 2409 18575 2467 18581
rect 3050 18572 3056 18584
rect 3108 18572 3114 18624
rect 3234 18572 3240 18624
rect 3292 18612 3298 18624
rect 3421 18615 3479 18621
rect 3421 18612 3433 18615
rect 3292 18584 3433 18612
rect 3292 18572 3298 18584
rect 3421 18581 3433 18584
rect 3467 18612 3479 18615
rect 3789 18615 3847 18621
rect 3789 18612 3801 18615
rect 3467 18584 3801 18612
rect 3467 18581 3479 18584
rect 3421 18575 3479 18581
rect 3789 18581 3801 18584
rect 3835 18581 3847 18615
rect 3789 18575 3847 18581
rect 3970 18572 3976 18624
rect 4028 18612 4034 18624
rect 4249 18615 4307 18621
rect 4249 18612 4261 18615
rect 4028 18584 4261 18612
rect 4028 18572 4034 18584
rect 4249 18581 4261 18584
rect 4295 18581 4307 18615
rect 5258 18612 5264 18624
rect 5219 18584 5264 18612
rect 4249 18575 4307 18581
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 6730 18572 6736 18624
rect 6788 18612 6794 18624
rect 7561 18615 7619 18621
rect 7561 18612 7573 18615
rect 6788 18584 7573 18612
rect 6788 18572 6794 18584
rect 7561 18581 7573 18584
rect 7607 18612 7619 18615
rect 7834 18612 7840 18624
rect 7607 18584 7840 18612
rect 7607 18581 7619 18584
rect 7561 18575 7619 18581
rect 7834 18572 7840 18584
rect 7892 18572 7898 18624
rect 7926 18572 7932 18624
rect 7984 18612 7990 18624
rect 9030 18612 9036 18624
rect 7984 18584 8029 18612
rect 8991 18584 9036 18612
rect 7984 18572 7990 18584
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 13357 18615 13415 18621
rect 13357 18581 13369 18615
rect 13403 18612 13415 18615
rect 13630 18612 13636 18624
rect 13403 18584 13636 18612
rect 13403 18581 13415 18584
rect 13357 18575 13415 18581
rect 13630 18572 13636 18584
rect 13688 18572 13694 18624
rect 14366 18612 14372 18624
rect 14327 18584 14372 18612
rect 14366 18572 14372 18584
rect 14424 18572 14430 18624
rect 17954 18572 17960 18624
rect 18012 18612 18018 18624
rect 18693 18615 18751 18621
rect 18693 18612 18705 18615
rect 18012 18584 18705 18612
rect 18012 18572 18018 18584
rect 18693 18581 18705 18584
rect 18739 18581 18751 18615
rect 18874 18612 18880 18624
rect 18835 18584 18880 18612
rect 18693 18575 18751 18581
rect 18874 18572 18880 18584
rect 18932 18572 18938 18624
rect 20349 18615 20407 18621
rect 20349 18581 20361 18615
rect 20395 18612 20407 18615
rect 20438 18612 20444 18624
rect 20395 18584 20444 18612
rect 20395 18581 20407 18584
rect 20349 18575 20407 18581
rect 20438 18572 20444 18584
rect 20496 18572 20502 18624
rect 21542 18572 21548 18624
rect 21600 18612 21606 18624
rect 22480 18612 22508 18779
rect 23014 18776 23020 18788
rect 23072 18776 23078 18828
rect 24118 18776 24124 18828
rect 24176 18816 24182 18828
rect 24302 18816 24308 18828
rect 24176 18788 24308 18816
rect 24176 18776 24182 18788
rect 24302 18776 24308 18788
rect 24360 18776 24366 18828
rect 24946 18816 24952 18828
rect 24907 18788 24952 18816
rect 24946 18776 24952 18788
rect 25004 18776 25010 18828
rect 22738 18612 22744 18624
rect 21600 18584 22744 18612
rect 21600 18572 21606 18584
rect 22738 18572 22744 18584
rect 22796 18572 22802 18624
rect 24210 18572 24216 18624
rect 24268 18612 24274 18624
rect 24397 18615 24455 18621
rect 24397 18612 24409 18615
rect 24268 18584 24409 18612
rect 24268 18572 24274 18584
rect 24397 18581 24409 18584
rect 24443 18581 24455 18615
rect 24397 18575 24455 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1857 18411 1915 18417
rect 1857 18377 1869 18411
rect 1903 18408 1915 18411
rect 2866 18408 2872 18420
rect 1903 18380 2872 18408
rect 1903 18377 1915 18380
rect 1857 18371 1915 18377
rect 2866 18368 2872 18380
rect 2924 18368 2930 18420
rect 4154 18408 4160 18420
rect 4115 18380 4160 18408
rect 4154 18368 4160 18380
rect 4212 18368 4218 18420
rect 5077 18411 5135 18417
rect 5077 18377 5089 18411
rect 5123 18408 5135 18411
rect 5534 18408 5540 18420
rect 5123 18380 5540 18408
rect 5123 18377 5135 18380
rect 5077 18371 5135 18377
rect 5534 18368 5540 18380
rect 5592 18368 5598 18420
rect 6273 18411 6331 18417
rect 6273 18377 6285 18411
rect 6319 18408 6331 18411
rect 6454 18408 6460 18420
rect 6319 18380 6460 18408
rect 6319 18377 6331 18380
rect 6273 18371 6331 18377
rect 6454 18368 6460 18380
rect 6512 18368 6518 18420
rect 7098 18408 7104 18420
rect 7059 18380 7104 18408
rect 7098 18368 7104 18380
rect 7156 18368 7162 18420
rect 8386 18368 8392 18420
rect 8444 18408 8450 18420
rect 9217 18411 9275 18417
rect 9217 18408 9229 18411
rect 8444 18380 9229 18408
rect 8444 18368 8450 18380
rect 9217 18377 9229 18380
rect 9263 18377 9275 18411
rect 9217 18371 9275 18377
rect 9674 18368 9680 18420
rect 9732 18408 9738 18420
rect 10229 18411 10287 18417
rect 10229 18408 10241 18411
rect 9732 18380 10241 18408
rect 9732 18368 9738 18380
rect 10229 18377 10241 18380
rect 10275 18377 10287 18411
rect 10229 18371 10287 18377
rect 10778 18368 10784 18420
rect 10836 18408 10842 18420
rect 11146 18408 11152 18420
rect 10836 18380 11152 18408
rect 10836 18368 10842 18380
rect 11146 18368 11152 18380
rect 11204 18368 11210 18420
rect 13354 18368 13360 18420
rect 13412 18408 13418 18420
rect 13449 18411 13507 18417
rect 13449 18408 13461 18411
rect 13412 18380 13461 18408
rect 13412 18368 13418 18380
rect 13449 18377 13461 18380
rect 13495 18377 13507 18411
rect 13449 18371 13507 18377
rect 13722 18368 13728 18420
rect 13780 18408 13786 18420
rect 13817 18411 13875 18417
rect 13817 18408 13829 18411
rect 13780 18380 13829 18408
rect 13780 18368 13786 18380
rect 13817 18377 13829 18380
rect 13863 18408 13875 18411
rect 13863 18380 14044 18408
rect 13863 18377 13875 18380
rect 13817 18371 13875 18377
rect 4338 18300 4344 18352
rect 4396 18340 4402 18352
rect 4433 18343 4491 18349
rect 4433 18340 4445 18343
rect 4396 18312 4445 18340
rect 4396 18300 4402 18312
rect 4433 18309 4445 18312
rect 4479 18309 4491 18343
rect 4433 18303 4491 18309
rect 7834 18300 7840 18352
rect 7892 18340 7898 18352
rect 8754 18340 8760 18352
rect 7892 18312 8760 18340
rect 7892 18300 7898 18312
rect 8754 18300 8760 18312
rect 8812 18340 8818 18352
rect 9125 18343 9183 18349
rect 9125 18340 9137 18343
rect 8812 18312 9137 18340
rect 8812 18300 8818 18312
rect 9125 18309 9137 18312
rect 9171 18340 9183 18343
rect 9171 18312 9812 18340
rect 9171 18309 9183 18312
rect 9125 18303 9183 18309
rect 5258 18232 5264 18284
rect 5316 18272 5322 18284
rect 5813 18275 5871 18281
rect 5813 18272 5825 18275
rect 5316 18244 5825 18272
rect 5316 18232 5322 18244
rect 5813 18241 5825 18244
rect 5859 18272 5871 18275
rect 6641 18275 6699 18281
rect 5859 18244 6132 18272
rect 5859 18241 5871 18244
rect 5813 18235 5871 18241
rect 1946 18204 1952 18216
rect 1907 18176 1952 18204
rect 1946 18164 1952 18176
rect 2004 18164 2010 18216
rect 6104 18204 6132 18244
rect 6641 18241 6653 18275
rect 6687 18272 6699 18275
rect 8110 18272 8116 18284
rect 6687 18244 8116 18272
rect 6687 18241 6699 18244
rect 6641 18235 6699 18241
rect 8110 18232 8116 18244
rect 8168 18232 8174 18284
rect 8202 18232 8208 18284
rect 8260 18272 8266 18284
rect 8260 18244 8305 18272
rect 8260 18232 8266 18244
rect 9582 18232 9588 18284
rect 9640 18272 9646 18284
rect 9784 18281 9812 18312
rect 9950 18300 9956 18352
rect 10008 18340 10014 18352
rect 10597 18343 10655 18349
rect 10597 18340 10609 18343
rect 10008 18312 10609 18340
rect 10008 18300 10014 18312
rect 10597 18309 10609 18312
rect 10643 18340 10655 18343
rect 10643 18312 11192 18340
rect 10643 18309 10655 18312
rect 10597 18303 10655 18309
rect 9677 18275 9735 18281
rect 9677 18272 9689 18275
rect 9640 18244 9689 18272
rect 9640 18232 9646 18244
rect 9677 18241 9689 18244
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 9769 18275 9827 18281
rect 9769 18241 9781 18275
rect 9815 18241 9827 18275
rect 9769 18235 9827 18241
rect 6730 18204 6736 18216
rect 6104 18176 6736 18204
rect 6730 18164 6736 18176
rect 6788 18164 6794 18216
rect 7650 18164 7656 18216
rect 7708 18204 7714 18216
rect 8021 18207 8079 18213
rect 8021 18204 8033 18207
rect 7708 18176 8033 18204
rect 7708 18164 7714 18176
rect 8021 18173 8033 18176
rect 8067 18173 8079 18207
rect 8021 18167 8079 18173
rect 8938 18164 8944 18216
rect 8996 18204 9002 18216
rect 11054 18204 11060 18216
rect 8996 18176 11060 18204
rect 8996 18164 9002 18176
rect 11054 18164 11060 18176
rect 11112 18164 11118 18216
rect 11164 18213 11192 18312
rect 11238 18232 11244 18284
rect 11296 18272 11302 18284
rect 11333 18275 11391 18281
rect 11333 18272 11345 18275
rect 11296 18244 11345 18272
rect 11296 18232 11302 18244
rect 11333 18241 11345 18244
rect 11379 18272 11391 18275
rect 11514 18272 11520 18284
rect 11379 18244 11520 18272
rect 11379 18241 11391 18244
rect 11333 18235 11391 18241
rect 11514 18232 11520 18244
rect 11572 18232 11578 18284
rect 12253 18275 12311 18281
rect 12253 18241 12265 18275
rect 12299 18272 12311 18275
rect 12618 18272 12624 18284
rect 12299 18244 12624 18272
rect 12299 18241 12311 18244
rect 12253 18235 12311 18241
rect 12618 18232 12624 18244
rect 12676 18272 12682 18284
rect 14016 18281 14044 18380
rect 14090 18368 14096 18420
rect 14148 18408 14154 18420
rect 14921 18411 14979 18417
rect 14921 18408 14933 18411
rect 14148 18380 14933 18408
rect 14148 18368 14154 18380
rect 14921 18377 14933 18380
rect 14967 18408 14979 18411
rect 15838 18408 15844 18420
rect 14967 18380 15844 18408
rect 14967 18377 14979 18380
rect 14921 18371 14979 18377
rect 12989 18275 13047 18281
rect 12989 18272 13001 18275
rect 12676 18244 13001 18272
rect 12676 18232 12682 18244
rect 12989 18241 13001 18244
rect 13035 18241 13047 18275
rect 12989 18235 13047 18241
rect 14001 18275 14059 18281
rect 14001 18241 14013 18275
rect 14047 18241 14059 18275
rect 14936 18272 14964 18371
rect 15838 18368 15844 18380
rect 15896 18408 15902 18420
rect 17037 18411 17095 18417
rect 17037 18408 17049 18411
rect 15896 18380 17049 18408
rect 15896 18368 15902 18380
rect 17037 18377 17049 18380
rect 17083 18377 17095 18411
rect 17402 18408 17408 18420
rect 17363 18380 17408 18408
rect 17037 18371 17095 18377
rect 15010 18272 15016 18284
rect 14923 18244 15016 18272
rect 14001 18235 14059 18241
rect 15010 18232 15016 18244
rect 15068 18272 15074 18284
rect 15105 18275 15163 18281
rect 15105 18272 15117 18275
rect 15068 18244 15117 18272
rect 15068 18232 15074 18244
rect 15105 18241 15117 18244
rect 15151 18241 15163 18275
rect 17052 18272 17080 18371
rect 17402 18368 17408 18380
rect 17460 18368 17466 18420
rect 18693 18411 18751 18417
rect 18693 18377 18705 18411
rect 18739 18408 18751 18411
rect 18966 18408 18972 18420
rect 18739 18380 18972 18408
rect 18739 18377 18751 18380
rect 18693 18371 18751 18377
rect 18966 18368 18972 18380
rect 19024 18408 19030 18420
rect 19426 18408 19432 18420
rect 19024 18380 19432 18408
rect 19024 18368 19030 18380
rect 19426 18368 19432 18380
rect 19484 18408 19490 18420
rect 20533 18411 20591 18417
rect 20533 18408 20545 18411
rect 19484 18380 20545 18408
rect 19484 18368 19490 18380
rect 20533 18377 20545 18380
rect 20579 18377 20591 18411
rect 21634 18408 21640 18420
rect 21595 18380 21640 18408
rect 20533 18371 20591 18377
rect 21634 18368 21640 18380
rect 21692 18368 21698 18420
rect 22738 18408 22744 18420
rect 22699 18380 22744 18408
rect 22738 18368 22744 18380
rect 22796 18368 22802 18420
rect 23014 18408 23020 18420
rect 22975 18380 23020 18408
rect 23014 18368 23020 18380
rect 23072 18368 23078 18420
rect 23661 18411 23719 18417
rect 23661 18377 23673 18411
rect 23707 18408 23719 18411
rect 24210 18408 24216 18420
rect 23707 18380 24216 18408
rect 23707 18377 23719 18380
rect 23661 18371 23719 18377
rect 24210 18368 24216 18380
rect 24268 18368 24274 18420
rect 25409 18411 25467 18417
rect 25409 18377 25421 18411
rect 25455 18408 25467 18411
rect 25498 18408 25504 18420
rect 25455 18380 25504 18408
rect 25455 18377 25467 18380
rect 25409 18371 25467 18377
rect 25498 18368 25504 18380
rect 25556 18368 25562 18420
rect 18322 18340 18328 18352
rect 18283 18312 18328 18340
rect 18322 18300 18328 18312
rect 18380 18300 18386 18352
rect 23566 18300 23572 18352
rect 23624 18340 23630 18352
rect 24394 18340 24400 18352
rect 23624 18312 24400 18340
rect 23624 18300 23630 18312
rect 24394 18300 24400 18312
rect 24452 18300 24458 18352
rect 24946 18300 24952 18352
rect 25004 18340 25010 18352
rect 25041 18343 25099 18349
rect 25041 18340 25053 18343
rect 25004 18312 25053 18340
rect 25004 18300 25010 18312
rect 25041 18309 25053 18312
rect 25087 18309 25099 18343
rect 25041 18303 25099 18309
rect 18506 18272 18512 18284
rect 17052 18244 18512 18272
rect 15105 18235 15163 18241
rect 18506 18232 18512 18244
rect 18564 18272 18570 18284
rect 18969 18275 19027 18281
rect 18969 18272 18981 18275
rect 18564 18244 18981 18272
rect 18564 18232 18570 18244
rect 18969 18241 18981 18244
rect 19015 18272 19027 18275
rect 19153 18275 19211 18281
rect 19153 18272 19165 18275
rect 19015 18244 19165 18272
rect 19015 18241 19027 18244
rect 18969 18235 19027 18241
rect 19153 18241 19165 18244
rect 19199 18241 19211 18275
rect 19153 18235 19211 18241
rect 21174 18232 21180 18284
rect 21232 18272 21238 18284
rect 21634 18272 21640 18284
rect 21232 18244 21640 18272
rect 21232 18232 21238 18244
rect 21634 18232 21640 18244
rect 21692 18272 21698 18284
rect 22189 18275 22247 18281
rect 22189 18272 22201 18275
rect 21692 18244 22201 18272
rect 21692 18232 21698 18244
rect 22189 18241 22201 18244
rect 22235 18241 22247 18275
rect 22189 18235 22247 18241
rect 24026 18232 24032 18284
rect 24084 18272 24090 18284
rect 24213 18275 24271 18281
rect 24213 18272 24225 18275
rect 24084 18244 24225 18272
rect 24084 18232 24090 18244
rect 24213 18241 24225 18244
rect 24259 18272 24271 18275
rect 24673 18275 24731 18281
rect 24673 18272 24685 18275
rect 24259 18244 24685 18272
rect 24259 18241 24271 18244
rect 24213 18235 24271 18241
rect 24673 18241 24685 18244
rect 24719 18241 24731 18275
rect 24673 18235 24731 18241
rect 11149 18207 11207 18213
rect 11149 18173 11161 18207
rect 11195 18204 11207 18207
rect 11606 18204 11612 18216
rect 11195 18176 11612 18204
rect 11195 18173 11207 18176
rect 11149 18167 11207 18173
rect 11606 18164 11612 18176
rect 11664 18164 11670 18216
rect 12805 18207 12863 18213
rect 12805 18173 12817 18207
rect 12851 18204 12863 18207
rect 13078 18204 13084 18216
rect 12851 18176 13084 18204
rect 12851 18173 12863 18176
rect 12805 18167 12863 18173
rect 13078 18164 13084 18176
rect 13136 18204 13142 18216
rect 13722 18204 13728 18216
rect 13136 18176 13728 18204
rect 13136 18164 13142 18176
rect 13722 18164 13728 18176
rect 13780 18164 13786 18216
rect 15372 18207 15430 18213
rect 15372 18204 15384 18207
rect 15304 18176 15384 18204
rect 2216 18139 2274 18145
rect 2216 18105 2228 18139
rect 2262 18136 2274 18139
rect 3602 18136 3608 18148
rect 2262 18108 3608 18136
rect 2262 18105 2274 18108
rect 2216 18099 2274 18105
rect 3602 18096 3608 18108
rect 3660 18096 3666 18148
rect 5442 18096 5448 18148
rect 5500 18136 5506 18148
rect 5537 18139 5595 18145
rect 5537 18136 5549 18139
rect 5500 18108 5549 18136
rect 5500 18096 5506 18108
rect 5537 18105 5549 18108
rect 5583 18136 5595 18139
rect 7834 18136 7840 18148
rect 5583 18108 7840 18136
rect 5583 18105 5595 18108
rect 5537 18099 5595 18105
rect 7834 18096 7840 18108
rect 7892 18096 7898 18148
rect 9398 18096 9404 18148
rect 9456 18136 9462 18148
rect 9585 18139 9643 18145
rect 9585 18136 9597 18139
rect 9456 18108 9597 18136
rect 9456 18096 9462 18108
rect 9585 18105 9597 18108
rect 9631 18136 9643 18139
rect 13998 18136 14004 18148
rect 9631 18108 10824 18136
rect 9631 18105 9643 18108
rect 9585 18099 9643 18105
rect 3326 18068 3332 18080
rect 3287 18040 3332 18068
rect 3326 18028 3332 18040
rect 3384 18028 3390 18080
rect 5166 18068 5172 18080
rect 5127 18040 5172 18068
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 5626 18068 5632 18080
rect 5587 18040 5632 18068
rect 5626 18028 5632 18040
rect 5684 18028 5690 18080
rect 7466 18068 7472 18080
rect 7427 18040 7472 18068
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 7650 18068 7656 18080
rect 7611 18040 7656 18068
rect 7650 18028 7656 18040
rect 7708 18028 7714 18080
rect 8757 18071 8815 18077
rect 8757 18037 8769 18071
rect 8803 18068 8815 18071
rect 8846 18068 8852 18080
rect 8803 18040 8852 18068
rect 8803 18037 8815 18040
rect 8757 18031 8815 18037
rect 8846 18028 8852 18040
rect 8904 18028 8910 18080
rect 10796 18077 10824 18108
rect 12820 18108 14004 18136
rect 10781 18071 10839 18077
rect 10781 18037 10793 18071
rect 10827 18037 10839 18071
rect 11238 18068 11244 18080
rect 11199 18040 11244 18068
rect 10781 18031 10839 18037
rect 11238 18028 11244 18040
rect 11296 18028 11302 18080
rect 11330 18028 11336 18080
rect 11388 18068 11394 18080
rect 11793 18071 11851 18077
rect 11793 18068 11805 18071
rect 11388 18040 11805 18068
rect 11388 18028 11394 18040
rect 11793 18037 11805 18040
rect 11839 18037 11851 18071
rect 11793 18031 11851 18037
rect 12437 18071 12495 18077
rect 12437 18037 12449 18071
rect 12483 18068 12495 18071
rect 12820 18068 12848 18108
rect 13998 18096 14004 18108
rect 14056 18096 14062 18148
rect 14645 18139 14703 18145
rect 14645 18105 14657 18139
rect 14691 18136 14703 18139
rect 15304 18136 15332 18176
rect 15372 18173 15384 18176
rect 15418 18204 15430 18207
rect 15654 18204 15660 18216
rect 15418 18176 15660 18204
rect 15418 18173 15430 18176
rect 15372 18167 15430 18173
rect 15654 18164 15660 18176
rect 15712 18164 15718 18216
rect 17865 18207 17923 18213
rect 17865 18173 17877 18207
rect 17911 18204 17923 18207
rect 18138 18204 18144 18216
rect 17911 18176 18144 18204
rect 17911 18173 17923 18176
rect 17865 18167 17923 18173
rect 18138 18164 18144 18176
rect 18196 18164 18202 18216
rect 19242 18164 19248 18216
rect 19300 18204 19306 18216
rect 19420 18207 19478 18213
rect 19420 18204 19432 18207
rect 19300 18176 19432 18204
rect 19300 18164 19306 18176
rect 19420 18173 19432 18176
rect 19466 18204 19478 18207
rect 21192 18204 21220 18232
rect 19466 18176 21220 18204
rect 19466 18173 19478 18176
rect 19420 18167 19478 18173
rect 23014 18164 23020 18216
rect 23072 18204 23078 18216
rect 24118 18204 24124 18216
rect 23072 18176 24124 18204
rect 23072 18164 23078 18176
rect 24118 18164 24124 18176
rect 24176 18164 24182 18216
rect 24854 18164 24860 18216
rect 24912 18204 24918 18216
rect 25225 18207 25283 18213
rect 25225 18204 25237 18207
rect 24912 18176 25237 18204
rect 24912 18164 24918 18176
rect 25225 18173 25237 18176
rect 25271 18204 25283 18207
rect 25777 18207 25835 18213
rect 25777 18204 25789 18207
rect 25271 18176 25789 18204
rect 25271 18173 25283 18176
rect 25225 18167 25283 18173
rect 25777 18173 25789 18176
rect 25823 18173 25835 18207
rect 25777 18167 25835 18173
rect 14691 18108 15332 18136
rect 14691 18105 14703 18108
rect 14645 18099 14703 18105
rect 17310 18096 17316 18148
rect 17368 18136 17374 18148
rect 20990 18136 20996 18148
rect 17368 18108 20996 18136
rect 17368 18096 17374 18108
rect 20990 18096 20996 18108
rect 21048 18136 21054 18148
rect 21085 18139 21143 18145
rect 21085 18136 21097 18139
rect 21048 18108 21097 18136
rect 21048 18096 21054 18108
rect 21085 18105 21097 18108
rect 21131 18105 21143 18139
rect 21085 18099 21143 18105
rect 21545 18139 21603 18145
rect 21545 18105 21557 18139
rect 21591 18136 21603 18139
rect 22097 18139 22155 18145
rect 22097 18136 22109 18139
rect 21591 18108 22109 18136
rect 21591 18105 21603 18108
rect 21545 18099 21603 18105
rect 22097 18105 22109 18108
rect 22143 18136 22155 18139
rect 22186 18136 22192 18148
rect 22143 18108 22192 18136
rect 22143 18105 22155 18108
rect 22097 18099 22155 18105
rect 12483 18040 12848 18068
rect 12897 18071 12955 18077
rect 12483 18037 12495 18040
rect 12437 18031 12495 18037
rect 12897 18037 12909 18071
rect 12943 18068 12955 18071
rect 13078 18068 13084 18080
rect 12943 18040 13084 18068
rect 12943 18037 12955 18040
rect 12897 18031 12955 18037
rect 13078 18028 13084 18040
rect 13136 18028 13142 18080
rect 16482 18068 16488 18080
rect 16443 18040 16488 18068
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 20898 18028 20904 18080
rect 20956 18068 20962 18080
rect 21560 18068 21588 18099
rect 22186 18096 22192 18108
rect 22244 18096 22250 18148
rect 23477 18139 23535 18145
rect 23477 18105 23489 18139
rect 23523 18136 23535 18139
rect 24029 18139 24087 18145
rect 24029 18136 24041 18139
rect 23523 18108 24041 18136
rect 23523 18105 23535 18108
rect 23477 18099 23535 18105
rect 24029 18105 24041 18108
rect 24075 18136 24087 18139
rect 24670 18136 24676 18148
rect 24075 18108 24676 18136
rect 24075 18105 24087 18108
rect 24029 18099 24087 18105
rect 24136 18080 24164 18108
rect 24670 18096 24676 18108
rect 24728 18096 24734 18148
rect 22002 18068 22008 18080
rect 20956 18040 21588 18068
rect 21963 18040 22008 18068
rect 20956 18028 20962 18040
rect 22002 18028 22008 18040
rect 22060 18068 22066 18080
rect 22370 18068 22376 18080
rect 22060 18040 22376 18068
rect 22060 18028 22066 18040
rect 22370 18028 22376 18040
rect 22428 18028 22434 18080
rect 24118 18028 24124 18080
rect 24176 18028 24182 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1578 17864 1584 17876
rect 1539 17836 1584 17864
rect 1578 17824 1584 17836
rect 1636 17824 1642 17876
rect 2317 17867 2375 17873
rect 2317 17833 2329 17867
rect 2363 17864 2375 17867
rect 2590 17864 2596 17876
rect 2363 17836 2596 17864
rect 2363 17833 2375 17836
rect 2317 17827 2375 17833
rect 2590 17824 2596 17836
rect 2648 17824 2654 17876
rect 4893 17867 4951 17873
rect 4893 17833 4905 17867
rect 4939 17864 4951 17867
rect 5442 17864 5448 17876
rect 4939 17836 5448 17864
rect 4939 17833 4951 17836
rect 4893 17827 4951 17833
rect 5442 17824 5448 17836
rect 5500 17824 5506 17876
rect 7650 17864 7656 17876
rect 5552 17836 7656 17864
rect 2774 17756 2780 17808
rect 2832 17796 2838 17808
rect 3418 17796 3424 17808
rect 2832 17768 3424 17796
rect 2832 17756 2838 17768
rect 3418 17756 3424 17768
rect 3476 17756 3482 17808
rect 3513 17799 3571 17805
rect 3513 17765 3525 17799
rect 3559 17796 3571 17799
rect 3602 17796 3608 17808
rect 3559 17768 3608 17796
rect 3559 17765 3571 17768
rect 3513 17759 3571 17765
rect 3602 17756 3608 17768
rect 3660 17756 3666 17808
rect 3881 17799 3939 17805
rect 3881 17765 3893 17799
rect 3927 17796 3939 17799
rect 5552 17796 5580 17836
rect 7650 17824 7656 17836
rect 7708 17824 7714 17876
rect 7745 17867 7803 17873
rect 7745 17833 7757 17867
rect 7791 17864 7803 17867
rect 8202 17864 8208 17876
rect 7791 17836 8208 17864
rect 7791 17833 7803 17836
rect 7745 17827 7803 17833
rect 8202 17824 8208 17836
rect 8260 17824 8266 17876
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 10045 17867 10103 17873
rect 10045 17864 10057 17867
rect 9732 17836 10057 17864
rect 9732 17824 9738 17836
rect 10045 17833 10057 17836
rect 10091 17833 10103 17867
rect 10870 17864 10876 17876
rect 10831 17836 10876 17864
rect 10045 17827 10103 17833
rect 10870 17824 10876 17836
rect 10928 17824 10934 17876
rect 11146 17864 11152 17876
rect 11107 17836 11152 17864
rect 11146 17824 11152 17836
rect 11204 17824 11210 17876
rect 11514 17864 11520 17876
rect 11475 17836 11520 17864
rect 11514 17824 11520 17836
rect 11572 17824 11578 17876
rect 12069 17867 12127 17873
rect 12069 17833 12081 17867
rect 12115 17864 12127 17867
rect 12621 17867 12679 17873
rect 12621 17864 12633 17867
rect 12115 17836 12633 17864
rect 12115 17833 12127 17836
rect 12069 17827 12127 17833
rect 12621 17833 12633 17836
rect 12667 17864 12679 17867
rect 12986 17864 12992 17876
rect 12667 17836 12992 17864
rect 12667 17833 12679 17836
rect 12621 17827 12679 17833
rect 12986 17824 12992 17836
rect 13044 17824 13050 17876
rect 13446 17864 13452 17876
rect 13407 17836 13452 17864
rect 13446 17824 13452 17836
rect 13504 17824 13510 17876
rect 13814 17824 13820 17876
rect 13872 17864 13878 17876
rect 14553 17867 14611 17873
rect 14553 17864 14565 17867
rect 13872 17836 14565 17864
rect 13872 17824 13878 17836
rect 14553 17833 14565 17836
rect 14599 17833 14611 17867
rect 15102 17864 15108 17876
rect 15063 17836 15108 17864
rect 14553 17827 14611 17833
rect 15102 17824 15108 17836
rect 15160 17824 15166 17876
rect 15746 17824 15752 17876
rect 15804 17864 15810 17876
rect 16390 17864 16396 17876
rect 15804 17836 16396 17864
rect 15804 17824 15810 17836
rect 16390 17824 16396 17836
rect 16448 17824 16454 17876
rect 18230 17864 18236 17876
rect 18191 17836 18236 17864
rect 18230 17824 18236 17836
rect 18288 17824 18294 17876
rect 18782 17864 18788 17876
rect 18743 17836 18788 17864
rect 18782 17824 18788 17836
rect 18840 17824 18846 17876
rect 19242 17864 19248 17876
rect 19203 17836 19248 17864
rect 19242 17824 19248 17836
rect 19300 17824 19306 17876
rect 19978 17824 19984 17876
rect 20036 17864 20042 17876
rect 20257 17867 20315 17873
rect 20257 17864 20269 17867
rect 20036 17836 20269 17864
rect 20036 17824 20042 17836
rect 20257 17833 20269 17836
rect 20303 17833 20315 17867
rect 20257 17827 20315 17833
rect 20717 17867 20775 17873
rect 20717 17833 20729 17867
rect 20763 17864 20775 17867
rect 21450 17864 21456 17876
rect 20763 17836 21456 17864
rect 20763 17833 20775 17836
rect 20717 17827 20775 17833
rect 21450 17824 21456 17836
rect 21508 17824 21514 17876
rect 22554 17864 22560 17876
rect 22515 17836 22560 17864
rect 22554 17824 22560 17836
rect 22612 17824 22618 17876
rect 23106 17824 23112 17876
rect 23164 17864 23170 17876
rect 23290 17864 23296 17876
rect 23164 17836 23296 17864
rect 23164 17824 23170 17836
rect 23290 17824 23296 17836
rect 23348 17824 23354 17876
rect 24121 17867 24179 17873
rect 24121 17833 24133 17867
rect 24167 17864 24179 17867
rect 24210 17864 24216 17876
rect 24167 17836 24216 17864
rect 24167 17833 24179 17836
rect 24121 17827 24179 17833
rect 24210 17824 24216 17836
rect 24268 17864 24274 17876
rect 24394 17864 24400 17876
rect 24268 17836 24400 17864
rect 24268 17824 24274 17836
rect 24394 17824 24400 17836
rect 24452 17824 24458 17876
rect 25406 17864 25412 17876
rect 25367 17836 25412 17864
rect 25406 17824 25412 17836
rect 25464 17824 25470 17876
rect 6822 17796 6828 17808
rect 3927 17768 5580 17796
rect 6735 17768 6828 17796
rect 3927 17765 3939 17768
rect 3881 17759 3939 17765
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17697 1455 17731
rect 3050 17728 3056 17740
rect 1397 17691 1455 17697
rect 2884 17700 3056 17728
rect 1412 17660 1440 17691
rect 2884 17672 2912 17700
rect 3050 17688 3056 17700
rect 3108 17688 3114 17740
rect 2866 17660 2872 17672
rect 1412 17632 2636 17660
rect 2827 17632 2872 17660
rect 1949 17595 2007 17601
rect 1949 17561 1961 17595
rect 1995 17592 2007 17595
rect 2498 17592 2504 17604
rect 1995 17564 2504 17592
rect 1995 17561 2007 17564
rect 1949 17555 2007 17561
rect 2498 17552 2504 17564
rect 2556 17552 2562 17604
rect 2314 17484 2320 17536
rect 2372 17524 2378 17536
rect 2409 17527 2467 17533
rect 2409 17524 2421 17527
rect 2372 17496 2421 17524
rect 2372 17484 2378 17496
rect 2409 17493 2421 17496
rect 2455 17493 2467 17527
rect 2608 17524 2636 17632
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 2961 17663 3019 17669
rect 2961 17629 2973 17663
rect 3007 17660 3019 17663
rect 3234 17660 3240 17672
rect 3007 17632 3240 17660
rect 3007 17629 3019 17632
rect 2961 17623 3019 17629
rect 3234 17620 3240 17632
rect 3292 17620 3298 17672
rect 3896 17524 3924 17759
rect 6822 17756 6828 17768
rect 6880 17796 6886 17808
rect 8938 17796 8944 17808
rect 6880 17768 8944 17796
rect 6880 17756 6886 17768
rect 8938 17756 8944 17768
rect 8996 17756 9002 17808
rect 14182 17796 14188 17808
rect 14143 17768 14188 17796
rect 14182 17756 14188 17768
rect 14240 17756 14246 17808
rect 15286 17756 15292 17808
rect 15344 17796 15350 17808
rect 15556 17799 15614 17805
rect 15556 17796 15568 17799
rect 15344 17768 15568 17796
rect 15344 17756 15350 17768
rect 15556 17765 15568 17768
rect 15602 17796 15614 17799
rect 16482 17796 16488 17808
rect 15602 17768 16488 17796
rect 15602 17765 15614 17768
rect 15556 17759 15614 17765
rect 16482 17756 16488 17768
rect 16540 17756 16546 17808
rect 22002 17796 22008 17808
rect 18156 17768 22008 17796
rect 4801 17731 4859 17737
rect 4801 17697 4813 17731
rect 4847 17728 4859 17731
rect 4982 17728 4988 17740
rect 4847 17700 4988 17728
rect 4847 17697 4859 17700
rect 4801 17691 4859 17697
rect 4982 17688 4988 17700
rect 5040 17728 5046 17740
rect 5261 17731 5319 17737
rect 5261 17728 5273 17731
rect 5040 17700 5273 17728
rect 5040 17688 5046 17700
rect 5261 17697 5273 17700
rect 5307 17697 5319 17731
rect 5261 17691 5319 17697
rect 6273 17731 6331 17737
rect 6273 17697 6285 17731
rect 6319 17728 6331 17731
rect 6319 17700 7236 17728
rect 6319 17697 6331 17700
rect 6273 17691 6331 17697
rect 5074 17620 5080 17672
rect 5132 17660 5138 17672
rect 5353 17663 5411 17669
rect 5353 17660 5365 17663
rect 5132 17632 5365 17660
rect 5132 17620 5138 17632
rect 5353 17629 5365 17632
rect 5399 17629 5411 17663
rect 5353 17623 5411 17629
rect 5445 17663 5503 17669
rect 5445 17629 5457 17663
rect 5491 17629 5503 17663
rect 6914 17660 6920 17672
rect 6875 17632 6920 17660
rect 5445 17623 5503 17629
rect 4433 17595 4491 17601
rect 4433 17561 4445 17595
rect 4479 17592 4491 17595
rect 5460 17592 5488 17623
rect 6914 17620 6920 17632
rect 6972 17620 6978 17672
rect 7009 17663 7067 17669
rect 7009 17629 7021 17663
rect 7055 17629 7067 17663
rect 7208 17660 7236 17700
rect 8294 17688 8300 17740
rect 8352 17728 8358 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 8352 17700 8401 17728
rect 8352 17688 8358 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 12529 17731 12587 17737
rect 12529 17697 12541 17731
rect 12575 17728 12587 17731
rect 12894 17728 12900 17740
rect 12575 17700 12900 17728
rect 12575 17697 12587 17700
rect 12529 17691 12587 17697
rect 12894 17688 12900 17700
rect 12952 17688 12958 17740
rect 13630 17688 13636 17740
rect 13688 17728 13694 17740
rect 13725 17731 13783 17737
rect 13725 17728 13737 17731
rect 13688 17700 13737 17728
rect 13688 17688 13694 17700
rect 13725 17697 13737 17700
rect 13771 17697 13783 17731
rect 13725 17691 13783 17697
rect 17494 17688 17500 17740
rect 17552 17728 17558 17740
rect 18156 17737 18184 17768
rect 22002 17756 22008 17768
rect 22060 17756 22066 17808
rect 22646 17756 22652 17808
rect 22704 17796 22710 17808
rect 22986 17799 23044 17805
rect 22986 17796 22998 17799
rect 22704 17768 22998 17796
rect 22704 17756 22710 17768
rect 22986 17765 22998 17768
rect 23032 17765 23044 17799
rect 22986 17759 23044 17765
rect 18141 17731 18199 17737
rect 18141 17728 18153 17731
rect 17552 17700 18153 17728
rect 17552 17688 17558 17700
rect 18141 17697 18153 17700
rect 18187 17697 18199 17731
rect 18141 17691 18199 17697
rect 19242 17688 19248 17740
rect 19300 17728 19306 17740
rect 19797 17731 19855 17737
rect 19797 17728 19809 17731
rect 19300 17700 19809 17728
rect 19300 17688 19306 17700
rect 19797 17697 19809 17700
rect 19843 17697 19855 17731
rect 19797 17691 19855 17697
rect 21174 17688 21180 17740
rect 21232 17728 21238 17740
rect 21269 17731 21327 17737
rect 21269 17728 21281 17731
rect 21232 17700 21281 17728
rect 21232 17688 21238 17700
rect 21269 17697 21281 17700
rect 21315 17697 21327 17731
rect 21269 17691 21327 17697
rect 21361 17731 21419 17737
rect 21361 17697 21373 17731
rect 21407 17728 21419 17731
rect 21910 17728 21916 17740
rect 21407 17700 21916 17728
rect 21407 17697 21419 17700
rect 21361 17691 21419 17697
rect 21910 17688 21916 17700
rect 21968 17688 21974 17740
rect 22738 17728 22744 17740
rect 22699 17700 22744 17728
rect 22738 17688 22744 17700
rect 22796 17688 22802 17740
rect 24946 17688 24952 17740
rect 25004 17728 25010 17740
rect 25225 17731 25283 17737
rect 25225 17728 25237 17731
rect 25004 17700 25237 17728
rect 25004 17688 25010 17700
rect 25225 17697 25237 17700
rect 25271 17697 25283 17731
rect 25225 17691 25283 17697
rect 8478 17660 8484 17672
rect 7208 17632 8484 17660
rect 7009 17623 7067 17629
rect 5534 17592 5540 17604
rect 4479 17564 5540 17592
rect 4479 17561 4491 17564
rect 4433 17555 4491 17561
rect 5534 17552 5540 17564
rect 5592 17592 5598 17604
rect 5905 17595 5963 17601
rect 5905 17592 5917 17595
rect 5592 17564 5917 17592
rect 5592 17552 5598 17564
rect 5905 17561 5917 17564
rect 5951 17592 5963 17595
rect 7024 17592 7052 17623
rect 8478 17620 8484 17632
rect 8536 17620 8542 17672
rect 8570 17620 8576 17672
rect 8628 17660 8634 17672
rect 10137 17663 10195 17669
rect 8628 17632 8673 17660
rect 8628 17620 8634 17632
rect 10137 17629 10149 17663
rect 10183 17629 10195 17663
rect 10137 17623 10195 17629
rect 10321 17663 10379 17669
rect 10321 17629 10333 17663
rect 10367 17660 10379 17663
rect 11146 17660 11152 17672
rect 10367 17632 11152 17660
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 5951 17564 7052 17592
rect 5951 17561 5963 17564
rect 5905 17555 5963 17561
rect 8754 17552 8760 17604
rect 8812 17592 8818 17604
rect 9125 17595 9183 17601
rect 9125 17592 9137 17595
rect 8812 17564 9137 17592
rect 8812 17552 8818 17564
rect 9125 17561 9137 17564
rect 9171 17592 9183 17595
rect 9677 17595 9735 17601
rect 9677 17592 9689 17595
rect 9171 17564 9689 17592
rect 9171 17561 9183 17564
rect 9125 17555 9183 17561
rect 9677 17561 9689 17564
rect 9723 17561 9735 17595
rect 9677 17555 9735 17561
rect 2608 17496 3924 17524
rect 2409 17487 2467 17493
rect 4522 17484 4528 17536
rect 4580 17524 4586 17536
rect 4798 17524 4804 17536
rect 4580 17496 4804 17524
rect 4580 17484 4586 17496
rect 4798 17484 4804 17496
rect 4856 17484 4862 17536
rect 6454 17524 6460 17536
rect 6415 17496 6460 17524
rect 6454 17484 6460 17496
rect 6512 17484 6518 17536
rect 8018 17524 8024 17536
rect 7979 17496 8024 17524
rect 8018 17484 8024 17496
rect 8076 17484 8082 17536
rect 9398 17524 9404 17536
rect 9359 17496 9404 17524
rect 9398 17484 9404 17496
rect 9456 17524 9462 17536
rect 10152 17524 10180 17623
rect 11146 17620 11152 17632
rect 11204 17620 11210 17672
rect 12805 17663 12863 17669
rect 12805 17629 12817 17663
rect 12851 17660 12863 17663
rect 13446 17660 13452 17672
rect 12851 17632 13452 17660
rect 12851 17629 12863 17632
rect 12805 17623 12863 17629
rect 13446 17620 13452 17632
rect 13504 17620 13510 17672
rect 15010 17620 15016 17672
rect 15068 17660 15074 17672
rect 15289 17663 15347 17669
rect 15289 17660 15301 17663
rect 15068 17632 15301 17660
rect 15068 17620 15074 17632
rect 15289 17629 15301 17632
rect 15335 17629 15347 17663
rect 15289 17623 15347 17629
rect 18417 17663 18475 17669
rect 18417 17629 18429 17663
rect 18463 17660 18475 17663
rect 18598 17660 18604 17672
rect 18463 17632 18604 17660
rect 18463 17629 18475 17632
rect 18417 17623 18475 17629
rect 13906 17592 13912 17604
rect 13867 17564 13912 17592
rect 13906 17552 13912 17564
rect 13964 17552 13970 17604
rect 9456 17496 10180 17524
rect 12161 17527 12219 17533
rect 9456 17484 9462 17496
rect 12161 17493 12173 17527
rect 12207 17524 12219 17527
rect 12342 17524 12348 17536
rect 12207 17496 12348 17524
rect 12207 17493 12219 17496
rect 12161 17487 12219 17493
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 15304 17524 15332 17623
rect 18598 17620 18604 17632
rect 18656 17620 18662 17672
rect 20070 17620 20076 17672
rect 20128 17660 20134 17672
rect 20346 17660 20352 17672
rect 20128 17632 20352 17660
rect 20128 17620 20134 17632
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 21450 17660 21456 17672
rect 21411 17632 21456 17660
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 16758 17552 16764 17604
rect 16816 17592 16822 17604
rect 17313 17595 17371 17601
rect 17313 17592 17325 17595
rect 16816 17564 17325 17592
rect 16816 17552 16822 17564
rect 17313 17561 17325 17564
rect 17359 17592 17371 17595
rect 17773 17595 17831 17601
rect 17773 17592 17785 17595
rect 17359 17564 17785 17592
rect 17359 17561 17371 17564
rect 17313 17555 17371 17561
rect 17773 17561 17785 17564
rect 17819 17561 17831 17595
rect 17773 17555 17831 17561
rect 19426 17552 19432 17604
rect 19484 17592 19490 17604
rect 20901 17595 20959 17601
rect 20901 17592 20913 17595
rect 19484 17564 20913 17592
rect 19484 17552 19490 17564
rect 20901 17561 20913 17564
rect 20947 17561 20959 17595
rect 20901 17555 20959 17561
rect 15654 17524 15660 17536
rect 15304 17496 15660 17524
rect 15654 17484 15660 17496
rect 15712 17484 15718 17536
rect 16666 17524 16672 17536
rect 16627 17496 16672 17524
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 17586 17524 17592 17536
rect 17547 17496 17592 17524
rect 17586 17484 17592 17496
rect 17644 17484 17650 17536
rect 19702 17524 19708 17536
rect 19663 17496 19708 17524
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 19978 17524 19984 17536
rect 19939 17496 19984 17524
rect 19978 17484 19984 17496
rect 20036 17484 20042 17536
rect 20438 17484 20444 17536
rect 20496 17524 20502 17536
rect 20622 17524 20628 17536
rect 20496 17496 20628 17524
rect 20496 17484 20502 17496
rect 20622 17484 20628 17496
rect 20680 17484 20686 17536
rect 24670 17524 24676 17536
rect 24631 17496 24676 17524
rect 24670 17484 24676 17496
rect 24728 17484 24734 17536
rect 24854 17484 24860 17536
rect 24912 17524 24918 17536
rect 25041 17527 25099 17533
rect 25041 17524 25053 17527
rect 24912 17496 25053 17524
rect 24912 17484 24918 17496
rect 25041 17493 25053 17496
rect 25087 17493 25099 17527
rect 25041 17487 25099 17493
rect 25406 17484 25412 17536
rect 25464 17524 25470 17536
rect 25958 17524 25964 17536
rect 25464 17496 25964 17524
rect 25464 17484 25470 17496
rect 25958 17484 25964 17496
rect 26016 17484 26022 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1949 17323 2007 17329
rect 1949 17289 1961 17323
rect 1995 17320 2007 17323
rect 2774 17320 2780 17332
rect 1995 17292 2780 17320
rect 1995 17289 2007 17292
rect 1949 17283 2007 17289
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 3786 17280 3792 17332
rect 3844 17320 3850 17332
rect 4249 17323 4307 17329
rect 4249 17320 4261 17323
rect 3844 17292 4261 17320
rect 3844 17280 3850 17292
rect 4249 17289 4261 17292
rect 4295 17320 4307 17323
rect 5074 17320 5080 17332
rect 4295 17292 5080 17320
rect 4295 17289 4307 17292
rect 4249 17283 4307 17289
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 5169 17323 5227 17329
rect 5169 17289 5181 17323
rect 5215 17320 5227 17323
rect 5442 17320 5448 17332
rect 5215 17292 5448 17320
rect 5215 17289 5227 17292
rect 5169 17283 5227 17289
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 6549 17323 6607 17329
rect 6549 17289 6561 17323
rect 6595 17320 6607 17323
rect 6822 17320 6828 17332
rect 6595 17292 6828 17320
rect 6595 17289 6607 17292
rect 6549 17283 6607 17289
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 8113 17323 8171 17329
rect 8113 17289 8125 17323
rect 8159 17320 8171 17323
rect 8570 17320 8576 17332
rect 8159 17292 8576 17320
rect 8159 17289 8171 17292
rect 8113 17283 8171 17289
rect 8570 17280 8576 17292
rect 8628 17280 8634 17332
rect 9401 17323 9459 17329
rect 9401 17289 9413 17323
rect 9447 17320 9459 17323
rect 11146 17320 11152 17332
rect 9447 17292 11152 17320
rect 9447 17289 9459 17292
rect 9401 17283 9459 17289
rect 11146 17280 11152 17292
rect 11204 17320 11210 17332
rect 11885 17323 11943 17329
rect 11885 17320 11897 17323
rect 11204 17292 11897 17320
rect 11204 17280 11210 17292
rect 11885 17289 11897 17292
rect 11931 17320 11943 17323
rect 13446 17320 13452 17332
rect 11931 17292 13452 17320
rect 11931 17289 11943 17292
rect 11885 17283 11943 17289
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 15286 17320 15292 17332
rect 15247 17292 15292 17320
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 15654 17280 15660 17332
rect 15712 17320 15718 17332
rect 15841 17323 15899 17329
rect 15841 17320 15853 17323
rect 15712 17292 15853 17320
rect 15712 17280 15718 17292
rect 15841 17289 15853 17292
rect 15887 17289 15899 17323
rect 17494 17320 17500 17332
rect 17455 17292 17500 17320
rect 15841 17283 15899 17289
rect 17494 17280 17500 17292
rect 17552 17280 17558 17332
rect 17865 17323 17923 17329
rect 17865 17289 17877 17323
rect 17911 17320 17923 17323
rect 18230 17320 18236 17332
rect 17911 17292 18236 17320
rect 17911 17289 17923 17292
rect 17865 17283 17923 17289
rect 18230 17280 18236 17292
rect 18288 17280 18294 17332
rect 19150 17320 19156 17332
rect 19111 17292 19156 17320
rect 19150 17280 19156 17292
rect 19208 17280 19214 17332
rect 21358 17280 21364 17332
rect 21416 17280 21422 17332
rect 21634 17320 21640 17332
rect 21595 17292 21640 17320
rect 21634 17280 21640 17292
rect 21692 17280 21698 17332
rect 22373 17323 22431 17329
rect 22373 17289 22385 17323
rect 22419 17320 22431 17323
rect 22646 17320 22652 17332
rect 22419 17292 22652 17320
rect 22419 17289 22431 17292
rect 22373 17283 22431 17289
rect 22646 17280 22652 17292
rect 22704 17280 22710 17332
rect 22738 17280 22744 17332
rect 22796 17320 22802 17332
rect 23017 17323 23075 17329
rect 23017 17320 23029 17323
rect 22796 17292 23029 17320
rect 22796 17280 22802 17292
rect 23017 17289 23029 17292
rect 23063 17289 23075 17323
rect 23474 17320 23480 17332
rect 23435 17292 23480 17320
rect 23017 17283 23075 17289
rect 23474 17280 23480 17292
rect 23532 17280 23538 17332
rect 23658 17320 23664 17332
rect 23619 17292 23664 17320
rect 23658 17280 23664 17292
rect 23716 17280 23722 17332
rect 25409 17323 25467 17329
rect 25409 17289 25421 17323
rect 25455 17320 25467 17323
rect 25774 17320 25780 17332
rect 25455 17292 25780 17320
rect 25455 17289 25467 17292
rect 25409 17283 25467 17289
rect 25774 17280 25780 17292
rect 25832 17280 25838 17332
rect 25869 17323 25927 17329
rect 25869 17289 25881 17323
rect 25915 17320 25927 17323
rect 26142 17320 26148 17332
rect 25915 17292 26148 17320
rect 25915 17289 25927 17292
rect 25869 17283 25927 17289
rect 1578 17212 1584 17264
rect 1636 17252 1642 17264
rect 1854 17252 1860 17264
rect 1636 17224 1860 17252
rect 1636 17212 1642 17224
rect 1854 17212 1860 17224
rect 1912 17212 1918 17264
rect 3878 17212 3884 17264
rect 3936 17252 3942 17264
rect 4338 17252 4344 17264
rect 3936 17224 4344 17252
rect 3936 17212 3942 17224
rect 4338 17212 4344 17224
rect 4396 17252 4402 17264
rect 4617 17255 4675 17261
rect 4617 17252 4629 17255
rect 4396 17224 4629 17252
rect 4396 17212 4402 17224
rect 4617 17221 4629 17224
rect 4663 17221 4675 17255
rect 9674 17252 9680 17264
rect 9635 17224 9680 17252
rect 4617 17215 4675 17221
rect 1302 17144 1308 17196
rect 1360 17184 1366 17196
rect 1486 17184 1492 17196
rect 1360 17156 1492 17184
rect 1360 17144 1366 17156
rect 1486 17144 1492 17156
rect 1544 17144 1550 17196
rect 1946 17144 1952 17196
rect 2004 17144 2010 17196
rect 1964 17116 1992 17144
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1964 17088 2053 17116
rect 2041 17085 2053 17088
rect 2087 17116 2099 17119
rect 2130 17116 2136 17128
rect 2087 17088 2136 17116
rect 2087 17085 2099 17088
rect 2041 17079 2099 17085
rect 2130 17076 2136 17088
rect 2188 17076 2194 17128
rect 1854 17008 1860 17060
rect 1912 17048 1918 17060
rect 2308 17051 2366 17057
rect 2308 17048 2320 17051
rect 1912 17020 2320 17048
rect 1912 17008 1918 17020
rect 2308 17017 2320 17020
rect 2354 17048 2366 17051
rect 3326 17048 3332 17060
rect 2354 17020 3332 17048
rect 2354 17017 2366 17020
rect 2308 17011 2366 17017
rect 3326 17008 3332 17020
rect 3384 17048 3390 17060
rect 3786 17048 3792 17060
rect 3384 17020 3792 17048
rect 3384 17008 3390 17020
rect 3786 17008 3792 17020
rect 3844 17008 3850 17060
rect 4632 17048 4660 17215
rect 9674 17212 9680 17224
rect 9732 17212 9738 17264
rect 11238 17252 11244 17264
rect 11199 17224 11244 17252
rect 11238 17212 11244 17224
rect 11296 17212 11302 17264
rect 4982 17144 4988 17196
rect 5040 17184 5046 17196
rect 5442 17184 5448 17196
rect 5040 17156 5448 17184
rect 5040 17144 5046 17156
rect 5442 17144 5448 17156
rect 5500 17144 5506 17196
rect 5534 17144 5540 17196
rect 5592 17184 5598 17196
rect 5721 17187 5779 17193
rect 5721 17184 5733 17187
rect 5592 17156 5733 17184
rect 5592 17144 5598 17156
rect 5721 17153 5733 17156
rect 5767 17153 5779 17187
rect 8754 17184 8760 17196
rect 8715 17156 8760 17184
rect 5721 17147 5779 17153
rect 8754 17144 8760 17156
rect 8812 17144 8818 17196
rect 8941 17187 8999 17193
rect 8941 17153 8953 17187
rect 8987 17184 8999 17187
rect 9490 17184 9496 17196
rect 8987 17156 9496 17184
rect 8987 17153 8999 17156
rect 8941 17147 8999 17153
rect 9490 17144 9496 17156
rect 9548 17144 9554 17196
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 12161 17187 12219 17193
rect 12161 17184 12173 17187
rect 11112 17156 12173 17184
rect 11112 17144 11118 17156
rect 12161 17153 12173 17156
rect 12207 17184 12219 17187
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12207 17156 12449 17184
rect 12207 17153 12219 17156
rect 12161 17147 12219 17153
rect 12437 17153 12449 17156
rect 12483 17153 12495 17187
rect 12437 17147 12495 17153
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17184 15439 17187
rect 16482 17184 16488 17196
rect 15427 17156 16488 17184
rect 15427 17153 15439 17156
rect 15381 17147 15439 17153
rect 16482 17144 16488 17156
rect 16540 17144 16546 17196
rect 16945 17187 17003 17193
rect 16945 17153 16957 17187
rect 16991 17153 17003 17187
rect 16945 17147 17003 17153
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 7377 17119 7435 17125
rect 7377 17116 7389 17119
rect 6871 17088 7389 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 7377 17085 7389 17088
rect 7423 17116 7435 17119
rect 8202 17116 8208 17128
rect 7423 17088 8208 17116
rect 7423 17085 7435 17088
rect 7377 17079 7435 17085
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 8665 17119 8723 17125
rect 8665 17085 8677 17119
rect 8711 17116 8723 17119
rect 9030 17116 9036 17128
rect 8711 17088 9036 17116
rect 8711 17085 8723 17088
rect 8665 17079 8723 17085
rect 9030 17076 9036 17088
rect 9088 17116 9094 17128
rect 9674 17116 9680 17128
rect 9088 17088 9680 17116
rect 9088 17076 9094 17088
rect 9674 17076 9680 17088
rect 9732 17076 9738 17128
rect 9861 17119 9919 17125
rect 9861 17085 9873 17119
rect 9907 17116 9919 17119
rect 9950 17116 9956 17128
rect 9907 17088 9956 17116
rect 9907 17085 9919 17088
rect 9861 17079 9919 17085
rect 9950 17076 9956 17088
rect 10008 17116 10014 17128
rect 11072 17116 11100 17144
rect 14366 17116 14372 17128
rect 10008 17088 11100 17116
rect 14327 17088 14372 17116
rect 10008 17076 10014 17088
rect 14366 17076 14372 17088
rect 14424 17076 14430 17128
rect 16758 17116 16764 17128
rect 16719 17088 16764 17116
rect 16758 17076 16764 17088
rect 16816 17076 16822 17128
rect 5537 17051 5595 17057
rect 5537 17048 5549 17051
rect 4632 17020 5549 17048
rect 5537 17017 5549 17020
rect 5583 17017 5595 17051
rect 5537 17011 5595 17017
rect 9490 17008 9496 17060
rect 9548 17048 9554 17060
rect 10128 17051 10186 17057
rect 10128 17048 10140 17051
rect 9548 17020 10140 17048
rect 9548 17008 9554 17020
rect 10128 17017 10140 17020
rect 10174 17048 10186 17051
rect 11698 17048 11704 17060
rect 10174 17020 11704 17048
rect 10174 17017 10186 17020
rect 10128 17011 10186 17017
rect 11698 17008 11704 17020
rect 11756 17008 11762 17060
rect 12526 17008 12532 17060
rect 12584 17048 12590 17060
rect 12682 17051 12740 17057
rect 12682 17048 12694 17051
rect 12584 17020 12694 17048
rect 12584 17008 12590 17020
rect 12682 17017 12694 17020
rect 12728 17017 12740 17051
rect 12682 17011 12740 17017
rect 16301 17051 16359 17057
rect 16301 17017 16313 17051
rect 16347 17048 16359 17051
rect 16574 17048 16580 17060
rect 16347 17020 16580 17048
rect 16347 17017 16359 17020
rect 16301 17011 16359 17017
rect 16574 17008 16580 17020
rect 16632 17048 16638 17060
rect 16960 17048 16988 17147
rect 18414 17144 18420 17196
rect 18472 17144 18478 17196
rect 18598 17184 18604 17196
rect 18559 17156 18604 17184
rect 18598 17144 18604 17156
rect 18656 17144 18662 17196
rect 21376 17184 21404 17280
rect 22756 17252 22784 17280
rect 21744 17224 22784 17252
rect 21634 17184 21640 17196
rect 21376 17156 21640 17184
rect 21634 17144 21640 17156
rect 21692 17144 21698 17196
rect 18432 17116 18460 17144
rect 18509 17119 18567 17125
rect 18509 17116 18521 17119
rect 18432 17088 18521 17116
rect 18509 17085 18521 17088
rect 18555 17085 18567 17119
rect 18509 17079 18567 17085
rect 19521 17119 19579 17125
rect 19521 17085 19533 17119
rect 19567 17116 19579 17119
rect 19613 17119 19671 17125
rect 19613 17116 19625 17119
rect 19567 17088 19625 17116
rect 19567 17085 19579 17088
rect 19521 17079 19579 17085
rect 19613 17085 19625 17088
rect 19659 17116 19671 17119
rect 21744 17116 21772 17224
rect 23492 17184 23520 17280
rect 24213 17187 24271 17193
rect 24213 17184 24225 17187
rect 23492 17156 24225 17184
rect 24213 17153 24225 17156
rect 24259 17153 24271 17187
rect 24213 17147 24271 17153
rect 22462 17116 22468 17128
rect 19659 17088 21772 17116
rect 22423 17088 22468 17116
rect 19659 17085 19671 17088
rect 19613 17079 19671 17085
rect 22462 17076 22468 17088
rect 22520 17076 22526 17128
rect 23658 17076 23664 17128
rect 23716 17116 23722 17128
rect 24029 17119 24087 17125
rect 24029 17116 24041 17119
rect 23716 17088 24041 17116
rect 23716 17076 23722 17088
rect 24029 17085 24041 17088
rect 24075 17116 24087 17119
rect 24670 17116 24676 17128
rect 24075 17088 24676 17116
rect 24075 17085 24087 17088
rect 24029 17079 24087 17085
rect 24670 17076 24676 17088
rect 24728 17076 24734 17128
rect 25225 17119 25283 17125
rect 25225 17085 25237 17119
rect 25271 17116 25283 17119
rect 25884 17116 25912 17283
rect 26142 17280 26148 17292
rect 26200 17280 26206 17332
rect 25271 17088 25912 17116
rect 25271 17085 25283 17088
rect 25225 17079 25283 17085
rect 16632 17020 16988 17048
rect 18417 17051 18475 17057
rect 16632 17008 16638 17020
rect 18417 17017 18429 17051
rect 18463 17048 18475 17051
rect 19150 17048 19156 17060
rect 18463 17020 19156 17048
rect 18463 17017 18475 17020
rect 18417 17011 18475 17017
rect 19150 17008 19156 17020
rect 19208 17008 19214 17060
rect 19702 17008 19708 17060
rect 19760 17048 19766 17060
rect 19858 17051 19916 17057
rect 19858 17048 19870 17051
rect 19760 17020 19870 17048
rect 19760 17008 19766 17020
rect 19858 17017 19870 17020
rect 19904 17048 19916 17051
rect 20622 17048 20628 17060
rect 19904 17020 20628 17048
rect 19904 17017 19916 17020
rect 19858 17011 19916 17017
rect 20622 17008 20628 17020
rect 20680 17008 20686 17060
rect 21726 17008 21732 17060
rect 21784 17048 21790 17060
rect 22554 17048 22560 17060
rect 21784 17020 22560 17048
rect 21784 17008 21790 17020
rect 22554 17008 22560 17020
rect 22612 17008 22618 17060
rect 23750 17008 23756 17060
rect 23808 17048 23814 17060
rect 24121 17051 24179 17057
rect 24121 17048 24133 17051
rect 23808 17020 24133 17048
rect 23808 17008 23814 17020
rect 24121 17017 24133 17020
rect 24167 17048 24179 17051
rect 24765 17051 24823 17057
rect 24765 17048 24777 17051
rect 24167 17020 24777 17048
rect 24167 17017 24179 17020
rect 24121 17011 24179 17017
rect 24765 17017 24777 17020
rect 24811 17017 24823 17051
rect 24765 17011 24823 17017
rect 25314 17008 25320 17060
rect 25372 17048 25378 17060
rect 26142 17048 26148 17060
rect 25372 17020 26148 17048
rect 25372 17008 25378 17020
rect 26142 17008 26148 17020
rect 26200 17008 26206 17060
rect 1302 16940 1308 16992
rect 1360 16980 1366 16992
rect 2038 16980 2044 16992
rect 1360 16952 2044 16980
rect 1360 16940 1366 16952
rect 2038 16940 2044 16952
rect 2096 16940 2102 16992
rect 3418 16980 3424 16992
rect 3331 16952 3424 16980
rect 3418 16940 3424 16952
rect 3476 16980 3482 16992
rect 4154 16980 4160 16992
rect 3476 16952 4160 16980
rect 3476 16940 3482 16952
rect 4154 16940 4160 16952
rect 4212 16940 4218 16992
rect 4982 16980 4988 16992
rect 4943 16952 4988 16980
rect 4982 16940 4988 16952
rect 5040 16980 5046 16992
rect 5629 16983 5687 16989
rect 5629 16980 5641 16983
rect 5040 16952 5641 16980
rect 5040 16940 5046 16952
rect 5629 16949 5641 16952
rect 5675 16949 5687 16983
rect 7006 16980 7012 16992
rect 6967 16952 7012 16980
rect 5629 16943 5687 16949
rect 7006 16940 7012 16952
rect 7064 16940 7070 16992
rect 8294 16980 8300 16992
rect 8255 16952 8300 16980
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 13446 16940 13452 16992
rect 13504 16980 13510 16992
rect 13817 16983 13875 16989
rect 13817 16980 13829 16983
rect 13504 16952 13829 16980
rect 13504 16940 13510 16952
rect 13817 16949 13829 16952
rect 13863 16949 13875 16983
rect 14918 16980 14924 16992
rect 14879 16952 14924 16980
rect 13817 16943 13875 16949
rect 14918 16940 14924 16952
rect 14976 16940 14982 16992
rect 16390 16980 16396 16992
rect 16351 16952 16396 16980
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 16850 16980 16856 16992
rect 16811 16952 16856 16980
rect 16850 16940 16856 16952
rect 16908 16940 16914 16992
rect 18046 16980 18052 16992
rect 18007 16952 18052 16980
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 20714 16940 20720 16992
rect 20772 16980 20778 16992
rect 20993 16983 21051 16989
rect 20993 16980 21005 16983
rect 20772 16952 21005 16980
rect 20772 16940 20778 16952
rect 20993 16949 21005 16952
rect 21039 16980 21051 16983
rect 21266 16980 21272 16992
rect 21039 16952 21272 16980
rect 21039 16949 21051 16952
rect 20993 16943 21051 16949
rect 21266 16940 21272 16952
rect 21324 16940 21330 16992
rect 22646 16980 22652 16992
rect 22607 16952 22652 16980
rect 22646 16940 22652 16952
rect 22704 16940 22710 16992
rect 23106 16940 23112 16992
rect 23164 16980 23170 16992
rect 24946 16980 24952 16992
rect 23164 16952 24952 16980
rect 23164 16940 23170 16952
rect 24946 16940 24952 16952
rect 25004 16980 25010 16992
rect 25041 16983 25099 16989
rect 25041 16980 25053 16983
rect 25004 16952 25053 16980
rect 25004 16940 25010 16952
rect 25041 16949 25053 16952
rect 25087 16949 25099 16983
rect 25041 16943 25099 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 3234 16776 3240 16788
rect 2832 16748 2877 16776
rect 3195 16748 3240 16776
rect 2832 16736 2838 16748
rect 3234 16736 3240 16748
rect 3292 16736 3298 16788
rect 3786 16776 3792 16788
rect 3747 16748 3792 16776
rect 3786 16736 3792 16748
rect 3844 16736 3850 16788
rect 4154 16736 4160 16788
rect 4212 16736 4218 16788
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 6365 16779 6423 16785
rect 6365 16776 6377 16779
rect 5592 16748 6377 16776
rect 5592 16736 5598 16748
rect 6365 16745 6377 16748
rect 6411 16745 6423 16779
rect 6365 16739 6423 16745
rect 8294 16736 8300 16788
rect 8352 16776 8358 16788
rect 8849 16779 8907 16785
rect 8849 16776 8861 16779
rect 8352 16748 8861 16776
rect 8352 16736 8358 16748
rect 8849 16745 8861 16748
rect 8895 16745 8907 16779
rect 9490 16776 9496 16788
rect 9451 16748 9496 16776
rect 8849 16739 8907 16745
rect 9490 16736 9496 16748
rect 9548 16736 9554 16788
rect 9950 16776 9956 16788
rect 9911 16748 9956 16776
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 12618 16736 12624 16788
rect 12676 16776 12682 16788
rect 12802 16776 12808 16788
rect 12676 16748 12808 16776
rect 12676 16736 12682 16748
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 14550 16776 14556 16788
rect 14511 16748 14556 16776
rect 14550 16736 14556 16748
rect 14608 16736 14614 16788
rect 15565 16779 15623 16785
rect 15565 16745 15577 16779
rect 15611 16776 15623 16779
rect 16117 16779 16175 16785
rect 16117 16776 16129 16779
rect 15611 16748 16129 16776
rect 15611 16745 15623 16748
rect 15565 16739 15623 16745
rect 16117 16745 16129 16748
rect 16163 16776 16175 16779
rect 16390 16776 16396 16788
rect 16163 16748 16396 16776
rect 16163 16745 16175 16748
rect 16117 16739 16175 16745
rect 16390 16736 16396 16748
rect 16448 16736 16454 16788
rect 18325 16779 18383 16785
rect 18325 16745 18337 16779
rect 18371 16776 18383 16779
rect 18414 16776 18420 16788
rect 18371 16748 18420 16776
rect 18371 16745 18383 16748
rect 18325 16739 18383 16745
rect 18414 16736 18420 16748
rect 18472 16736 18478 16788
rect 19242 16776 19248 16788
rect 19203 16748 19248 16776
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 19426 16736 19432 16788
rect 19484 16776 19490 16788
rect 19705 16779 19763 16785
rect 19705 16776 19717 16779
rect 19484 16748 19717 16776
rect 19484 16736 19490 16748
rect 19705 16745 19717 16748
rect 19751 16745 19763 16779
rect 20254 16776 20260 16788
rect 20215 16748 20260 16776
rect 19705 16739 19763 16745
rect 20254 16736 20260 16748
rect 20312 16736 20318 16788
rect 20622 16776 20628 16788
rect 20583 16748 20628 16776
rect 20622 16736 20628 16748
rect 20680 16736 20686 16788
rect 20901 16779 20959 16785
rect 20901 16745 20913 16779
rect 20947 16745 20959 16779
rect 21266 16776 21272 16788
rect 21227 16748 21272 16776
rect 20901 16739 20959 16745
rect 2130 16708 2136 16720
rect 2043 16680 2136 16708
rect 2130 16668 2136 16680
rect 2188 16708 2194 16720
rect 4172 16708 4200 16736
rect 4310 16711 4368 16717
rect 4310 16708 4322 16711
rect 2188 16680 4108 16708
rect 4172 16680 4322 16708
rect 2188 16668 2194 16680
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 1670 16640 1676 16652
rect 1443 16612 1676 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 1670 16600 1676 16612
rect 1728 16600 1734 16652
rect 2869 16643 2927 16649
rect 2869 16609 2881 16643
rect 2915 16640 2927 16643
rect 3786 16640 3792 16652
rect 2915 16612 3792 16640
rect 2915 16609 2927 16612
rect 2869 16603 2927 16609
rect 3786 16600 3792 16612
rect 3844 16600 3850 16652
rect 4080 16649 4108 16680
rect 4310 16677 4322 16680
rect 4356 16677 4368 16711
rect 6086 16708 6092 16720
rect 6047 16680 6092 16708
rect 4310 16671 4368 16677
rect 6086 16668 6092 16680
rect 6144 16668 6150 16720
rect 6730 16668 6736 16720
rect 6788 16717 6794 16720
rect 6788 16711 6852 16717
rect 6788 16677 6806 16711
rect 6840 16677 6852 16711
rect 6788 16671 6852 16677
rect 8573 16711 8631 16717
rect 8573 16677 8585 16711
rect 8619 16708 8631 16711
rect 9508 16708 9536 16736
rect 8619 16680 9536 16708
rect 8619 16677 8631 16680
rect 8573 16671 8631 16677
rect 6788 16668 6794 16671
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16640 4123 16643
rect 4798 16640 4804 16652
rect 4111 16612 4804 16640
rect 4111 16609 4123 16612
rect 4065 16603 4123 16609
rect 4798 16600 4804 16612
rect 4856 16600 4862 16652
rect 9968 16640 9996 16736
rect 10588 16711 10646 16717
rect 10588 16677 10600 16711
rect 10634 16708 10646 16711
rect 11146 16708 11152 16720
rect 10634 16680 11152 16708
rect 10634 16677 10646 16680
rect 10588 16671 10646 16677
rect 11146 16668 11152 16680
rect 11204 16668 11210 16720
rect 12894 16668 12900 16720
rect 12952 16708 12958 16720
rect 13909 16711 13967 16717
rect 13909 16708 13921 16711
rect 12952 16680 13921 16708
rect 12952 16668 12958 16680
rect 13909 16677 13921 16680
rect 13955 16708 13967 16711
rect 14826 16708 14832 16720
rect 13955 16680 14832 16708
rect 13955 16677 13967 16680
rect 13909 16671 13967 16677
rect 14826 16668 14832 16680
rect 14884 16668 14890 16720
rect 17494 16668 17500 16720
rect 17552 16708 17558 16720
rect 18598 16708 18604 16720
rect 17552 16680 18604 16708
rect 17552 16668 17558 16680
rect 10318 16640 10324 16652
rect 9968 16612 10324 16640
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 12526 16640 12532 16652
rect 12487 16612 12532 16640
rect 12526 16600 12532 16612
rect 12584 16600 12590 16652
rect 13170 16640 13176 16652
rect 13131 16612 13176 16640
rect 13170 16600 13176 16612
rect 13228 16600 13234 16652
rect 13722 16600 13728 16652
rect 13780 16640 13786 16652
rect 14185 16643 14243 16649
rect 14185 16640 14197 16643
rect 13780 16612 14197 16640
rect 13780 16600 13786 16612
rect 14185 16609 14197 16612
rect 14231 16609 14243 16643
rect 15102 16640 15108 16652
rect 15063 16612 15108 16640
rect 14185 16603 14243 16609
rect 15102 16600 15108 16612
rect 15160 16600 15166 16652
rect 16022 16640 16028 16652
rect 15983 16612 16028 16640
rect 16022 16600 16028 16612
rect 16080 16600 16086 16652
rect 16850 16640 16856 16652
rect 16592 16612 16856 16640
rect 2774 16532 2780 16584
rect 2832 16572 2838 16584
rect 2961 16575 3019 16581
rect 2961 16572 2973 16575
rect 2832 16544 2973 16572
rect 2832 16532 2838 16544
rect 2961 16541 2973 16544
rect 3007 16572 3019 16575
rect 6546 16572 6552 16584
rect 3007 16544 4108 16572
rect 6507 16544 6552 16572
rect 3007 16541 3019 16544
rect 2961 16535 3019 16541
rect 1581 16507 1639 16513
rect 1581 16473 1593 16507
rect 1627 16504 1639 16507
rect 3510 16504 3516 16516
rect 1627 16476 3516 16504
rect 1627 16473 1639 16476
rect 1581 16467 1639 16473
rect 3510 16464 3516 16476
rect 3568 16464 3574 16516
rect 2406 16436 2412 16448
rect 2367 16408 2412 16436
rect 2406 16396 2412 16408
rect 2464 16396 2470 16448
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 3237 16439 3295 16445
rect 3237 16436 3249 16439
rect 2832 16408 3249 16436
rect 2832 16396 2838 16408
rect 3237 16405 3249 16408
rect 3283 16436 3295 16439
rect 3421 16439 3479 16445
rect 3421 16436 3433 16439
rect 3283 16408 3433 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 3421 16405 3433 16408
rect 3467 16405 3479 16439
rect 4080 16436 4108 16544
rect 6546 16532 6552 16544
rect 6604 16532 6610 16584
rect 13262 16572 13268 16584
rect 13223 16544 13268 16572
rect 13262 16532 13268 16544
rect 13320 16532 13326 16584
rect 13446 16572 13452 16584
rect 13407 16544 13452 16572
rect 13446 16532 13452 16544
rect 13504 16532 13510 16584
rect 13906 16532 13912 16584
rect 13964 16572 13970 16584
rect 14642 16572 14648 16584
rect 13964 16544 14648 16572
rect 13964 16532 13970 16544
rect 14642 16532 14648 16544
rect 14700 16532 14706 16584
rect 15562 16532 15568 16584
rect 15620 16572 15626 16584
rect 16209 16575 16267 16581
rect 16209 16572 16221 16575
rect 15620 16544 16221 16572
rect 15620 16532 15626 16544
rect 16209 16541 16221 16544
rect 16255 16541 16267 16575
rect 16209 16535 16267 16541
rect 16390 16532 16396 16584
rect 16448 16572 16454 16584
rect 16592 16572 16620 16612
rect 16850 16600 16856 16612
rect 16908 16640 16914 16652
rect 17037 16643 17095 16649
rect 17037 16640 17049 16643
rect 16908 16612 17049 16640
rect 16908 16600 16914 16612
rect 17037 16609 17049 16612
rect 17083 16609 17095 16643
rect 17037 16603 17095 16609
rect 17126 16600 17132 16652
rect 17184 16640 17190 16652
rect 17589 16643 17647 16649
rect 17589 16640 17601 16643
rect 17184 16612 17601 16640
rect 17184 16600 17190 16612
rect 17589 16609 17601 16612
rect 17635 16609 17647 16643
rect 17589 16603 17647 16609
rect 17678 16572 17684 16584
rect 16448 16544 16620 16572
rect 17591 16544 17684 16572
rect 16448 16532 16454 16544
rect 17678 16532 17684 16544
rect 17736 16532 17742 16584
rect 17788 16581 17816 16680
rect 18598 16668 18604 16680
rect 18656 16668 18662 16720
rect 20916 16708 20944 16739
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 21910 16776 21916 16788
rect 21871 16748 21916 16776
rect 21910 16736 21916 16748
rect 21968 16736 21974 16788
rect 22462 16776 22468 16788
rect 22423 16748 22468 16776
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 24121 16779 24179 16785
rect 24121 16745 24133 16779
rect 24167 16776 24179 16779
rect 24670 16776 24676 16788
rect 24167 16748 24676 16776
rect 24167 16745 24179 16748
rect 24121 16739 24179 16745
rect 24670 16736 24676 16748
rect 24728 16736 24734 16788
rect 25038 16776 25044 16788
rect 24999 16748 25044 16776
rect 25038 16736 25044 16748
rect 25096 16736 25102 16788
rect 25409 16779 25467 16785
rect 25409 16745 25421 16779
rect 25455 16776 25467 16779
rect 25682 16776 25688 16788
rect 25455 16748 25688 16776
rect 25455 16745 25467 16748
rect 25409 16739 25467 16745
rect 25682 16736 25688 16748
rect 25740 16736 25746 16788
rect 19628 16680 20944 16708
rect 19628 16652 19656 16680
rect 20990 16668 20996 16720
rect 21048 16708 21054 16720
rect 21361 16711 21419 16717
rect 21361 16708 21373 16711
rect 21048 16680 21373 16708
rect 21048 16668 21054 16680
rect 21361 16677 21373 16680
rect 21407 16677 21419 16711
rect 21361 16671 21419 16677
rect 23008 16711 23066 16717
rect 23008 16677 23020 16711
rect 23054 16708 23066 16711
rect 23290 16708 23296 16720
rect 23054 16680 23296 16708
rect 23054 16677 23066 16680
rect 23008 16671 23066 16677
rect 23290 16668 23296 16680
rect 23348 16708 23354 16720
rect 24210 16708 24216 16720
rect 23348 16680 24216 16708
rect 23348 16668 23354 16680
rect 24210 16668 24216 16680
rect 24268 16668 24274 16720
rect 18966 16600 18972 16652
rect 19024 16640 19030 16652
rect 19150 16640 19156 16652
rect 19024 16612 19156 16640
rect 19024 16600 19030 16612
rect 19150 16600 19156 16612
rect 19208 16600 19214 16652
rect 19610 16640 19616 16652
rect 19571 16612 19616 16640
rect 19610 16600 19616 16612
rect 19668 16600 19674 16652
rect 22738 16640 22744 16652
rect 22699 16612 22744 16640
rect 22738 16600 22744 16612
rect 22796 16600 22802 16652
rect 23750 16600 23756 16652
rect 23808 16640 23814 16652
rect 23934 16640 23940 16652
rect 23808 16612 23940 16640
rect 23808 16600 23814 16612
rect 23934 16600 23940 16612
rect 23992 16600 23998 16652
rect 25225 16643 25283 16649
rect 25225 16609 25237 16643
rect 25271 16640 25283 16643
rect 25314 16640 25320 16652
rect 25271 16612 25320 16640
rect 25271 16609 25283 16612
rect 25225 16603 25283 16609
rect 25314 16600 25320 16612
rect 25372 16600 25378 16652
rect 17773 16575 17831 16581
rect 17773 16541 17785 16575
rect 17819 16541 17831 16575
rect 17773 16535 17831 16541
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16572 19855 16575
rect 20714 16572 20720 16584
rect 19843 16544 20720 16572
rect 19843 16541 19855 16544
rect 19797 16535 19855 16541
rect 17696 16504 17724 16532
rect 17862 16504 17868 16516
rect 5276 16476 6040 16504
rect 17696 16476 17868 16504
rect 5276 16436 5304 16476
rect 5442 16436 5448 16448
rect 4080 16408 5304 16436
rect 5403 16408 5448 16436
rect 3421 16399 3479 16405
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 6012 16436 6040 16476
rect 17862 16464 17868 16476
rect 17920 16464 17926 16516
rect 19334 16464 19340 16516
rect 19392 16504 19398 16516
rect 19812 16504 19840 16535
rect 20714 16532 20720 16544
rect 20772 16532 20778 16584
rect 21545 16575 21603 16581
rect 21545 16541 21557 16575
rect 21591 16541 21603 16575
rect 21545 16535 21603 16541
rect 19392 16476 19840 16504
rect 19392 16464 19398 16476
rect 20622 16464 20628 16516
rect 20680 16504 20686 16516
rect 21450 16504 21456 16516
rect 20680 16476 21456 16504
rect 20680 16464 20686 16476
rect 21450 16464 21456 16476
rect 21508 16504 21514 16516
rect 21560 16504 21588 16535
rect 21508 16476 21588 16504
rect 21508 16464 21514 16476
rect 23934 16464 23940 16516
rect 23992 16504 23998 16516
rect 24673 16507 24731 16513
rect 24673 16504 24685 16507
rect 23992 16476 24685 16504
rect 23992 16464 23998 16476
rect 24673 16473 24685 16476
rect 24719 16473 24731 16507
rect 24673 16467 24731 16473
rect 7929 16439 7987 16445
rect 7929 16436 7941 16439
rect 6012 16408 7941 16436
rect 7929 16405 7941 16408
rect 7975 16436 7987 16439
rect 8110 16436 8116 16448
rect 7975 16408 8116 16436
rect 7975 16405 7987 16408
rect 7929 16399 7987 16405
rect 8110 16396 8116 16408
rect 8168 16396 8174 16448
rect 11698 16436 11704 16448
rect 11659 16408 11704 16436
rect 11698 16396 11704 16408
rect 11756 16396 11762 16448
rect 12802 16436 12808 16448
rect 12763 16408 12808 16436
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 15654 16436 15660 16448
rect 15615 16408 15660 16436
rect 15654 16396 15660 16408
rect 15712 16396 15718 16448
rect 16758 16436 16764 16448
rect 16719 16408 16764 16436
rect 16758 16396 16764 16408
rect 16816 16396 16822 16448
rect 17218 16436 17224 16448
rect 17179 16408 17224 16436
rect 17218 16396 17224 16408
rect 17276 16396 17282 16448
rect 22646 16396 22652 16448
rect 22704 16436 22710 16448
rect 25777 16439 25835 16445
rect 25777 16436 25789 16439
rect 22704 16408 25789 16436
rect 22704 16396 22710 16408
rect 25777 16405 25789 16408
rect 25823 16405 25835 16439
rect 25777 16399 25835 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2038 16232 2044 16244
rect 1999 16204 2044 16232
rect 2038 16192 2044 16204
rect 2096 16192 2102 16244
rect 2130 16192 2136 16244
rect 2188 16232 2194 16244
rect 3418 16232 3424 16244
rect 2188 16204 3424 16232
rect 2188 16192 2194 16204
rect 3418 16192 3424 16204
rect 3476 16192 3482 16244
rect 5077 16235 5135 16241
rect 5077 16201 5089 16235
rect 5123 16232 5135 16235
rect 5534 16232 5540 16244
rect 5123 16204 5540 16232
rect 5123 16201 5135 16204
rect 5077 16195 5135 16201
rect 5534 16192 5540 16204
rect 5592 16192 5598 16244
rect 6730 16192 6736 16244
rect 6788 16232 6794 16244
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 6788 16204 8217 16232
rect 6788 16192 6794 16204
rect 8205 16201 8217 16204
rect 8251 16201 8263 16235
rect 8205 16195 8263 16201
rect 9122 16192 9128 16244
rect 9180 16232 9186 16244
rect 9493 16235 9551 16241
rect 9493 16232 9505 16235
rect 9180 16204 9505 16232
rect 9180 16192 9186 16204
rect 9493 16201 9505 16204
rect 9539 16201 9551 16235
rect 9674 16232 9680 16244
rect 9635 16204 9680 16232
rect 9493 16195 9551 16201
rect 3605 16167 3663 16173
rect 3605 16133 3617 16167
rect 3651 16164 3663 16167
rect 3786 16164 3792 16176
rect 3651 16136 3792 16164
rect 3651 16133 3663 16136
rect 3605 16127 3663 16133
rect 3786 16124 3792 16136
rect 3844 16124 3850 16176
rect 2498 16096 2504 16108
rect 2459 16068 2504 16096
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16096 2743 16099
rect 2774 16096 2780 16108
rect 2731 16068 2780 16096
rect 2731 16065 2743 16068
rect 2685 16059 2743 16065
rect 2774 16056 2780 16068
rect 2832 16056 2838 16108
rect 3878 16056 3884 16108
rect 3936 16096 3942 16108
rect 4157 16099 4215 16105
rect 4157 16096 4169 16099
rect 3936 16068 4169 16096
rect 3936 16056 3942 16068
rect 4157 16065 4169 16068
rect 4203 16065 4215 16099
rect 5552 16096 5580 16192
rect 5721 16099 5779 16105
rect 5721 16096 5733 16099
rect 5552 16068 5733 16096
rect 4157 16059 4215 16065
rect 5721 16065 5733 16068
rect 5767 16096 5779 16099
rect 6086 16096 6092 16108
rect 5767 16068 6092 16096
rect 5767 16065 5779 16068
rect 5721 16059 5779 16065
rect 6086 16056 6092 16068
rect 6144 16096 6150 16108
rect 9508 16096 9536 16195
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 10689 16235 10747 16241
rect 10689 16232 10701 16235
rect 10376 16204 10701 16232
rect 10376 16192 10382 16204
rect 10689 16201 10701 16204
rect 10735 16232 10747 16235
rect 10870 16232 10876 16244
rect 10735 16204 10876 16232
rect 10735 16201 10747 16204
rect 10689 16195 10747 16201
rect 10870 16192 10876 16204
rect 10928 16192 10934 16244
rect 11146 16232 11152 16244
rect 11107 16204 11152 16232
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 11882 16232 11888 16244
rect 11843 16204 11888 16232
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 12342 16192 12348 16244
rect 12400 16232 12406 16244
rect 12437 16235 12495 16241
rect 12437 16232 12449 16235
rect 12400 16204 12449 16232
rect 12400 16192 12406 16204
rect 12437 16201 12449 16204
rect 12483 16201 12495 16235
rect 13446 16232 13452 16244
rect 13407 16204 13452 16232
rect 12437 16195 12495 16201
rect 13446 16192 13452 16204
rect 13504 16192 13510 16244
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 14001 16235 14059 16241
rect 14001 16232 14013 16235
rect 13872 16204 14013 16232
rect 13872 16192 13878 16204
rect 14001 16201 14013 16204
rect 14047 16201 14059 16235
rect 14001 16195 14059 16201
rect 14274 16192 14280 16244
rect 14332 16232 14338 16244
rect 14550 16232 14556 16244
rect 14332 16204 14556 16232
rect 14332 16192 14338 16204
rect 14550 16192 14556 16204
rect 14608 16192 14614 16244
rect 16390 16232 16396 16244
rect 16351 16204 16396 16232
rect 16390 16192 16396 16204
rect 16448 16192 16454 16244
rect 18601 16235 18659 16241
rect 18601 16201 18613 16235
rect 18647 16232 18659 16235
rect 19058 16232 19064 16244
rect 18647 16204 19064 16232
rect 18647 16201 18659 16204
rect 18601 16195 18659 16201
rect 19058 16192 19064 16204
rect 19116 16192 19122 16244
rect 20441 16235 20499 16241
rect 20441 16201 20453 16235
rect 20487 16232 20499 16235
rect 20622 16232 20628 16244
rect 20487 16204 20628 16232
rect 20487 16201 20499 16204
rect 20441 16195 20499 16201
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 20898 16192 20904 16244
rect 20956 16232 20962 16244
rect 21085 16235 21143 16241
rect 21085 16232 21097 16235
rect 20956 16204 21097 16232
rect 20956 16192 20962 16204
rect 21085 16201 21097 16204
rect 21131 16201 21143 16235
rect 21085 16195 21143 16201
rect 11164 16164 11192 16192
rect 16298 16164 16304 16176
rect 10336 16136 11192 16164
rect 16259 16136 16304 16164
rect 10336 16105 10364 16136
rect 16298 16124 16304 16136
rect 16356 16124 16362 16176
rect 17862 16164 17868 16176
rect 17823 16136 17868 16164
rect 17862 16124 17868 16136
rect 17920 16124 17926 16176
rect 18506 16124 18512 16176
rect 18564 16164 18570 16176
rect 18690 16164 18696 16176
rect 18564 16136 18696 16164
rect 18564 16124 18570 16136
rect 18690 16124 18696 16136
rect 18748 16164 18754 16176
rect 18877 16167 18935 16173
rect 18877 16164 18889 16167
rect 18748 16136 18889 16164
rect 18748 16124 18754 16136
rect 18877 16133 18889 16136
rect 18923 16164 18935 16167
rect 18923 16136 19104 16164
rect 18923 16133 18935 16136
rect 18877 16127 18935 16133
rect 10137 16099 10195 16105
rect 10137 16096 10149 16099
rect 6144 16068 6960 16096
rect 9508 16068 10149 16096
rect 6144 16056 6150 16068
rect 3694 15988 3700 16040
rect 3752 16028 3758 16040
rect 3973 16031 4031 16037
rect 3973 16028 3985 16031
rect 3752 16000 3985 16028
rect 3752 15988 3758 16000
rect 3973 15997 3985 16000
rect 4019 15997 4031 16031
rect 3973 15991 4031 15997
rect 6546 15988 6552 16040
rect 6604 16028 6610 16040
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6604 16000 6837 16028
rect 6604 15988 6610 16000
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 6932 16028 6960 16068
rect 10137 16065 10149 16068
rect 10183 16065 10195 16099
rect 10137 16059 10195 16065
rect 10321 16099 10379 16105
rect 10321 16065 10333 16099
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 7081 16031 7139 16037
rect 7081 16028 7093 16031
rect 6932 16000 7093 16028
rect 6825 15991 6883 15997
rect 7081 15997 7093 16000
rect 7127 15997 7139 16031
rect 7081 15991 7139 15997
rect 8849 16031 8907 16037
rect 8849 15997 8861 16031
rect 8895 16028 8907 16031
rect 10336 16028 10364 16059
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 12253 16099 12311 16105
rect 12253 16096 12265 16099
rect 11756 16068 12265 16096
rect 11756 16056 11762 16068
rect 12253 16065 12265 16068
rect 12299 16096 12311 16099
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 12299 16068 13001 16096
rect 12299 16065 12311 16068
rect 12253 16059 12311 16065
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 13170 16056 13176 16108
rect 13228 16096 13234 16108
rect 13446 16096 13452 16108
rect 13228 16068 13452 16096
rect 13228 16056 13234 16068
rect 13446 16056 13452 16068
rect 13504 16056 13510 16108
rect 13814 16056 13820 16108
rect 13872 16096 13878 16108
rect 14553 16099 14611 16105
rect 14553 16096 14565 16099
rect 13872 16068 14565 16096
rect 13872 16056 13878 16068
rect 14553 16065 14565 16068
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 16758 16056 16764 16108
rect 16816 16096 16822 16108
rect 16945 16099 17003 16105
rect 16945 16096 16957 16099
rect 16816 16068 16957 16096
rect 16816 16056 16822 16068
rect 16945 16065 16957 16068
rect 16991 16096 17003 16099
rect 17494 16096 17500 16108
rect 16991 16068 17500 16096
rect 16991 16065 17003 16068
rect 16945 16059 17003 16065
rect 17494 16056 17500 16068
rect 17552 16056 17558 16108
rect 19076 16105 19104 16136
rect 19061 16099 19119 16105
rect 19061 16065 19073 16099
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 11238 16028 11244 16040
rect 8895 16000 10364 16028
rect 11199 16000 11244 16028
rect 8895 15997 8907 16000
rect 8849 15991 8907 15997
rect 11238 15988 11244 16000
rect 11296 15988 11302 16040
rect 12802 16028 12808 16040
rect 12715 16000 12808 16028
rect 12802 15988 12808 16000
rect 12860 16028 12866 16040
rect 15013 16031 15071 16037
rect 15013 16028 15025 16031
rect 12860 16000 15025 16028
rect 12860 15988 12866 16000
rect 15013 15997 15025 16000
rect 15059 15997 15071 16031
rect 15013 15991 15071 15997
rect 15933 16031 15991 16037
rect 15933 15997 15945 16031
rect 15979 16028 15991 16031
rect 16853 16031 16911 16037
rect 16853 16028 16865 16031
rect 15979 16000 16865 16028
rect 15979 15997 15991 16000
rect 15933 15991 15991 15997
rect 16853 15997 16865 16000
rect 16899 16028 16911 16031
rect 17034 16028 17040 16040
rect 16899 16000 17040 16028
rect 16899 15997 16911 16000
rect 16853 15991 16911 15997
rect 17034 15988 17040 16000
rect 17092 16028 17098 16040
rect 17678 16028 17684 16040
rect 17092 16000 17684 16028
rect 17092 15988 17098 16000
rect 17678 15988 17684 16000
rect 17736 15988 17742 16040
rect 2682 15920 2688 15972
rect 2740 15960 2746 15972
rect 3053 15963 3111 15969
rect 3053 15960 3065 15963
rect 2740 15932 3065 15960
rect 2740 15920 2746 15932
rect 3053 15929 3065 15932
rect 3099 15929 3111 15963
rect 3053 15923 3111 15929
rect 4065 15963 4123 15969
rect 4065 15929 4077 15963
rect 4111 15960 4123 15963
rect 5537 15963 5595 15969
rect 4111 15932 5212 15960
rect 4111 15929 4123 15932
rect 4065 15923 4123 15929
rect 5184 15904 5212 15932
rect 5537 15929 5549 15963
rect 5583 15960 5595 15963
rect 9217 15963 9275 15969
rect 5583 15932 6868 15960
rect 5583 15929 5595 15932
rect 5537 15923 5595 15929
rect 6840 15904 6868 15932
rect 9217 15929 9229 15963
rect 9263 15960 9275 15963
rect 10045 15963 10103 15969
rect 10045 15960 10057 15963
rect 9263 15932 10057 15960
rect 9263 15929 9275 15932
rect 9217 15923 9275 15929
rect 10045 15929 10057 15932
rect 10091 15960 10103 15963
rect 10962 15960 10968 15972
rect 10091 15932 10968 15960
rect 10091 15929 10103 15932
rect 10045 15923 10103 15929
rect 10962 15920 10968 15932
rect 11020 15920 11026 15972
rect 12434 15920 12440 15972
rect 12492 15960 12498 15972
rect 12897 15963 12955 15969
rect 12897 15960 12909 15963
rect 12492 15932 12909 15960
rect 12492 15920 12498 15932
rect 12897 15929 12909 15932
rect 12943 15960 12955 15963
rect 13722 15960 13728 15972
rect 12943 15932 13728 15960
rect 12943 15929 12955 15932
rect 12897 15923 12955 15929
rect 13722 15920 13728 15932
rect 13780 15920 13786 15972
rect 13906 15920 13912 15972
rect 13964 15960 13970 15972
rect 14461 15963 14519 15969
rect 14461 15960 14473 15963
rect 13964 15932 14473 15960
rect 13964 15920 13970 15932
rect 14461 15929 14473 15932
rect 14507 15960 14519 15963
rect 14918 15960 14924 15972
rect 14507 15932 14924 15960
rect 14507 15929 14519 15932
rect 14461 15923 14519 15929
rect 14918 15920 14924 15932
rect 14976 15920 14982 15972
rect 16298 15920 16304 15972
rect 16356 15960 16362 15972
rect 16666 15960 16672 15972
rect 16356 15932 16672 15960
rect 16356 15920 16362 15932
rect 16666 15920 16672 15932
rect 16724 15960 16730 15972
rect 16761 15963 16819 15969
rect 16761 15960 16773 15963
rect 16724 15932 16773 15960
rect 16724 15920 16730 15932
rect 16761 15929 16773 15932
rect 16807 15929 16819 15963
rect 16761 15923 16819 15929
rect 19150 15920 19156 15972
rect 19208 15960 19214 15972
rect 19306 15963 19364 15969
rect 19306 15960 19318 15963
rect 19208 15932 19318 15960
rect 19208 15920 19214 15932
rect 19306 15929 19318 15932
rect 19352 15929 19364 15963
rect 19306 15923 19364 15929
rect 19426 15920 19432 15972
rect 19484 15960 19490 15972
rect 20070 15960 20076 15972
rect 19484 15932 20076 15960
rect 19484 15920 19490 15932
rect 20070 15920 20076 15932
rect 20128 15920 20134 15972
rect 21100 15960 21128 16195
rect 22462 16192 22468 16244
rect 22520 16232 22526 16244
rect 22738 16232 22744 16244
rect 22520 16204 22744 16232
rect 22520 16192 22526 16204
rect 22738 16192 22744 16204
rect 22796 16192 22802 16244
rect 23201 16235 23259 16241
rect 23201 16201 23213 16235
rect 23247 16232 23259 16235
rect 23290 16232 23296 16244
rect 23247 16204 23296 16232
rect 23247 16201 23259 16204
rect 23201 16195 23259 16201
rect 22094 16056 22100 16108
rect 22152 16096 22158 16108
rect 22281 16099 22339 16105
rect 22281 16096 22293 16099
rect 22152 16068 22293 16096
rect 22152 16056 22158 16068
rect 22281 16065 22293 16068
rect 22327 16096 22339 16099
rect 23216 16096 23244 16195
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 23658 16232 23664 16244
rect 23619 16204 23664 16232
rect 23658 16192 23664 16204
rect 23716 16192 23722 16244
rect 24854 16192 24860 16244
rect 24912 16232 24918 16244
rect 25409 16235 25467 16241
rect 25409 16232 25421 16235
rect 24912 16204 25421 16232
rect 24912 16192 24918 16204
rect 25409 16201 25421 16204
rect 25455 16201 25467 16235
rect 25409 16195 25467 16201
rect 25498 16192 25504 16244
rect 25556 16232 25562 16244
rect 25774 16232 25780 16244
rect 25556 16204 25780 16232
rect 25556 16192 25562 16204
rect 25774 16192 25780 16204
rect 25832 16192 25838 16244
rect 22327 16068 23244 16096
rect 22327 16065 22339 16068
rect 22281 16059 22339 16065
rect 24026 16056 24032 16108
rect 24084 16096 24090 16108
rect 24305 16099 24363 16105
rect 24305 16096 24317 16099
rect 24084 16068 24317 16096
rect 24084 16056 24090 16068
rect 24305 16065 24317 16068
rect 24351 16096 24363 16099
rect 24673 16099 24731 16105
rect 24673 16096 24685 16099
rect 24351 16068 24685 16096
rect 24351 16065 24363 16068
rect 24305 16059 24363 16065
rect 24673 16065 24685 16068
rect 24719 16065 24731 16099
rect 24673 16059 24731 16065
rect 21545 16031 21603 16037
rect 21545 15997 21557 16031
rect 21591 16028 21603 16031
rect 22002 16028 22008 16040
rect 21591 16000 22008 16028
rect 21591 15997 21603 16000
rect 21545 15991 21603 15997
rect 22002 15988 22008 16000
rect 22060 15988 22066 16040
rect 24854 15988 24860 16040
rect 24912 16028 24918 16040
rect 25225 16031 25283 16037
rect 25225 16028 25237 16031
rect 24912 16000 25237 16028
rect 24912 15988 24918 16000
rect 25225 15997 25237 16000
rect 25271 16028 25283 16031
rect 25777 16031 25835 16037
rect 25777 16028 25789 16031
rect 25271 16000 25789 16028
rect 25271 15997 25283 16000
rect 25225 15991 25283 15997
rect 25777 15997 25789 16000
rect 25823 15997 25835 16031
rect 26234 16028 26240 16040
rect 26195 16000 26240 16028
rect 25777 15991 25835 15997
rect 26234 15988 26240 16000
rect 26292 15988 26298 16040
rect 22097 15963 22155 15969
rect 22097 15960 22109 15963
rect 21100 15932 22109 15960
rect 22097 15929 22109 15932
rect 22143 15929 22155 15963
rect 22097 15923 22155 15929
rect 23934 15920 23940 15972
rect 23992 15960 23998 15972
rect 24121 15963 24179 15969
rect 24121 15960 24133 15963
rect 23992 15932 24133 15960
rect 23992 15920 23998 15932
rect 24121 15929 24133 15932
rect 24167 15929 24179 15963
rect 24121 15923 24179 15929
rect 25133 15963 25191 15969
rect 25133 15929 25145 15963
rect 25179 15960 25191 15963
rect 25314 15960 25320 15972
rect 25179 15932 25320 15960
rect 25179 15929 25191 15932
rect 25133 15923 25191 15929
rect 25314 15920 25320 15932
rect 25372 15960 25378 15972
rect 25866 15960 25872 15972
rect 25372 15932 25872 15960
rect 25372 15920 25378 15932
rect 25866 15920 25872 15932
rect 25924 15920 25930 15972
rect 1762 15852 1768 15904
rect 1820 15892 1826 15904
rect 1949 15895 2007 15901
rect 1949 15892 1961 15895
rect 1820 15864 1961 15892
rect 1820 15852 1826 15864
rect 1949 15861 1961 15864
rect 1995 15892 2007 15895
rect 2409 15895 2467 15901
rect 2409 15892 2421 15895
rect 1995 15864 2421 15892
rect 1995 15861 2007 15864
rect 1949 15855 2007 15861
rect 2409 15861 2421 15864
rect 2455 15892 2467 15895
rect 3326 15892 3332 15904
rect 2455 15864 3332 15892
rect 2455 15861 2467 15864
rect 2409 15855 2467 15861
rect 3326 15852 3332 15864
rect 3384 15852 3390 15904
rect 4709 15895 4767 15901
rect 4709 15861 4721 15895
rect 4755 15892 4767 15895
rect 4798 15892 4804 15904
rect 4755 15864 4804 15892
rect 4755 15861 4767 15864
rect 4709 15855 4767 15861
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 5166 15892 5172 15904
rect 5127 15864 5172 15892
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5626 15852 5632 15904
rect 5684 15892 5690 15904
rect 6273 15895 6331 15901
rect 5684 15864 5729 15892
rect 5684 15852 5690 15864
rect 6273 15861 6285 15895
rect 6319 15892 6331 15895
rect 6546 15892 6552 15904
rect 6319 15864 6552 15892
rect 6319 15861 6331 15864
rect 6273 15855 6331 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 6822 15852 6828 15904
rect 6880 15852 6886 15904
rect 13814 15892 13820 15904
rect 13775 15864 13820 15892
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 14366 15892 14372 15904
rect 14327 15864 14372 15892
rect 14366 15852 14372 15864
rect 14424 15852 14430 15904
rect 15562 15892 15568 15904
rect 15523 15864 15568 15892
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 17126 15852 17132 15904
rect 17184 15892 17190 15904
rect 17405 15895 17463 15901
rect 17405 15892 17417 15895
rect 17184 15864 17417 15892
rect 17184 15852 17190 15864
rect 17405 15861 17417 15864
rect 17451 15861 17463 15895
rect 17405 15855 17463 15861
rect 18049 15895 18107 15901
rect 18049 15861 18061 15895
rect 18095 15892 18107 15895
rect 18138 15892 18144 15904
rect 18095 15864 18144 15892
rect 18095 15861 18107 15864
rect 18049 15855 18107 15861
rect 18138 15852 18144 15864
rect 18196 15852 18202 15904
rect 21637 15895 21695 15901
rect 21637 15861 21649 15895
rect 21683 15892 21695 15895
rect 23290 15892 23296 15904
rect 21683 15864 23296 15892
rect 21683 15861 21695 15864
rect 21637 15855 21695 15861
rect 23290 15852 23296 15864
rect 23348 15852 23354 15904
rect 24026 15892 24032 15904
rect 23987 15864 24032 15892
rect 24026 15852 24032 15864
rect 24084 15852 24090 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2133 15691 2191 15697
rect 2133 15657 2145 15691
rect 2179 15688 2191 15691
rect 2498 15688 2504 15700
rect 2179 15660 2504 15688
rect 2179 15657 2191 15660
rect 2133 15651 2191 15657
rect 2498 15648 2504 15660
rect 2556 15688 2562 15700
rect 3418 15688 3424 15700
rect 2556 15660 3424 15688
rect 2556 15648 2562 15660
rect 3418 15648 3424 15660
rect 3476 15648 3482 15700
rect 3878 15688 3884 15700
rect 3839 15660 3884 15688
rect 3878 15648 3884 15660
rect 3936 15688 3942 15700
rect 3936 15660 5580 15688
rect 3936 15648 3942 15660
rect 2777 15623 2835 15629
rect 2777 15589 2789 15623
rect 2823 15620 2835 15623
rect 4062 15620 4068 15632
rect 2823 15592 4068 15620
rect 2823 15589 2835 15592
rect 2777 15583 2835 15589
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 2406 15552 2412 15564
rect 1443 15524 2412 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 2406 15512 2412 15524
rect 2464 15512 2470 15564
rect 2682 15512 2688 15564
rect 2740 15552 2746 15564
rect 2792 15552 2820 15583
rect 4062 15580 4068 15592
rect 4120 15580 4126 15632
rect 4617 15623 4675 15629
rect 4617 15589 4629 15623
rect 4663 15620 4675 15623
rect 4976 15623 5034 15629
rect 4976 15620 4988 15623
rect 4663 15592 4988 15620
rect 4663 15589 4675 15592
rect 4617 15583 4675 15589
rect 4976 15589 4988 15592
rect 5022 15620 5034 15623
rect 5442 15620 5448 15632
rect 5022 15592 5448 15620
rect 5022 15589 5034 15592
rect 4976 15583 5034 15589
rect 5442 15580 5448 15592
rect 5500 15580 5506 15632
rect 5552 15620 5580 15660
rect 5626 15648 5632 15700
rect 5684 15688 5690 15700
rect 8021 15691 8079 15697
rect 8021 15688 8033 15691
rect 5684 15660 8033 15688
rect 5684 15648 5690 15660
rect 8021 15657 8033 15660
rect 8067 15688 8079 15691
rect 10597 15691 10655 15697
rect 10597 15688 10609 15691
rect 8067 15660 10609 15688
rect 8067 15657 8079 15660
rect 8021 15651 8079 15657
rect 10597 15657 10609 15660
rect 10643 15657 10655 15691
rect 12158 15688 12164 15700
rect 12119 15660 12164 15688
rect 10597 15651 10655 15657
rect 12158 15648 12164 15660
rect 12216 15648 12222 15700
rect 12805 15691 12863 15697
rect 12805 15657 12817 15691
rect 12851 15688 12863 15691
rect 13078 15688 13084 15700
rect 12851 15660 13084 15688
rect 12851 15657 12863 15660
rect 12805 15651 12863 15657
rect 13078 15648 13084 15660
rect 13136 15688 13142 15700
rect 13354 15688 13360 15700
rect 13136 15660 13360 15688
rect 13136 15648 13142 15660
rect 13354 15648 13360 15660
rect 13412 15648 13418 15700
rect 13538 15648 13544 15700
rect 13596 15688 13602 15700
rect 13633 15691 13691 15697
rect 13633 15688 13645 15691
rect 13596 15660 13645 15688
rect 13596 15648 13602 15660
rect 13633 15657 13645 15660
rect 13679 15688 13691 15691
rect 13722 15688 13728 15700
rect 13679 15660 13728 15688
rect 13679 15657 13691 15660
rect 13633 15651 13691 15657
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 14274 15688 14280 15700
rect 14235 15660 14280 15688
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 14642 15688 14648 15700
rect 14603 15660 14648 15688
rect 14642 15648 14648 15660
rect 14700 15648 14706 15700
rect 17129 15691 17187 15697
rect 17129 15657 17141 15691
rect 17175 15688 17187 15691
rect 17402 15688 17408 15700
rect 17175 15660 17408 15688
rect 17175 15657 17187 15660
rect 17129 15651 17187 15657
rect 17402 15648 17408 15660
rect 17460 15648 17466 15700
rect 18046 15648 18052 15700
rect 18104 15688 18110 15700
rect 18414 15688 18420 15700
rect 18104 15660 18420 15688
rect 18104 15648 18110 15660
rect 18414 15648 18420 15660
rect 18472 15688 18478 15700
rect 18693 15691 18751 15697
rect 18693 15688 18705 15691
rect 18472 15660 18705 15688
rect 18472 15648 18478 15660
rect 18693 15657 18705 15660
rect 18739 15657 18751 15691
rect 19334 15688 19340 15700
rect 19295 15660 19340 15688
rect 18693 15651 18751 15657
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 20346 15688 20352 15700
rect 20307 15660 20352 15688
rect 20346 15648 20352 15660
rect 20404 15648 20410 15700
rect 20622 15688 20628 15700
rect 20583 15660 20628 15688
rect 20622 15648 20628 15660
rect 20680 15648 20686 15700
rect 20901 15691 20959 15697
rect 20901 15657 20913 15691
rect 20947 15688 20959 15691
rect 21266 15688 21272 15700
rect 20947 15660 21272 15688
rect 20947 15657 20959 15660
rect 20901 15651 20959 15657
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 21361 15691 21419 15697
rect 21361 15657 21373 15691
rect 21407 15688 21419 15691
rect 21542 15688 21548 15700
rect 21407 15660 21548 15688
rect 21407 15657 21419 15660
rect 21361 15651 21419 15657
rect 6641 15623 6699 15629
rect 6641 15620 6653 15623
rect 5552 15592 6653 15620
rect 6641 15589 6653 15592
rect 6687 15620 6699 15623
rect 6730 15620 6736 15632
rect 6687 15592 6736 15620
rect 6687 15589 6699 15592
rect 6641 15583 6699 15589
rect 6730 15580 6736 15592
rect 6788 15580 6794 15632
rect 7101 15623 7159 15629
rect 7101 15589 7113 15623
rect 7147 15620 7159 15623
rect 7466 15620 7472 15632
rect 7147 15592 7472 15620
rect 7147 15589 7159 15592
rect 7101 15583 7159 15589
rect 7466 15580 7472 15592
rect 7524 15580 7530 15632
rect 8110 15580 8116 15632
rect 8168 15620 8174 15632
rect 8386 15620 8392 15632
rect 8168 15592 8392 15620
rect 8168 15580 8174 15592
rect 8386 15580 8392 15592
rect 8444 15580 8450 15632
rect 9858 15580 9864 15632
rect 9916 15620 9922 15632
rect 10229 15623 10287 15629
rect 10229 15620 10241 15623
rect 9916 15592 10241 15620
rect 9916 15580 9922 15592
rect 10229 15589 10241 15592
rect 10275 15589 10287 15623
rect 10229 15583 10287 15589
rect 11048 15623 11106 15629
rect 11048 15589 11060 15623
rect 11094 15620 11106 15623
rect 11146 15620 11152 15632
rect 11094 15592 11152 15620
rect 11094 15589 11106 15592
rect 11048 15583 11106 15589
rect 11146 15580 11152 15592
rect 11204 15580 11210 15632
rect 13173 15623 13231 15629
rect 13173 15589 13185 15623
rect 13219 15620 13231 15623
rect 13262 15620 13268 15632
rect 13219 15592 13268 15620
rect 13219 15589 13231 15592
rect 13173 15583 13231 15589
rect 13262 15580 13268 15592
rect 13320 15620 13326 15632
rect 13320 15592 17908 15620
rect 13320 15580 13326 15592
rect 2740 15524 2820 15552
rect 2740 15512 2746 15524
rect 4338 15512 4344 15564
rect 4396 15552 4402 15564
rect 4709 15555 4767 15561
rect 4709 15552 4721 15555
rect 4396 15524 4721 15552
rect 4396 15512 4402 15524
rect 4709 15521 4721 15524
rect 4755 15552 4767 15555
rect 4798 15552 4804 15564
rect 4755 15524 4804 15552
rect 4755 15521 4767 15524
rect 4709 15515 4767 15521
rect 4798 15512 4804 15524
rect 4856 15552 4862 15564
rect 6546 15552 6552 15564
rect 4856 15524 6552 15552
rect 4856 15512 4862 15524
rect 6546 15512 6552 15524
rect 6604 15512 6610 15564
rect 8294 15512 8300 15564
rect 8352 15552 8358 15564
rect 8481 15555 8539 15561
rect 8481 15552 8493 15555
rect 8352 15524 8493 15552
rect 8352 15512 8358 15524
rect 8481 15521 8493 15524
rect 8527 15521 8539 15555
rect 8481 15515 8539 15521
rect 9677 15555 9735 15561
rect 9677 15521 9689 15555
rect 9723 15552 9735 15555
rect 10686 15552 10692 15564
rect 9723 15524 10692 15552
rect 9723 15521 9735 15524
rect 9677 15515 9735 15521
rect 10686 15512 10692 15524
rect 10744 15512 10750 15564
rect 10781 15555 10839 15561
rect 10781 15521 10793 15555
rect 10827 15552 10839 15555
rect 10870 15552 10876 15564
rect 10827 15524 10876 15552
rect 10827 15521 10839 15524
rect 10781 15515 10839 15521
rect 10870 15512 10876 15524
rect 10928 15512 10934 15564
rect 15562 15512 15568 15564
rect 15620 15552 15626 15564
rect 16016 15555 16074 15561
rect 16016 15552 16028 15555
rect 15620 15524 16028 15552
rect 15620 15512 15626 15524
rect 16016 15521 16028 15524
rect 16062 15552 16074 15555
rect 16390 15552 16396 15564
rect 16062 15524 16396 15552
rect 16062 15521 16074 15524
rect 16016 15515 16074 15521
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 1578 15444 1584 15496
rect 1636 15484 1642 15496
rect 2038 15484 2044 15496
rect 1636 15456 2044 15484
rect 1636 15444 1642 15456
rect 2038 15444 2044 15456
rect 2096 15444 2102 15496
rect 2498 15444 2504 15496
rect 2556 15484 2562 15496
rect 2869 15487 2927 15493
rect 2869 15484 2881 15487
rect 2556 15456 2881 15484
rect 2556 15444 2562 15456
rect 2869 15453 2881 15456
rect 2915 15453 2927 15487
rect 2869 15447 2927 15453
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 3099 15456 3556 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 2774 15376 2780 15428
rect 2832 15416 2838 15428
rect 3068 15416 3096 15447
rect 2832 15388 3096 15416
rect 2832 15376 2838 15388
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 2406 15348 2412 15360
rect 2367 15320 2412 15348
rect 2406 15308 2412 15320
rect 2464 15308 2470 15360
rect 3528 15357 3556 15456
rect 8570 15444 8576 15496
rect 8628 15484 8634 15496
rect 8849 15487 8907 15493
rect 8628 15456 8673 15484
rect 8628 15444 8634 15456
rect 8849 15453 8861 15487
rect 8895 15484 8907 15487
rect 9401 15487 9459 15493
rect 9401 15484 9413 15487
rect 8895 15456 9413 15484
rect 8895 15453 8907 15456
rect 8849 15447 8907 15453
rect 9401 15453 9413 15456
rect 9447 15453 9459 15487
rect 9401 15447 9459 15453
rect 13538 15444 13544 15496
rect 13596 15484 13602 15496
rect 13725 15487 13783 15493
rect 13725 15484 13737 15487
rect 13596 15456 13737 15484
rect 13596 15444 13602 15456
rect 13725 15453 13737 15456
rect 13771 15453 13783 15487
rect 13906 15484 13912 15496
rect 13867 15456 13912 15484
rect 13725 15447 13783 15453
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 15102 15484 15108 15496
rect 15063 15456 15108 15484
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 15749 15487 15807 15493
rect 15749 15484 15761 15487
rect 15488 15456 15761 15484
rect 6086 15416 6092 15428
rect 6047 15388 6092 15416
rect 6086 15376 6092 15388
rect 6144 15416 6150 15428
rect 7377 15419 7435 15425
rect 7377 15416 7389 15419
rect 6144 15388 7389 15416
rect 6144 15376 6150 15388
rect 7377 15385 7389 15388
rect 7423 15385 7435 15419
rect 7742 15416 7748 15428
rect 7703 15388 7748 15416
rect 7377 15379 7435 15385
rect 7742 15376 7748 15388
rect 7800 15376 7806 15428
rect 8478 15376 8484 15428
rect 8536 15416 8542 15428
rect 9306 15416 9312 15428
rect 8536 15388 9312 15416
rect 8536 15376 8542 15388
rect 9306 15376 9312 15388
rect 9364 15376 9370 15428
rect 9674 15376 9680 15428
rect 9732 15416 9738 15428
rect 9861 15419 9919 15425
rect 9861 15416 9873 15419
rect 9732 15388 9873 15416
rect 9732 15376 9738 15388
rect 9861 15385 9873 15388
rect 9907 15385 9919 15419
rect 9861 15379 9919 15385
rect 15488 15360 15516 15456
rect 15749 15453 15761 15456
rect 15795 15453 15807 15487
rect 17880 15484 17908 15592
rect 19242 15580 19248 15632
rect 19300 15620 19306 15632
rect 19705 15623 19763 15629
rect 19705 15620 19717 15623
rect 19300 15592 19717 15620
rect 19300 15580 19306 15592
rect 19705 15589 19717 15592
rect 19751 15620 19763 15623
rect 20990 15620 20996 15632
rect 19751 15592 20996 15620
rect 19751 15589 19763 15592
rect 19705 15583 19763 15589
rect 20990 15580 20996 15592
rect 21048 15580 21054 15632
rect 21174 15580 21180 15632
rect 21232 15620 21238 15632
rect 21376 15620 21404 15651
rect 21542 15648 21548 15660
rect 21600 15648 21606 15700
rect 22005 15691 22063 15697
rect 22005 15657 22017 15691
rect 22051 15688 22063 15691
rect 22094 15688 22100 15700
rect 22051 15660 22100 15688
rect 22051 15657 22063 15660
rect 22005 15651 22063 15657
rect 22094 15648 22100 15660
rect 22152 15648 22158 15700
rect 22186 15648 22192 15700
rect 22244 15688 22250 15700
rect 22281 15691 22339 15697
rect 22281 15688 22293 15691
rect 22244 15660 22293 15688
rect 22244 15648 22250 15660
rect 22281 15657 22293 15660
rect 22327 15657 22339 15691
rect 22281 15651 22339 15657
rect 24026 15648 24032 15700
rect 24084 15688 24090 15700
rect 24765 15691 24823 15697
rect 24765 15688 24777 15691
rect 24084 15660 24777 15688
rect 24084 15648 24090 15660
rect 24765 15657 24777 15660
rect 24811 15657 24823 15691
rect 24765 15651 24823 15657
rect 25133 15691 25191 15697
rect 25133 15657 25145 15691
rect 25179 15688 25191 15691
rect 25222 15688 25228 15700
rect 25179 15660 25228 15688
rect 25179 15657 25191 15660
rect 25133 15651 25191 15657
rect 25222 15648 25228 15660
rect 25280 15648 25286 15700
rect 25498 15620 25504 15632
rect 21232 15592 21404 15620
rect 25459 15592 25504 15620
rect 21232 15580 21238 15592
rect 25498 15580 25504 15592
rect 25556 15580 25562 15632
rect 17954 15512 17960 15564
rect 18012 15552 18018 15564
rect 18601 15555 18659 15561
rect 18601 15552 18613 15555
rect 18012 15524 18613 15552
rect 18012 15512 18018 15524
rect 18601 15521 18613 15524
rect 18647 15521 18659 15555
rect 18601 15515 18659 15521
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 19518 15552 19524 15564
rect 19392 15524 19524 15552
rect 19392 15512 19398 15524
rect 19518 15512 19524 15524
rect 19576 15512 19582 15564
rect 19797 15555 19855 15561
rect 19797 15521 19809 15555
rect 19843 15552 19855 15555
rect 21269 15555 21327 15561
rect 21269 15552 21281 15555
rect 19843 15524 21281 15552
rect 19843 15521 19855 15524
rect 19797 15515 19855 15521
rect 21269 15521 21281 15524
rect 21315 15552 21327 15555
rect 21910 15552 21916 15564
rect 21315 15524 21916 15552
rect 21315 15521 21327 15524
rect 21269 15515 21327 15521
rect 21910 15512 21916 15524
rect 21968 15512 21974 15564
rect 22370 15512 22376 15564
rect 22428 15552 22434 15564
rect 22721 15555 22779 15561
rect 22721 15552 22733 15555
rect 22428 15524 22733 15552
rect 22428 15512 22434 15524
rect 22721 15521 22733 15524
rect 22767 15521 22779 15555
rect 24946 15552 24952 15564
rect 24907 15524 24952 15552
rect 22721 15515 22779 15521
rect 24946 15512 24952 15524
rect 25004 15512 25010 15564
rect 18782 15484 18788 15496
rect 17880 15456 18460 15484
rect 18743 15456 18788 15484
rect 15749 15447 15807 15453
rect 18230 15416 18236 15428
rect 18191 15388 18236 15416
rect 18230 15376 18236 15388
rect 18288 15376 18294 15428
rect 18432 15416 18460 15456
rect 18782 15444 18788 15456
rect 18840 15444 18846 15496
rect 20622 15444 20628 15496
rect 20680 15484 20686 15496
rect 21453 15487 21511 15493
rect 21453 15484 21465 15487
rect 20680 15456 21465 15484
rect 20680 15444 20686 15456
rect 21453 15453 21465 15456
rect 21499 15453 21511 15487
rect 22462 15484 22468 15496
rect 22423 15456 22468 15484
rect 21453 15447 21511 15453
rect 22462 15444 22468 15456
rect 22520 15444 22526 15496
rect 20990 15416 20996 15428
rect 18432 15388 20996 15416
rect 20990 15376 20996 15388
rect 21048 15376 21054 15428
rect 21100 15388 22232 15416
rect 3513 15351 3571 15357
rect 3513 15317 3525 15351
rect 3559 15348 3571 15351
rect 3694 15348 3700 15360
rect 3559 15320 3700 15348
rect 3559 15317 3571 15320
rect 3513 15311 3571 15317
rect 3694 15308 3700 15320
rect 3752 15308 3758 15360
rect 3970 15308 3976 15360
rect 4028 15348 4034 15360
rect 8849 15351 8907 15357
rect 8849 15348 8861 15351
rect 4028 15320 8861 15348
rect 4028 15308 4034 15320
rect 8849 15317 8861 15320
rect 8895 15317 8907 15351
rect 9030 15348 9036 15360
rect 8991 15320 9036 15348
rect 8849 15311 8907 15317
rect 9030 15308 9036 15320
rect 9088 15308 9094 15360
rect 13265 15351 13323 15357
rect 13265 15317 13277 15351
rect 13311 15348 13323 15351
rect 14090 15348 14096 15360
rect 13311 15320 14096 15348
rect 13311 15317 13323 15320
rect 13265 15311 13323 15317
rect 14090 15308 14096 15320
rect 14148 15308 14154 15360
rect 15470 15348 15476 15360
rect 15431 15320 15476 15348
rect 15470 15308 15476 15320
rect 15528 15308 15534 15360
rect 15562 15308 15568 15360
rect 15620 15348 15626 15360
rect 17310 15348 17316 15360
rect 15620 15320 17316 15348
rect 15620 15308 15626 15320
rect 17310 15308 17316 15320
rect 17368 15308 17374 15360
rect 17494 15308 17500 15360
rect 17552 15348 17558 15360
rect 17681 15351 17739 15357
rect 17681 15348 17693 15351
rect 17552 15320 17693 15348
rect 17552 15308 17558 15320
rect 17681 15317 17693 15320
rect 17727 15317 17739 15351
rect 17681 15311 17739 15317
rect 18141 15351 18199 15357
rect 18141 15317 18153 15351
rect 18187 15348 18199 15351
rect 18598 15348 18604 15360
rect 18187 15320 18604 15348
rect 18187 15317 18199 15320
rect 18141 15311 18199 15317
rect 18598 15308 18604 15320
rect 18656 15308 18662 15360
rect 19886 15308 19892 15360
rect 19944 15348 19950 15360
rect 21100 15348 21128 15388
rect 19944 15320 21128 15348
rect 19944 15308 19950 15320
rect 21634 15308 21640 15360
rect 21692 15348 21698 15360
rect 21818 15348 21824 15360
rect 21692 15320 21824 15348
rect 21692 15308 21698 15320
rect 21818 15308 21824 15320
rect 21876 15308 21882 15360
rect 22204 15348 22232 15388
rect 22830 15348 22836 15360
rect 22204 15320 22836 15348
rect 22830 15308 22836 15320
rect 22888 15308 22894 15360
rect 23474 15308 23480 15360
rect 23532 15348 23538 15360
rect 23845 15351 23903 15357
rect 23845 15348 23857 15351
rect 23532 15320 23857 15348
rect 23532 15308 23538 15320
rect 23845 15317 23857 15320
rect 23891 15317 23903 15351
rect 23845 15311 23903 15317
rect 24118 15308 24124 15360
rect 24176 15348 24182 15360
rect 24397 15351 24455 15357
rect 24397 15348 24409 15351
rect 24176 15320 24409 15348
rect 24176 15308 24182 15320
rect 24397 15317 24409 15320
rect 24443 15317 24455 15351
rect 24397 15311 24455 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1949 15147 2007 15153
rect 1949 15113 1961 15147
rect 1995 15144 2007 15147
rect 2682 15144 2688 15156
rect 1995 15116 2688 15144
rect 1995 15113 2007 15116
rect 1949 15107 2007 15113
rect 2682 15104 2688 15116
rect 2740 15104 2746 15156
rect 7009 15147 7067 15153
rect 7009 15113 7021 15147
rect 7055 15144 7067 15147
rect 7190 15144 7196 15156
rect 7055 15116 7196 15144
rect 7055 15113 7067 15116
rect 7009 15107 7067 15113
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 8110 15144 8116 15156
rect 8071 15116 8116 15144
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 8389 15147 8447 15153
rect 8389 15144 8401 15147
rect 8352 15116 8401 15144
rect 8352 15104 8358 15116
rect 8389 15113 8401 15116
rect 8435 15144 8447 15147
rect 9306 15144 9312 15156
rect 8435 15116 9312 15144
rect 8435 15113 8447 15116
rect 8389 15107 8447 15113
rect 9306 15104 9312 15116
rect 9364 15104 9370 15156
rect 10870 15144 10876 15156
rect 10831 15116 10876 15144
rect 10870 15104 10876 15116
rect 10928 15144 10934 15156
rect 11698 15144 11704 15156
rect 10928 15116 11704 15144
rect 10928 15104 10934 15116
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 12713 15147 12771 15153
rect 12713 15113 12725 15147
rect 12759 15144 12771 15147
rect 13722 15144 13728 15156
rect 12759 15116 13728 15144
rect 12759 15113 12771 15116
rect 12713 15107 12771 15113
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 14458 15144 14464 15156
rect 14419 15116 14464 15144
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 17218 15104 17224 15156
rect 17276 15144 17282 15156
rect 17405 15147 17463 15153
rect 17405 15144 17417 15147
rect 17276 15116 17417 15144
rect 17276 15104 17282 15116
rect 17405 15113 17417 15116
rect 17451 15144 17463 15147
rect 17862 15144 17868 15156
rect 17451 15116 17868 15144
rect 17451 15113 17463 15116
rect 17405 15107 17463 15113
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 19521 15147 19579 15153
rect 19521 15113 19533 15147
rect 19567 15144 19579 15147
rect 20254 15144 20260 15156
rect 19567 15116 20260 15144
rect 19567 15113 19579 15116
rect 19521 15107 19579 15113
rect 20254 15104 20260 15116
rect 20312 15104 20318 15156
rect 21910 15144 21916 15156
rect 21871 15116 21916 15144
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 22094 15104 22100 15156
rect 22152 15144 22158 15156
rect 22462 15144 22468 15156
rect 22152 15116 22468 15144
rect 22152 15104 22158 15116
rect 22462 15104 22468 15116
rect 22520 15104 22526 15156
rect 22554 15104 22560 15156
rect 22612 15144 22618 15156
rect 24946 15144 24952 15156
rect 22612 15116 24952 15144
rect 22612 15104 22618 15116
rect 24946 15104 24952 15116
rect 25004 15104 25010 15156
rect 25409 15147 25467 15153
rect 25409 15113 25421 15147
rect 25455 15144 25467 15147
rect 25958 15144 25964 15156
rect 25455 15116 25964 15144
rect 25455 15113 25467 15116
rect 25409 15107 25467 15113
rect 25958 15104 25964 15116
rect 26016 15104 26022 15156
rect 2409 15079 2467 15085
rect 2409 15045 2421 15079
rect 2455 15076 2467 15079
rect 2774 15076 2780 15088
rect 2455 15048 2780 15076
rect 2455 15045 2467 15048
rect 2409 15039 2467 15045
rect 2774 15036 2780 15048
rect 2832 15036 2838 15088
rect 3970 15076 3976 15088
rect 2884 15048 3976 15076
rect 1486 14968 1492 15020
rect 1544 15008 1550 15020
rect 1762 15008 1768 15020
rect 1544 14980 1768 15008
rect 1544 14968 1550 14980
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 2314 14968 2320 15020
rect 2372 15008 2378 15020
rect 2884 15017 2912 15048
rect 3970 15036 3976 15048
rect 4028 15036 4034 15088
rect 5997 15079 6055 15085
rect 5997 15045 6009 15079
rect 6043 15076 6055 15079
rect 6546 15076 6552 15088
rect 6043 15048 6552 15076
rect 6043 15045 6055 15048
rect 5997 15039 6055 15045
rect 6546 15036 6552 15048
rect 6604 15076 6610 15088
rect 6604 15048 8616 15076
rect 6604 15036 6610 15048
rect 2869 15011 2927 15017
rect 2869 15008 2881 15011
rect 2372 14980 2881 15008
rect 2372 14968 2378 14980
rect 2869 14977 2881 14980
rect 2915 14977 2927 15011
rect 2869 14971 2927 14977
rect 3053 15011 3111 15017
rect 3053 14977 3065 15011
rect 3099 15008 3111 15011
rect 3602 15008 3608 15020
rect 3099 14980 3608 15008
rect 3099 14977 3111 14980
rect 3053 14971 3111 14977
rect 3602 14968 3608 14980
rect 3660 14968 3666 15020
rect 7558 15008 7564 15020
rect 7519 14980 7564 15008
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 1946 14940 1952 14952
rect 1443 14912 1952 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 1946 14900 1952 14912
rect 2004 14900 2010 14952
rect 2777 14943 2835 14949
rect 2777 14909 2789 14943
rect 2823 14940 2835 14943
rect 3142 14940 3148 14952
rect 2823 14912 3148 14940
rect 2823 14909 2835 14912
rect 2777 14903 2835 14909
rect 3142 14900 3148 14912
rect 3200 14900 3206 14952
rect 3881 14943 3939 14949
rect 3881 14909 3893 14943
rect 3927 14940 3939 14943
rect 3973 14943 4031 14949
rect 3973 14940 3985 14943
rect 3927 14912 3985 14940
rect 3927 14909 3939 14912
rect 3881 14903 3939 14909
rect 3973 14909 3985 14912
rect 4019 14940 4031 14943
rect 4019 14912 4384 14940
rect 4019 14909 4031 14912
rect 3973 14903 4031 14909
rect 4356 14884 4384 14912
rect 4614 14900 4620 14952
rect 4672 14940 4678 14952
rect 7190 14940 7196 14952
rect 4672 14912 7196 14940
rect 4672 14900 4678 14912
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 7469 14943 7527 14949
rect 7469 14909 7481 14943
rect 7515 14940 7527 14943
rect 7742 14940 7748 14952
rect 7515 14912 7748 14940
rect 7515 14909 7527 14912
rect 7469 14903 7527 14909
rect 4246 14881 4252 14884
rect 4240 14872 4252 14881
rect 4207 14844 4252 14872
rect 4240 14835 4252 14844
rect 4246 14832 4252 14835
rect 4304 14832 4310 14884
rect 4338 14832 4344 14884
rect 4396 14832 4402 14884
rect 6641 14875 6699 14881
rect 6641 14841 6653 14875
rect 6687 14872 6699 14875
rect 7484 14872 7512 14903
rect 7742 14900 7748 14912
rect 7800 14900 7806 14952
rect 8588 14949 8616 15048
rect 10134 15036 10140 15088
rect 10192 15076 10198 15088
rect 11238 15076 11244 15088
rect 10192 15048 11244 15076
rect 10192 15036 10198 15048
rect 11238 15036 11244 15048
rect 11296 15036 11302 15088
rect 11716 15076 11744 15104
rect 14185 15079 14243 15085
rect 11716 15048 14136 15076
rect 11054 15008 11060 15020
rect 11015 14980 11060 15008
rect 11054 14968 11060 14980
rect 11112 14968 11118 15020
rect 13265 15011 13323 15017
rect 13265 15008 13277 15011
rect 12452 14980 13277 15008
rect 8573 14943 8631 14949
rect 8573 14909 8585 14943
rect 8619 14940 8631 14943
rect 9582 14940 9588 14952
rect 8619 14912 9588 14940
rect 8619 14909 8631 14912
rect 8573 14903 8631 14909
rect 9582 14900 9588 14912
rect 9640 14900 9646 14952
rect 10134 14900 10140 14952
rect 10192 14940 10198 14952
rect 10594 14940 10600 14952
rect 10192 14912 10600 14940
rect 10192 14900 10198 14912
rect 10594 14900 10600 14912
rect 10652 14900 10658 14952
rect 12452 14940 12480 14980
rect 13265 14977 13277 14980
rect 13311 14977 13323 15011
rect 14108 15008 14136 15048
rect 14185 15045 14197 15079
rect 14231 15076 14243 15079
rect 14642 15076 14648 15088
rect 14231 15048 14648 15076
rect 14231 15045 14243 15048
rect 14185 15039 14243 15045
rect 14642 15036 14648 15048
rect 14700 15036 14706 15088
rect 17788 15048 18644 15076
rect 15289 15011 15347 15017
rect 15289 15008 15301 15011
rect 14108 14980 15301 15008
rect 13265 14971 13323 14977
rect 15289 14977 15301 14980
rect 15335 15008 15347 15011
rect 15470 15008 15476 15020
rect 15335 14980 15476 15008
rect 15335 14977 15347 14980
rect 15289 14971 15347 14977
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 17402 14968 17408 15020
rect 17460 15008 17466 15020
rect 17788 15017 17816 15048
rect 17773 15011 17831 15017
rect 17773 15008 17785 15011
rect 17460 14980 17785 15008
rect 17460 14968 17466 14980
rect 17773 14977 17785 14980
rect 17819 14977 17831 15011
rect 18506 15008 18512 15020
rect 18467 14980 18512 15008
rect 17773 14971 17831 14977
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 18616 15017 18644 15048
rect 18782 15036 18788 15088
rect 18840 15076 18846 15088
rect 18877 15079 18935 15085
rect 18877 15076 18889 15079
rect 18840 15048 18889 15076
rect 18840 15036 18846 15048
rect 18877 15045 18889 15048
rect 18923 15045 18935 15079
rect 22370 15076 22376 15088
rect 22331 15048 22376 15076
rect 18877 15039 18935 15045
rect 22370 15036 22376 15048
rect 22428 15036 22434 15088
rect 22738 15036 22744 15088
rect 22796 15076 22802 15088
rect 23017 15079 23075 15085
rect 23017 15076 23029 15079
rect 22796 15048 23029 15076
rect 22796 15036 22802 15048
rect 23017 15045 23029 15048
rect 23063 15045 23075 15079
rect 23017 15039 23075 15045
rect 24026 15036 24032 15088
rect 24084 15076 24090 15088
rect 26234 15076 26240 15088
rect 24084 15048 24900 15076
rect 26195 15048 26240 15076
rect 24084 15036 24090 15048
rect 18601 15011 18659 15017
rect 18601 14977 18613 15011
rect 18647 14977 18659 15011
rect 24118 15008 24124 15020
rect 24079 14980 24124 15008
rect 18601 14971 18659 14977
rect 24118 14968 24124 14980
rect 24176 14968 24182 15020
rect 24213 15011 24271 15017
rect 24213 14977 24225 15011
rect 24259 14977 24271 15011
rect 24213 14971 24271 14977
rect 13078 14940 13084 14952
rect 12268 14912 12480 14940
rect 13039 14912 13084 14940
rect 6687 14844 7512 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 8386 14832 8392 14884
rect 8444 14872 8450 14884
rect 8818 14875 8876 14881
rect 8818 14872 8830 14875
rect 8444 14844 8830 14872
rect 8444 14832 8450 14844
rect 8818 14841 8830 14844
rect 8864 14872 8876 14875
rect 9030 14872 9036 14884
rect 8864 14844 9036 14872
rect 8864 14841 8876 14844
rect 8818 14835 8876 14841
rect 9030 14832 9036 14844
rect 9088 14832 9094 14884
rect 12268 14816 12296 14912
rect 13078 14900 13084 14912
rect 13136 14900 13142 14952
rect 13173 14943 13231 14949
rect 13173 14909 13185 14943
rect 13219 14940 13231 14943
rect 13446 14940 13452 14952
rect 13219 14912 13452 14940
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 13446 14900 13452 14912
rect 13504 14900 13510 14952
rect 13998 14900 14004 14952
rect 14056 14940 14062 14952
rect 14277 14943 14335 14949
rect 14277 14940 14289 14943
rect 14056 14912 14289 14940
rect 14056 14900 14062 14912
rect 14277 14909 14289 14912
rect 14323 14940 14335 14943
rect 14918 14940 14924 14952
rect 14323 14912 14924 14940
rect 14323 14909 14335 14912
rect 14277 14903 14335 14909
rect 14918 14900 14924 14912
rect 14976 14900 14982 14952
rect 17034 14900 17040 14952
rect 17092 14940 17098 14952
rect 19886 14940 19892 14952
rect 17092 14912 19892 14940
rect 17092 14900 17098 14912
rect 19886 14900 19892 14912
rect 19944 14900 19950 14952
rect 19981 14943 20039 14949
rect 19981 14909 19993 14943
rect 20027 14909 20039 14943
rect 19981 14903 20039 14909
rect 15746 14881 15752 14884
rect 15013 14875 15071 14881
rect 15013 14841 15025 14875
rect 15059 14872 15071 14875
rect 15740 14872 15752 14881
rect 15059 14844 15752 14872
rect 15059 14841 15071 14844
rect 15013 14835 15071 14841
rect 15740 14835 15752 14844
rect 15746 14832 15752 14835
rect 15804 14832 15810 14884
rect 17862 14832 17868 14884
rect 17920 14872 17926 14884
rect 18877 14875 18935 14881
rect 18877 14872 18889 14875
rect 17920 14844 18889 14872
rect 17920 14832 17926 14844
rect 18877 14841 18889 14844
rect 18923 14872 18935 14875
rect 19061 14875 19119 14881
rect 19061 14872 19073 14875
rect 18923 14844 19073 14872
rect 18923 14841 18935 14844
rect 18877 14835 18935 14841
rect 19061 14841 19073 14844
rect 19107 14841 19119 14875
rect 19996 14872 20024 14903
rect 22186 14900 22192 14952
rect 22244 14940 22250 14952
rect 22465 14943 22523 14949
rect 22465 14940 22477 14943
rect 22244 14912 22477 14940
rect 22244 14900 22250 14912
rect 22465 14909 22477 14912
rect 22511 14909 22523 14943
rect 23474 14940 23480 14952
rect 23435 14912 23480 14940
rect 22465 14903 22523 14909
rect 23474 14900 23480 14912
rect 23532 14940 23538 14952
rect 24228 14940 24256 14971
rect 23532 14912 24256 14940
rect 24872 14940 24900 15048
rect 26234 15036 26240 15048
rect 26292 15036 26298 15088
rect 25225 14943 25283 14949
rect 25225 14940 25237 14943
rect 24872 14912 25237 14940
rect 23532 14900 23538 14912
rect 25225 14909 25237 14912
rect 25271 14940 25283 14943
rect 25777 14943 25835 14949
rect 25777 14940 25789 14943
rect 25271 14912 25789 14940
rect 25271 14909 25283 14912
rect 25225 14903 25283 14909
rect 25777 14909 25789 14912
rect 25823 14909 25835 14943
rect 25777 14903 25835 14909
rect 20254 14881 20260 14884
rect 20248 14872 20260 14881
rect 19061 14835 19119 14841
rect 19812 14844 20024 14872
rect 20215 14844 20260 14872
rect 1486 14764 1492 14816
rect 1544 14804 1550 14816
rect 1581 14807 1639 14813
rect 1581 14804 1593 14807
rect 1544 14776 1593 14804
rect 1544 14764 1550 14776
rect 1581 14773 1593 14776
rect 1627 14773 1639 14807
rect 1581 14767 1639 14773
rect 2317 14807 2375 14813
rect 2317 14773 2329 14807
rect 2363 14804 2375 14807
rect 2498 14804 2504 14816
rect 2363 14776 2504 14804
rect 2363 14773 2375 14776
rect 2317 14767 2375 14773
rect 2498 14764 2504 14776
rect 2556 14804 2562 14816
rect 2866 14804 2872 14816
rect 2556 14776 2872 14804
rect 2556 14764 2562 14776
rect 2866 14764 2872 14776
rect 2924 14764 2930 14816
rect 3513 14807 3571 14813
rect 3513 14773 3525 14807
rect 3559 14804 3571 14807
rect 3694 14804 3700 14816
rect 3559 14776 3700 14804
rect 3559 14773 3571 14776
rect 3513 14767 3571 14773
rect 3694 14764 3700 14776
rect 3752 14804 3758 14816
rect 5166 14804 5172 14816
rect 3752 14776 5172 14804
rect 3752 14764 3758 14776
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 5350 14804 5356 14816
rect 5311 14776 5356 14804
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 6362 14804 6368 14816
rect 5500 14776 6368 14804
rect 5500 14764 5506 14776
rect 6362 14764 6368 14776
rect 6420 14764 6426 14816
rect 7377 14807 7435 14813
rect 7377 14773 7389 14807
rect 7423 14804 7435 14807
rect 7466 14804 7472 14816
rect 7423 14776 7472 14804
rect 7423 14773 7435 14776
rect 7377 14767 7435 14773
rect 7466 14764 7472 14776
rect 7524 14764 7530 14816
rect 9953 14807 10011 14813
rect 9953 14773 9965 14807
rect 9999 14804 10011 14807
rect 10042 14804 10048 14816
rect 9999 14776 10048 14804
rect 9999 14773 10011 14776
rect 9953 14767 10011 14773
rect 10042 14764 10048 14776
rect 10100 14764 10106 14816
rect 10597 14807 10655 14813
rect 10597 14773 10609 14807
rect 10643 14804 10655 14807
rect 10686 14804 10692 14816
rect 10643 14776 10692 14804
rect 10643 14773 10655 14776
rect 10597 14767 10655 14773
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 11609 14807 11667 14813
rect 11609 14804 11621 14807
rect 11204 14776 11621 14804
rect 11204 14764 11210 14776
rect 11609 14773 11621 14776
rect 11655 14804 11667 14807
rect 12250 14804 12256 14816
rect 11655 14776 12256 14804
rect 11655 14773 11667 14776
rect 11609 14767 11667 14773
rect 12250 14764 12256 14776
rect 12308 14764 12314 14816
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 13170 14804 13176 14816
rect 12676 14776 13176 14804
rect 12676 14764 12682 14776
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 13814 14804 13820 14816
rect 13775 14776 13820 14804
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 16850 14804 16856 14816
rect 16811 14776 16856 14804
rect 16850 14764 16856 14776
rect 16908 14764 16914 14816
rect 18046 14804 18052 14816
rect 18007 14776 18052 14804
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 18417 14807 18475 14813
rect 18417 14773 18429 14807
rect 18463 14804 18475 14807
rect 18598 14804 18604 14816
rect 18463 14776 18604 14804
rect 18463 14773 18475 14776
rect 18417 14767 18475 14773
rect 18598 14764 18604 14776
rect 18656 14764 18662 14816
rect 18690 14764 18696 14816
rect 18748 14804 18754 14816
rect 19812 14813 19840 14844
rect 20248 14835 20260 14844
rect 20254 14832 20260 14835
rect 20312 14832 20318 14884
rect 20806 14832 20812 14884
rect 20864 14872 20870 14884
rect 21818 14872 21824 14884
rect 20864 14844 21824 14872
rect 20864 14832 20870 14844
rect 21818 14832 21824 14844
rect 21876 14832 21882 14884
rect 19797 14807 19855 14813
rect 19797 14804 19809 14807
rect 18748 14776 19809 14804
rect 18748 14764 18754 14776
rect 19797 14773 19809 14776
rect 19843 14773 19855 14807
rect 19797 14767 19855 14773
rect 20438 14764 20444 14816
rect 20496 14804 20502 14816
rect 21361 14807 21419 14813
rect 21361 14804 21373 14807
rect 20496 14776 21373 14804
rect 20496 14764 20502 14776
rect 21361 14773 21373 14776
rect 21407 14773 21419 14807
rect 22646 14804 22652 14816
rect 22607 14776 22652 14804
rect 21361 14767 21419 14773
rect 22646 14764 22652 14776
rect 22704 14764 22710 14816
rect 23658 14804 23664 14816
rect 23619 14776 23664 14804
rect 23658 14764 23664 14776
rect 23716 14764 23722 14816
rect 24026 14804 24032 14816
rect 23987 14776 24032 14804
rect 24026 14764 24032 14776
rect 24084 14764 24090 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1946 14600 1952 14612
rect 1907 14572 1952 14600
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 2406 14600 2412 14612
rect 2367 14572 2412 14600
rect 2406 14560 2412 14572
rect 2464 14560 2470 14612
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 2832 14572 2912 14600
rect 2832 14560 2838 14572
rect 2884 14541 2912 14572
rect 3050 14560 3056 14612
rect 3108 14600 3114 14612
rect 3421 14603 3479 14609
rect 3421 14600 3433 14603
rect 3108 14572 3433 14600
rect 3108 14560 3114 14572
rect 3421 14569 3433 14572
rect 3467 14569 3479 14603
rect 3421 14563 3479 14569
rect 3881 14603 3939 14609
rect 3881 14569 3893 14603
rect 3927 14600 3939 14603
rect 4246 14600 4252 14612
rect 3927 14572 4252 14600
rect 3927 14569 3939 14572
rect 3881 14563 3939 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 6178 14600 6184 14612
rect 6139 14572 6184 14600
rect 6178 14560 6184 14572
rect 6236 14560 6242 14612
rect 6914 14560 6920 14612
rect 6972 14600 6978 14612
rect 8018 14600 8024 14612
rect 6972 14572 8024 14600
rect 6972 14560 6978 14572
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 8294 14560 8300 14612
rect 8352 14600 8358 14612
rect 8389 14603 8447 14609
rect 8389 14600 8401 14603
rect 8352 14572 8401 14600
rect 8352 14560 8358 14572
rect 8389 14569 8401 14572
rect 8435 14569 8447 14603
rect 8389 14563 8447 14569
rect 10134 14560 10140 14612
rect 10192 14600 10198 14612
rect 10229 14603 10287 14609
rect 10229 14600 10241 14603
rect 10192 14572 10241 14600
rect 10192 14560 10198 14572
rect 10229 14569 10241 14572
rect 10275 14569 10287 14603
rect 10870 14600 10876 14612
rect 10831 14572 10876 14600
rect 10229 14563 10287 14569
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 13354 14600 13360 14612
rect 13315 14572 13360 14600
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 13906 14600 13912 14612
rect 13867 14572 13912 14600
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 14274 14600 14280 14612
rect 14235 14572 14280 14600
rect 14274 14560 14280 14572
rect 14332 14560 14338 14612
rect 14366 14560 14372 14612
rect 14424 14600 14430 14612
rect 15102 14600 15108 14612
rect 14424 14572 15108 14600
rect 14424 14560 14430 14572
rect 15102 14560 15108 14572
rect 15160 14560 15166 14612
rect 15746 14560 15752 14612
rect 15804 14600 15810 14612
rect 16574 14600 16580 14612
rect 15804 14572 16580 14600
rect 15804 14560 15810 14572
rect 16574 14560 16580 14572
rect 16632 14600 16638 14612
rect 17862 14600 17868 14612
rect 16632 14572 17868 14600
rect 16632 14560 16638 14572
rect 17862 14560 17868 14572
rect 17920 14560 17926 14612
rect 18414 14600 18420 14612
rect 18375 14572 18420 14600
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 19242 14600 19248 14612
rect 19203 14572 19248 14600
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 19518 14560 19524 14612
rect 19576 14600 19582 14612
rect 19613 14603 19671 14609
rect 19613 14600 19625 14603
rect 19576 14572 19625 14600
rect 19576 14560 19582 14572
rect 19613 14569 19625 14572
rect 19659 14569 19671 14603
rect 21082 14600 21088 14612
rect 21043 14572 21088 14600
rect 19613 14563 19671 14569
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 21266 14560 21272 14612
rect 21324 14600 21330 14612
rect 21453 14603 21511 14609
rect 21453 14600 21465 14603
rect 21324 14572 21465 14600
rect 21324 14560 21330 14572
rect 21453 14569 21465 14572
rect 21499 14569 21511 14603
rect 21453 14563 21511 14569
rect 22370 14560 22376 14612
rect 22428 14600 22434 14612
rect 23474 14600 23480 14612
rect 22428 14572 23480 14600
rect 22428 14560 22434 14572
rect 23474 14560 23480 14572
rect 23532 14600 23538 14612
rect 23661 14603 23719 14609
rect 23661 14600 23673 14603
rect 23532 14572 23673 14600
rect 23532 14560 23538 14572
rect 23661 14569 23673 14572
rect 23707 14569 23719 14603
rect 23661 14563 23719 14569
rect 24118 14560 24124 14612
rect 24176 14600 24182 14612
rect 24765 14603 24823 14609
rect 24765 14600 24777 14603
rect 24176 14572 24777 14600
rect 24176 14560 24182 14572
rect 24765 14569 24777 14572
rect 24811 14569 24823 14603
rect 24765 14563 24823 14569
rect 2869 14535 2927 14541
rect 2869 14501 2881 14535
rect 2915 14532 2927 14535
rect 6362 14532 6368 14544
rect 2915 14504 6368 14532
rect 2915 14501 2927 14504
rect 2869 14495 2927 14501
rect 6362 14492 6368 14504
rect 6420 14492 6426 14544
rect 7377 14535 7435 14541
rect 7377 14501 7389 14535
rect 7423 14532 7435 14535
rect 7558 14532 7564 14544
rect 7423 14504 7564 14532
rect 7423 14501 7435 14504
rect 7377 14495 7435 14501
rect 7558 14492 7564 14504
rect 7616 14532 7622 14544
rect 7837 14535 7895 14541
rect 7837 14532 7849 14535
rect 7616 14504 7849 14532
rect 7616 14492 7622 14504
rect 7837 14501 7849 14504
rect 7883 14501 7895 14535
rect 7837 14495 7895 14501
rect 8481 14535 8539 14541
rect 8481 14501 8493 14535
rect 8527 14532 8539 14535
rect 9122 14532 9128 14544
rect 8527 14504 9128 14532
rect 8527 14501 8539 14504
rect 8481 14495 8539 14501
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 1762 14464 1768 14476
rect 1443 14436 1768 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 1762 14424 1768 14436
rect 1820 14464 1826 14476
rect 1946 14464 1952 14476
rect 1820 14436 1952 14464
rect 1820 14424 1826 14436
rect 1946 14424 1952 14436
rect 2004 14424 2010 14476
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 2832 14436 2877 14464
rect 2832 14424 2838 14436
rect 4154 14424 4160 14476
rect 4212 14464 4218 14476
rect 4505 14467 4563 14473
rect 4505 14464 4517 14467
rect 4212 14436 4517 14464
rect 4212 14424 4218 14436
rect 4505 14433 4517 14436
rect 4551 14464 4563 14467
rect 5350 14464 5356 14476
rect 4551 14436 5356 14464
rect 4551 14433 4563 14436
rect 4505 14427 4563 14433
rect 5350 14424 5356 14436
rect 5408 14424 5414 14476
rect 6730 14464 6736 14476
rect 6691 14436 6736 14464
rect 6730 14424 6736 14436
rect 6788 14424 6794 14476
rect 7852 14464 7880 14495
rect 9122 14492 9128 14504
rect 9180 14492 9186 14544
rect 11885 14535 11943 14541
rect 11885 14501 11897 14535
rect 11931 14532 11943 14535
rect 12158 14532 12164 14544
rect 11931 14504 12164 14532
rect 11931 14501 11943 14504
rect 11885 14495 11943 14501
rect 12158 14492 12164 14504
rect 12216 14541 12222 14544
rect 12216 14535 12280 14541
rect 12216 14501 12234 14535
rect 12268 14501 12280 14535
rect 12216 14495 12280 14501
rect 12216 14492 12222 14495
rect 14550 14492 14556 14544
rect 14608 14532 14614 14544
rect 15930 14532 15936 14544
rect 14608 14504 15936 14532
rect 14608 14492 14614 14504
rect 15930 14492 15936 14504
rect 15988 14492 15994 14544
rect 16390 14532 16396 14544
rect 16303 14504 16396 14532
rect 16390 14492 16396 14504
rect 16448 14532 16454 14544
rect 16850 14532 16856 14544
rect 16448 14504 16856 14532
rect 16448 14492 16454 14504
rect 16850 14492 16856 14504
rect 16908 14492 16914 14544
rect 21358 14492 21364 14544
rect 21416 14532 21422 14544
rect 21913 14535 21971 14541
rect 21913 14532 21925 14535
rect 21416 14504 21925 14532
rect 21416 14492 21422 14504
rect 21913 14501 21925 14504
rect 21959 14532 21971 14535
rect 22094 14532 22100 14544
rect 21959 14504 22100 14532
rect 21959 14501 21971 14504
rect 21913 14495 21971 14501
rect 22094 14492 22100 14504
rect 22152 14492 22158 14544
rect 7852 14436 8616 14464
rect 1854 14356 1860 14408
rect 1912 14396 1918 14408
rect 2682 14396 2688 14408
rect 1912 14368 2688 14396
rect 1912 14356 1918 14368
rect 2682 14356 2688 14368
rect 2740 14396 2746 14408
rect 2961 14399 3019 14405
rect 2961 14396 2973 14399
rect 2740 14368 2973 14396
rect 2740 14356 2746 14368
rect 2961 14365 2973 14368
rect 3007 14365 3019 14399
rect 4246 14396 4252 14408
rect 4207 14368 4252 14396
rect 2961 14359 3019 14365
rect 4246 14356 4252 14368
rect 4304 14356 4310 14408
rect 8588 14405 8616 14436
rect 11698 14424 11704 14476
rect 11756 14464 11762 14476
rect 11977 14467 12035 14473
rect 11977 14464 11989 14467
rect 11756 14436 11989 14464
rect 11756 14424 11762 14436
rect 11977 14433 11989 14436
rect 12023 14433 12035 14467
rect 11977 14427 12035 14433
rect 12526 14424 12532 14476
rect 12584 14464 12590 14476
rect 12986 14464 12992 14476
rect 12584 14436 12992 14464
rect 12584 14424 12590 14436
rect 12986 14424 12992 14436
rect 13044 14424 13050 14476
rect 15470 14424 15476 14476
rect 15528 14464 15534 14476
rect 16482 14464 16488 14476
rect 15528 14436 16488 14464
rect 15528 14424 15534 14436
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 16758 14473 16764 14476
rect 16752 14464 16764 14473
rect 16719 14436 16764 14464
rect 16752 14427 16764 14436
rect 16758 14424 16764 14427
rect 16816 14424 16822 14476
rect 20070 14464 20076 14476
rect 19720 14436 20076 14464
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14396 8631 14399
rect 8662 14396 8668 14408
rect 8619 14368 8668 14396
rect 8619 14365 8631 14368
rect 8573 14359 8631 14365
rect 8662 14356 8668 14368
rect 8720 14356 8726 14408
rect 9950 14356 9956 14408
rect 10008 14396 10014 14408
rect 10321 14399 10379 14405
rect 10321 14396 10333 14399
rect 10008 14368 10333 14396
rect 10008 14356 10014 14368
rect 10321 14365 10333 14368
rect 10367 14365 10379 14399
rect 10321 14359 10379 14365
rect 10505 14399 10563 14405
rect 10505 14365 10517 14399
rect 10551 14396 10563 14399
rect 10870 14396 10876 14408
rect 10551 14368 10876 14396
rect 10551 14365 10563 14368
rect 10505 14359 10563 14365
rect 2317 14331 2375 14337
rect 2317 14297 2329 14331
rect 2363 14328 2375 14331
rect 3602 14328 3608 14340
rect 2363 14300 3608 14328
rect 2363 14297 2375 14300
rect 2317 14291 2375 14297
rect 3602 14288 3608 14300
rect 3660 14288 3666 14340
rect 6914 14328 6920 14340
rect 6875 14300 6920 14328
rect 6914 14288 6920 14300
rect 6972 14288 6978 14340
rect 9493 14331 9551 14337
rect 9493 14297 9505 14331
rect 9539 14328 9551 14331
rect 10520 14328 10548 14359
rect 10870 14356 10876 14368
rect 10928 14356 10934 14408
rect 11238 14396 11244 14408
rect 11199 14368 11244 14396
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 15286 14396 15292 14408
rect 15247 14368 15292 14396
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 18598 14356 18604 14408
rect 18656 14396 18662 14408
rect 18966 14396 18972 14408
rect 18656 14368 18972 14396
rect 18656 14356 18662 14368
rect 18966 14356 18972 14368
rect 19024 14356 19030 14408
rect 19242 14356 19248 14408
rect 19300 14396 19306 14408
rect 19720 14405 19748 14436
rect 20070 14424 20076 14436
rect 20128 14424 20134 14476
rect 20714 14424 20720 14476
rect 20772 14464 20778 14476
rect 20901 14467 20959 14473
rect 20901 14464 20913 14467
rect 20772 14436 20913 14464
rect 20772 14424 20778 14436
rect 20901 14433 20913 14436
rect 20947 14433 20959 14467
rect 20901 14427 20959 14433
rect 21450 14424 21456 14476
rect 21508 14464 21514 14476
rect 22548 14467 22606 14473
rect 22548 14464 22560 14467
rect 21508 14436 22560 14464
rect 21508 14424 21514 14436
rect 22548 14433 22560 14436
rect 22594 14464 22606 14467
rect 23382 14464 23388 14476
rect 22594 14436 23388 14464
rect 22594 14433 22606 14436
rect 22548 14427 22606 14433
rect 23382 14424 23388 14436
rect 23440 14424 23446 14476
rect 25133 14467 25191 14473
rect 25133 14433 25145 14467
rect 25179 14464 25191 14467
rect 25498 14464 25504 14476
rect 25179 14436 25504 14464
rect 25179 14433 25191 14436
rect 25133 14427 25191 14433
rect 25498 14424 25504 14436
rect 25556 14424 25562 14476
rect 19705 14399 19763 14405
rect 19705 14396 19717 14399
rect 19300 14368 19717 14396
rect 19300 14356 19306 14368
rect 19705 14365 19717 14368
rect 19751 14365 19763 14399
rect 19705 14359 19763 14365
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14396 19947 14399
rect 20622 14396 20628 14408
rect 19935 14368 20628 14396
rect 19935 14365 19947 14368
rect 19889 14359 19947 14365
rect 19150 14328 19156 14340
rect 9539 14300 10548 14328
rect 19063 14300 19156 14328
rect 9539 14297 9551 14300
rect 9493 14291 9551 14297
rect 19150 14288 19156 14300
rect 19208 14328 19214 14340
rect 19904 14328 19932 14359
rect 20622 14356 20628 14368
rect 20680 14356 20686 14408
rect 22281 14399 22339 14405
rect 22281 14365 22293 14399
rect 22327 14365 22339 14399
rect 22281 14359 22339 14365
rect 19208 14300 19932 14328
rect 19208 14288 19214 14300
rect 20254 14288 20260 14340
rect 20312 14328 20318 14340
rect 20530 14328 20536 14340
rect 20312 14300 20536 14328
rect 20312 14288 20318 14300
rect 20530 14288 20536 14300
rect 20588 14288 20594 14340
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14260 1639 14263
rect 1762 14260 1768 14272
rect 1627 14232 1768 14260
rect 1627 14229 1639 14232
rect 1581 14223 1639 14229
rect 1762 14220 1768 14232
rect 1820 14220 1826 14272
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 5629 14263 5687 14269
rect 5629 14260 5641 14263
rect 5592 14232 5641 14260
rect 5592 14220 5598 14232
rect 5629 14229 5641 14232
rect 5675 14229 5687 14263
rect 6546 14260 6552 14272
rect 6507 14232 6552 14260
rect 5629 14223 5687 14229
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 9125 14263 9183 14269
rect 9125 14229 9137 14263
rect 9171 14260 9183 14263
rect 9582 14260 9588 14272
rect 9171 14232 9588 14260
rect 9171 14229 9183 14232
rect 9125 14223 9183 14229
rect 9582 14220 9588 14232
rect 9640 14220 9646 14272
rect 9861 14263 9919 14269
rect 9861 14229 9873 14263
rect 9907 14260 9919 14263
rect 10594 14260 10600 14272
rect 9907 14232 10600 14260
rect 9907 14229 9919 14232
rect 9861 14223 9919 14229
rect 10594 14220 10600 14232
rect 10652 14220 10658 14272
rect 12342 14220 12348 14272
rect 12400 14260 12406 14272
rect 14645 14263 14703 14269
rect 14645 14260 14657 14263
rect 12400 14232 14657 14260
rect 12400 14220 12406 14232
rect 14645 14229 14657 14232
rect 14691 14229 14703 14263
rect 20346 14260 20352 14272
rect 20307 14232 20352 14260
rect 14645 14223 14703 14229
rect 20346 14220 20352 14232
rect 20404 14220 20410 14272
rect 22296 14260 22324 14359
rect 24946 14356 24952 14408
rect 25004 14396 25010 14408
rect 25225 14399 25283 14405
rect 25225 14396 25237 14399
rect 25004 14368 25237 14396
rect 25004 14356 25010 14368
rect 25225 14365 25237 14368
rect 25271 14365 25283 14399
rect 25225 14359 25283 14365
rect 25317 14399 25375 14405
rect 25317 14365 25329 14399
rect 25363 14365 25375 14399
rect 26234 14396 26240 14408
rect 26195 14368 26240 14396
rect 25317 14359 25375 14365
rect 24026 14288 24032 14340
rect 24084 14328 24090 14340
rect 24581 14331 24639 14337
rect 24581 14328 24593 14331
rect 24084 14300 24593 14328
rect 24084 14288 24090 14300
rect 24581 14297 24593 14300
rect 24627 14297 24639 14331
rect 24581 14291 24639 14297
rect 25038 14288 25044 14340
rect 25096 14328 25102 14340
rect 25332 14328 25360 14359
rect 26234 14356 26240 14368
rect 26292 14356 26298 14408
rect 25096 14300 25360 14328
rect 25096 14288 25102 14300
rect 22646 14260 22652 14272
rect 22296 14232 22652 14260
rect 22646 14220 22652 14232
rect 22704 14220 22710 14272
rect 24118 14220 24124 14272
rect 24176 14260 24182 14272
rect 24213 14263 24271 14269
rect 24213 14260 24225 14263
rect 24176 14232 24225 14260
rect 24176 14220 24182 14232
rect 24213 14229 24225 14232
rect 24259 14229 24271 14263
rect 25774 14260 25780 14272
rect 25735 14232 25780 14260
rect 24213 14223 24271 14229
rect 25774 14220 25780 14232
rect 25832 14220 25838 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2038 14016 2044 14068
rect 2096 14056 2102 14068
rect 2409 14059 2467 14065
rect 2409 14056 2421 14059
rect 2096 14028 2421 14056
rect 2096 14016 2102 14028
rect 2409 14025 2421 14028
rect 2455 14025 2467 14059
rect 2682 14056 2688 14068
rect 2643 14028 2688 14056
rect 2409 14019 2467 14025
rect 2682 14016 2688 14028
rect 2740 14016 2746 14068
rect 2774 14016 2780 14068
rect 2832 14056 2838 14068
rect 3421 14059 3479 14065
rect 3421 14056 3433 14059
rect 2832 14028 3433 14056
rect 2832 14016 2838 14028
rect 3421 14025 3433 14028
rect 3467 14025 3479 14059
rect 8478 14056 8484 14068
rect 3421 14019 3479 14025
rect 6472 14028 8484 14056
rect 1946 13880 1952 13932
rect 2004 13880 2010 13932
rect 2038 13880 2044 13932
rect 2096 13920 2102 13932
rect 2225 13923 2283 13929
rect 2225 13920 2237 13923
rect 2096 13892 2237 13920
rect 2096 13880 2102 13892
rect 2225 13889 2237 13892
rect 2271 13920 2283 13923
rect 2700 13920 2728 14016
rect 3329 13991 3387 13997
rect 3329 13957 3341 13991
rect 3375 13988 3387 13991
rect 3602 13988 3608 14000
rect 3375 13960 3608 13988
rect 3375 13957 3387 13960
rect 3329 13951 3387 13957
rect 3602 13948 3608 13960
rect 3660 13948 3666 14000
rect 4982 13988 4988 14000
rect 3896 13960 4988 13988
rect 2271 13892 2728 13920
rect 2271 13889 2283 13892
rect 2225 13883 2283 13889
rect 1964 13852 1992 13880
rect 2682 13852 2688 13864
rect 1964 13824 2688 13852
rect 2682 13812 2688 13824
rect 2740 13812 2746 13864
rect 3620 13852 3648 13948
rect 3896 13929 3924 13960
rect 4982 13948 4988 13960
rect 5040 13948 5046 14000
rect 5166 13948 5172 14000
rect 5224 13988 5230 14000
rect 5224 13960 5672 13988
rect 5224 13948 5230 13960
rect 3881 13923 3939 13929
rect 3881 13889 3893 13923
rect 3927 13889 3939 13923
rect 3881 13883 3939 13889
rect 3973 13923 4031 13929
rect 3973 13889 3985 13923
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 4893 13923 4951 13929
rect 4893 13889 4905 13923
rect 4939 13920 4951 13923
rect 5442 13920 5448 13932
rect 4939 13892 5448 13920
rect 4939 13889 4951 13892
rect 4893 13883 4951 13889
rect 3988 13852 4016 13883
rect 5442 13880 5448 13892
rect 5500 13880 5506 13932
rect 5644 13929 5672 13960
rect 5629 13923 5687 13929
rect 5629 13889 5641 13923
rect 5675 13920 5687 13923
rect 5997 13923 6055 13929
rect 5997 13920 6009 13923
rect 5675 13892 6009 13920
rect 5675 13889 5687 13892
rect 5629 13883 5687 13889
rect 5997 13889 6009 13892
rect 6043 13889 6055 13923
rect 5997 13883 6055 13889
rect 3620 13824 4016 13852
rect 4525 13855 4583 13861
rect 4525 13821 4537 13855
rect 4571 13852 4583 13855
rect 5353 13855 5411 13861
rect 5353 13852 5365 13855
rect 4571 13824 5365 13852
rect 4571 13821 4583 13824
rect 4525 13815 4583 13821
rect 5353 13821 5365 13824
rect 5399 13852 5411 13855
rect 6472 13852 6500 14028
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 10870 14016 10876 14068
rect 10928 14056 10934 14068
rect 11241 14059 11299 14065
rect 11241 14056 11253 14059
rect 10928 14028 11253 14056
rect 10928 14016 10934 14028
rect 11241 14025 11253 14028
rect 11287 14056 11299 14059
rect 12250 14056 12256 14068
rect 11287 14028 12256 14056
rect 11287 14025 11299 14028
rect 11241 14019 11299 14025
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 12437 14059 12495 14065
rect 12437 14025 12449 14059
rect 12483 14056 12495 14059
rect 12526 14056 12532 14068
rect 12483 14028 12532 14056
rect 12483 14025 12495 14028
rect 12437 14019 12495 14025
rect 12526 14016 12532 14028
rect 12584 14016 12590 14068
rect 16482 14016 16488 14068
rect 16540 14056 16546 14068
rect 16945 14059 17003 14065
rect 16945 14056 16957 14059
rect 16540 14028 16957 14056
rect 16540 14016 16546 14028
rect 16945 14025 16957 14028
rect 16991 14025 17003 14059
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 16945 14019 17003 14025
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 17770 14056 17776 14068
rect 17731 14028 17776 14056
rect 17770 14016 17776 14028
rect 17828 14016 17834 14068
rect 18325 14059 18383 14065
rect 18325 14025 18337 14059
rect 18371 14056 18383 14059
rect 18506 14056 18512 14068
rect 18371 14028 18512 14056
rect 18371 14025 18383 14028
rect 18325 14019 18383 14025
rect 18506 14016 18512 14028
rect 18564 14016 18570 14068
rect 19061 14059 19119 14065
rect 19061 14025 19073 14059
rect 19107 14056 19119 14059
rect 19242 14056 19248 14068
rect 19107 14028 19248 14056
rect 19107 14025 19119 14028
rect 19061 14019 19119 14025
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 19337 14059 19395 14065
rect 19337 14025 19349 14059
rect 19383 14056 19395 14059
rect 19610 14056 19616 14068
rect 19383 14028 19616 14056
rect 19383 14025 19395 14028
rect 19337 14019 19395 14025
rect 19610 14016 19616 14028
rect 19668 14056 19674 14068
rect 20806 14056 20812 14068
rect 19668 14028 20668 14056
rect 20767 14028 20812 14056
rect 19668 14016 19674 14028
rect 8386 13988 8392 14000
rect 8347 13960 8392 13988
rect 8386 13948 8392 13960
rect 8444 13948 8450 14000
rect 11698 13948 11704 14000
rect 11756 13988 11762 14000
rect 11977 13991 12035 13997
rect 11977 13988 11989 13991
rect 11756 13960 11989 13988
rect 11756 13948 11762 13960
rect 11977 13957 11989 13960
rect 12023 13957 12035 13991
rect 13998 13988 14004 14000
rect 13959 13960 14004 13988
rect 11977 13951 12035 13957
rect 13998 13948 14004 13960
rect 14056 13948 14062 14000
rect 15286 13948 15292 14000
rect 15344 13988 15350 14000
rect 15933 13991 15991 13997
rect 15933 13988 15945 13991
rect 15344 13960 15945 13988
rect 15344 13948 15350 13960
rect 15933 13957 15945 13960
rect 15979 13957 15991 13991
rect 15933 13951 15991 13957
rect 6546 13880 6552 13932
rect 6604 13920 6610 13932
rect 6604 13892 7144 13920
rect 6604 13880 6610 13892
rect 7009 13855 7067 13861
rect 7009 13852 7021 13855
rect 5399 13824 6500 13852
rect 6564 13824 7021 13852
rect 5399 13821 5411 13824
rect 5353 13815 5411 13821
rect 1946 13784 1952 13796
rect 1859 13756 1952 13784
rect 1946 13744 1952 13756
rect 2004 13784 2010 13796
rect 2222 13784 2228 13796
rect 2004 13756 2228 13784
rect 2004 13744 2010 13756
rect 2222 13744 2228 13756
rect 2280 13744 2286 13796
rect 1581 13719 1639 13725
rect 1581 13685 1593 13719
rect 1627 13716 1639 13719
rect 1854 13716 1860 13728
rect 1627 13688 1860 13716
rect 1627 13685 1639 13688
rect 1581 13679 1639 13685
rect 1854 13676 1860 13688
rect 1912 13676 1918 13728
rect 2041 13719 2099 13725
rect 2041 13685 2053 13719
rect 2087 13716 2099 13719
rect 2409 13719 2467 13725
rect 2409 13716 2421 13719
rect 2087 13688 2421 13716
rect 2087 13685 2099 13688
rect 2041 13679 2099 13685
rect 2409 13685 2421 13688
rect 2455 13716 2467 13719
rect 3142 13716 3148 13728
rect 2455 13688 3148 13716
rect 2455 13685 2467 13688
rect 2409 13679 2467 13685
rect 3142 13676 3148 13688
rect 3200 13676 3206 13728
rect 3786 13716 3792 13728
rect 3747 13688 3792 13716
rect 3786 13676 3792 13688
rect 3844 13676 3850 13728
rect 6270 13676 6276 13728
rect 6328 13716 6334 13728
rect 6564 13725 6592 13824
rect 7009 13821 7021 13824
rect 7055 13821 7067 13855
rect 7116 13852 7144 13892
rect 7265 13855 7323 13861
rect 7265 13852 7277 13855
rect 7116 13824 7277 13852
rect 7009 13815 7067 13821
rect 7265 13821 7277 13824
rect 7311 13852 7323 13855
rect 7742 13852 7748 13864
rect 7311 13824 7748 13852
rect 7311 13821 7323 13824
rect 7265 13815 7323 13821
rect 7742 13812 7748 13824
rect 7800 13812 7806 13864
rect 9033 13855 9091 13861
rect 9033 13821 9045 13855
rect 9079 13852 9091 13855
rect 9122 13852 9128 13864
rect 9079 13824 9128 13852
rect 9079 13821 9091 13824
rect 9033 13815 9091 13821
rect 9122 13812 9128 13824
rect 9180 13812 9186 13864
rect 9582 13812 9588 13864
rect 9640 13852 9646 13864
rect 9769 13855 9827 13861
rect 9769 13852 9781 13855
rect 9640 13824 9781 13852
rect 9640 13812 9646 13824
rect 9769 13821 9781 13824
rect 9815 13852 9827 13855
rect 9861 13855 9919 13861
rect 9861 13852 9873 13855
rect 9815 13824 9873 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 9861 13821 9873 13824
rect 9907 13852 9919 13855
rect 11716 13852 11744 13948
rect 12158 13880 12164 13932
rect 12216 13920 12222 13932
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 12216 13892 13093 13920
rect 12216 13880 12222 13892
rect 13081 13889 13093 13892
rect 13127 13920 13139 13923
rect 13449 13923 13507 13929
rect 13449 13920 13461 13923
rect 13127 13892 13461 13920
rect 13127 13889 13139 13892
rect 13081 13883 13139 13889
rect 13449 13889 13461 13892
rect 13495 13889 13507 13923
rect 14016 13920 14044 13948
rect 14458 13920 14464 13932
rect 13449 13883 13507 13889
rect 13648 13892 14044 13920
rect 14419 13892 14464 13920
rect 12894 13852 12900 13864
rect 9907 13824 11744 13852
rect 12855 13824 12900 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 9401 13787 9459 13793
rect 9401 13753 9413 13787
rect 9447 13784 9459 13787
rect 9490 13784 9496 13796
rect 9447 13756 9496 13784
rect 9447 13753 9459 13756
rect 9401 13747 9459 13753
rect 9490 13744 9496 13756
rect 9548 13784 9554 13796
rect 10042 13784 10048 13796
rect 9548 13756 10048 13784
rect 9548 13744 9554 13756
rect 10042 13744 10048 13756
rect 10100 13793 10106 13796
rect 10100 13787 10164 13793
rect 10100 13753 10118 13787
rect 10152 13753 10164 13787
rect 10100 13747 10164 13753
rect 12805 13787 12863 13793
rect 12805 13753 12817 13787
rect 12851 13784 12863 13787
rect 13648 13784 13676 13892
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 14553 13923 14611 13929
rect 14553 13889 14565 13923
rect 14599 13889 14611 13923
rect 14553 13883 14611 13889
rect 15381 13923 15439 13929
rect 15381 13889 15393 13923
rect 15427 13920 15439 13923
rect 16577 13923 16635 13929
rect 16577 13920 16589 13923
rect 15427 13892 16589 13920
rect 15427 13889 15439 13892
rect 15381 13883 15439 13889
rect 16577 13889 16589 13892
rect 16623 13920 16635 13923
rect 16758 13920 16764 13932
rect 16623 13892 16764 13920
rect 16623 13889 16635 13892
rect 16577 13883 16635 13889
rect 13722 13812 13728 13864
rect 13780 13852 13786 13864
rect 13909 13855 13967 13861
rect 13909 13852 13921 13855
rect 13780 13824 13921 13852
rect 13780 13812 13786 13824
rect 13909 13821 13921 13824
rect 13955 13852 13967 13855
rect 14568 13852 14596 13883
rect 16758 13880 16764 13892
rect 16816 13920 16822 13932
rect 17420 13920 17448 14016
rect 18874 13948 18880 14000
rect 18932 13988 18938 14000
rect 19153 13991 19211 13997
rect 19153 13988 19165 13991
rect 18932 13960 19165 13988
rect 18932 13948 18938 13960
rect 19153 13957 19165 13960
rect 19199 13957 19211 13991
rect 20640 13988 20668 14028
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 21450 14056 21456 14068
rect 21411 14028 21456 14056
rect 21450 14016 21456 14028
rect 21508 14016 21514 14068
rect 21913 14059 21971 14065
rect 21913 14025 21925 14059
rect 21959 14056 21971 14059
rect 22002 14056 22008 14068
rect 21959 14028 22008 14056
rect 21959 14025 21971 14028
rect 21913 14019 21971 14025
rect 22002 14016 22008 14028
rect 22060 14016 22066 14068
rect 22738 14016 22744 14068
rect 22796 14056 22802 14068
rect 22925 14059 22983 14065
rect 22925 14056 22937 14059
rect 22796 14028 22937 14056
rect 22796 14016 22802 14028
rect 22925 14025 22937 14028
rect 22971 14025 22983 14059
rect 23474 14056 23480 14068
rect 23435 14028 23480 14056
rect 22925 14019 22983 14025
rect 23474 14016 23480 14028
rect 23532 14016 23538 14068
rect 23661 14059 23719 14065
rect 23661 14025 23673 14059
rect 23707 14056 23719 14059
rect 24026 14056 24032 14068
rect 23707 14028 24032 14056
rect 23707 14025 23719 14028
rect 23661 14019 23719 14025
rect 24026 14016 24032 14028
rect 24084 14016 24090 14068
rect 25406 14056 25412 14068
rect 25367 14028 25412 14056
rect 25406 14016 25412 14028
rect 25464 14016 25470 14068
rect 26237 14059 26295 14065
rect 26237 14025 26249 14059
rect 26283 14056 26295 14059
rect 26602 14056 26608 14068
rect 26283 14028 26608 14056
rect 26283 14025 26295 14028
rect 26237 14019 26295 14025
rect 26602 14016 26608 14028
rect 26660 14016 26666 14068
rect 22370 13988 22376 14000
rect 20640 13960 22376 13988
rect 19153 13951 19211 13957
rect 22370 13948 22376 13960
rect 22428 13948 22434 14000
rect 23492 13988 23520 14016
rect 24765 13991 24823 13997
rect 24765 13988 24777 13991
rect 23492 13960 24777 13988
rect 16816 13892 17448 13920
rect 16816 13880 16822 13892
rect 18046 13880 18052 13932
rect 18104 13920 18110 13932
rect 18104 13892 19564 13920
rect 18104 13880 18110 13892
rect 13955 13824 14596 13852
rect 13955 13821 13967 13824
rect 13909 13815 13967 13821
rect 15470 13812 15476 13864
rect 15528 13852 15534 13864
rect 15749 13855 15807 13861
rect 15749 13852 15761 13855
rect 15528 13824 15761 13852
rect 15528 13812 15534 13824
rect 15749 13821 15761 13824
rect 15795 13852 15807 13855
rect 16393 13855 16451 13861
rect 16393 13852 16405 13855
rect 15795 13824 16405 13852
rect 15795 13821 15807 13824
rect 15749 13815 15807 13821
rect 16393 13821 16405 13824
rect 16439 13821 16451 13855
rect 16393 13815 16451 13821
rect 19153 13855 19211 13861
rect 19153 13821 19165 13855
rect 19199 13821 19211 13855
rect 19153 13815 19211 13821
rect 19429 13855 19487 13861
rect 19429 13821 19441 13855
rect 19475 13821 19487 13855
rect 19536 13852 19564 13892
rect 20622 13880 20628 13932
rect 20680 13920 20686 13932
rect 20680 13892 21956 13920
rect 20680 13880 20686 13892
rect 20438 13852 20444 13864
rect 19536 13824 20444 13852
rect 19429 13815 19487 13821
rect 12851 13756 13676 13784
rect 12851 13753 12863 13756
rect 12805 13747 12863 13753
rect 10100 13744 10106 13747
rect 14090 13744 14096 13796
rect 14148 13784 14154 13796
rect 14369 13787 14427 13793
rect 14369 13784 14381 13787
rect 14148 13756 14381 13784
rect 14148 13744 14154 13756
rect 14369 13753 14381 13756
rect 14415 13784 14427 13787
rect 17954 13784 17960 13796
rect 14415 13756 17960 13784
rect 14415 13753 14427 13756
rect 14369 13747 14427 13753
rect 17954 13744 17960 13756
rect 18012 13744 18018 13796
rect 18506 13744 18512 13796
rect 18564 13784 18570 13796
rect 18877 13787 18935 13793
rect 18877 13784 18889 13787
rect 18564 13756 18889 13784
rect 18564 13744 18570 13756
rect 18877 13753 18889 13756
rect 18923 13784 18935 13787
rect 19061 13787 19119 13793
rect 19061 13784 19073 13787
rect 18923 13756 19073 13784
rect 18923 13753 18935 13756
rect 18877 13747 18935 13753
rect 19061 13753 19073 13756
rect 19107 13753 19119 13787
rect 19168 13784 19196 13815
rect 19444 13784 19472 13815
rect 20438 13812 20444 13824
rect 20496 13812 20502 13864
rect 21358 13812 21364 13864
rect 21416 13852 21422 13864
rect 21729 13855 21787 13861
rect 21729 13852 21741 13855
rect 21416 13824 21741 13852
rect 21416 13812 21422 13824
rect 21729 13821 21741 13824
rect 21775 13852 21787 13855
rect 21928 13852 21956 13892
rect 22002 13880 22008 13932
rect 22060 13920 22066 13932
rect 22465 13923 22523 13929
rect 22465 13920 22477 13923
rect 22060 13892 22477 13920
rect 22060 13880 22066 13892
rect 22465 13889 22477 13892
rect 22511 13889 22523 13923
rect 24118 13920 24124 13932
rect 24079 13892 24124 13920
rect 22465 13883 22523 13889
rect 24118 13880 24124 13892
rect 24176 13880 24182 13932
rect 24228 13929 24256 13960
rect 24765 13957 24777 13960
rect 24811 13988 24823 13991
rect 25038 13988 25044 14000
rect 24811 13960 25044 13988
rect 24811 13957 24823 13960
rect 24765 13951 24823 13957
rect 25038 13948 25044 13960
rect 25096 13948 25102 14000
rect 25222 13948 25228 14000
rect 25280 13948 25286 14000
rect 24213 13923 24271 13929
rect 24213 13889 24225 13923
rect 24259 13889 24271 13923
rect 24213 13883 24271 13889
rect 24302 13880 24308 13932
rect 24360 13920 24366 13932
rect 25240 13920 25268 13948
rect 24360 13892 25268 13920
rect 24360 13880 24366 13892
rect 25406 13880 25412 13932
rect 25464 13920 25470 13932
rect 25866 13920 25872 13932
rect 25464 13892 25872 13920
rect 25464 13880 25470 13892
rect 25866 13880 25872 13892
rect 25924 13880 25930 13932
rect 25222 13852 25228 13864
rect 21775 13824 21864 13852
rect 21928 13824 22692 13852
rect 25183 13824 25228 13852
rect 21775 13821 21787 13824
rect 21729 13815 21787 13821
rect 19168 13756 19472 13784
rect 19696 13787 19754 13793
rect 19061 13747 19119 13753
rect 19696 13753 19708 13787
rect 19742 13784 19754 13787
rect 20346 13784 20352 13796
rect 19742 13756 20352 13784
rect 19742 13753 19754 13756
rect 19696 13747 19754 13753
rect 20346 13744 20352 13756
rect 20404 13744 20410 13796
rect 6549 13719 6607 13725
rect 6549 13716 6561 13719
rect 6328 13688 6561 13716
rect 6328 13676 6334 13688
rect 6549 13685 6561 13688
rect 6595 13685 6607 13719
rect 6549 13679 6607 13685
rect 10686 13676 10692 13728
rect 10744 13716 10750 13728
rect 10962 13716 10968 13728
rect 10744 13688 10968 13716
rect 10744 13676 10750 13688
rect 10962 13676 10968 13688
rect 11020 13676 11026 13728
rect 11054 13676 11060 13728
rect 11112 13716 11118 13728
rect 12894 13716 12900 13728
rect 11112 13688 12900 13716
rect 11112 13676 11118 13688
rect 12894 13676 12900 13688
rect 12952 13716 12958 13728
rect 15013 13719 15071 13725
rect 15013 13716 15025 13719
rect 12952 13688 15025 13716
rect 12952 13676 12958 13688
rect 15013 13685 15025 13688
rect 15059 13685 15071 13719
rect 15013 13679 15071 13685
rect 15930 13676 15936 13728
rect 15988 13716 15994 13728
rect 16301 13719 16359 13725
rect 16301 13716 16313 13719
rect 15988 13688 16313 13716
rect 15988 13676 15994 13688
rect 16301 13685 16313 13688
rect 16347 13685 16359 13719
rect 16301 13679 16359 13685
rect 18417 13719 18475 13725
rect 18417 13685 18429 13719
rect 18463 13716 18475 13719
rect 18782 13716 18788 13728
rect 18463 13688 18788 13716
rect 18463 13685 18475 13688
rect 18417 13679 18475 13685
rect 18782 13676 18788 13688
rect 18840 13676 18846 13728
rect 19150 13676 19156 13728
rect 19208 13716 19214 13728
rect 20070 13716 20076 13728
rect 19208 13688 20076 13716
rect 19208 13676 19214 13688
rect 20070 13676 20076 13688
rect 20128 13676 20134 13728
rect 21836 13716 21864 13824
rect 22094 13744 22100 13796
rect 22152 13784 22158 13796
rect 22281 13787 22339 13793
rect 22281 13784 22293 13787
rect 22152 13756 22293 13784
rect 22152 13744 22158 13756
rect 22281 13753 22293 13756
rect 22327 13753 22339 13787
rect 22664 13784 22692 13824
rect 25222 13812 25228 13824
rect 25280 13852 25286 13864
rect 25777 13855 25835 13861
rect 25777 13852 25789 13855
rect 25280 13824 25789 13852
rect 25280 13812 25286 13824
rect 25777 13821 25789 13824
rect 25823 13821 25835 13855
rect 25777 13815 25835 13821
rect 25866 13784 25872 13796
rect 22664 13756 25872 13784
rect 22281 13747 22339 13753
rect 25866 13744 25872 13756
rect 25924 13744 25930 13796
rect 22373 13719 22431 13725
rect 22373 13716 22385 13719
rect 21836 13688 22385 13716
rect 22373 13685 22385 13688
rect 22419 13716 22431 13719
rect 22646 13716 22652 13728
rect 22419 13688 22652 13716
rect 22419 13685 22431 13688
rect 22373 13679 22431 13685
rect 22646 13676 22652 13688
rect 22704 13676 22710 13728
rect 24026 13716 24032 13728
rect 23987 13688 24032 13716
rect 24026 13676 24032 13688
rect 24084 13676 24090 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1854 13472 1860 13524
rect 1912 13512 1918 13524
rect 2222 13512 2228 13524
rect 1912 13484 2228 13512
rect 1912 13472 1918 13484
rect 2222 13472 2228 13484
rect 2280 13472 2286 13524
rect 2317 13515 2375 13521
rect 2317 13481 2329 13515
rect 2363 13512 2375 13515
rect 2406 13512 2412 13524
rect 2363 13484 2412 13512
rect 2363 13481 2375 13484
rect 2317 13475 2375 13481
rect 2406 13472 2412 13484
rect 2464 13472 2470 13524
rect 3142 13472 3148 13524
rect 3200 13512 3206 13524
rect 3605 13515 3663 13521
rect 3605 13512 3617 13515
rect 3200 13484 3617 13512
rect 3200 13472 3206 13484
rect 3605 13481 3617 13484
rect 3651 13481 3663 13515
rect 4798 13512 4804 13524
rect 4759 13484 4804 13512
rect 3605 13475 3663 13481
rect 4798 13472 4804 13484
rect 4856 13472 4862 13524
rect 5166 13472 5172 13524
rect 5224 13512 5230 13524
rect 5261 13515 5319 13521
rect 5261 13512 5273 13515
rect 5224 13484 5273 13512
rect 5224 13472 5230 13484
rect 5261 13481 5273 13484
rect 5307 13481 5319 13515
rect 7742 13512 7748 13524
rect 7703 13484 7748 13512
rect 5261 13475 5319 13481
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 8110 13472 8116 13524
rect 8168 13512 8174 13524
rect 8294 13512 8300 13524
rect 8168 13484 8300 13512
rect 8168 13472 8174 13484
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 8662 13512 8668 13524
rect 8623 13484 8668 13512
rect 8662 13472 8668 13484
rect 8720 13472 8726 13524
rect 9030 13512 9036 13524
rect 8991 13484 9036 13512
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 9490 13512 9496 13524
rect 9451 13484 9496 13512
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13512 9735 13515
rect 10134 13512 10140 13524
rect 9723 13484 10140 13512
rect 9723 13481 9735 13484
rect 9677 13475 9735 13481
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 11238 13512 11244 13524
rect 11199 13484 11244 13512
rect 11238 13472 11244 13484
rect 11296 13472 11302 13524
rect 11606 13512 11612 13524
rect 11567 13484 11612 13512
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 12713 13515 12771 13521
rect 12713 13481 12725 13515
rect 12759 13512 12771 13515
rect 13170 13512 13176 13524
rect 12759 13484 13176 13512
rect 12759 13481 12771 13484
rect 12713 13475 12771 13481
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 13906 13512 13912 13524
rect 13867 13484 13912 13512
rect 13906 13472 13912 13484
rect 13964 13472 13970 13524
rect 14182 13512 14188 13524
rect 14143 13484 14188 13512
rect 14182 13472 14188 13484
rect 14240 13472 14246 13524
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 17037 13515 17095 13521
rect 17037 13512 17049 13515
rect 16632 13484 17049 13512
rect 16632 13472 16638 13484
rect 17037 13481 17049 13484
rect 17083 13512 17095 13515
rect 17862 13512 17868 13524
rect 17083 13484 17868 13512
rect 17083 13481 17095 13484
rect 17037 13475 17095 13481
rect 17862 13472 17868 13484
rect 17920 13472 17926 13524
rect 19058 13512 19064 13524
rect 19019 13484 19064 13512
rect 19058 13472 19064 13484
rect 19116 13472 19122 13524
rect 19242 13472 19248 13524
rect 19300 13512 19306 13524
rect 19521 13515 19579 13521
rect 19521 13512 19533 13515
rect 19300 13484 19533 13512
rect 19300 13472 19306 13484
rect 19521 13481 19533 13484
rect 19567 13512 19579 13515
rect 21818 13512 21824 13524
rect 19567 13484 21824 13512
rect 19567 13481 19579 13484
rect 19521 13475 19579 13481
rect 21818 13472 21824 13484
rect 21876 13472 21882 13524
rect 22002 13472 22008 13524
rect 22060 13512 22066 13524
rect 22833 13515 22891 13521
rect 22833 13512 22845 13515
rect 22060 13484 22845 13512
rect 22060 13472 22066 13484
rect 22833 13481 22845 13484
rect 22879 13481 22891 13515
rect 22833 13475 22891 13481
rect 23293 13515 23351 13521
rect 23293 13481 23305 13515
rect 23339 13512 23351 13515
rect 23385 13515 23443 13521
rect 23385 13512 23397 13515
rect 23339 13484 23397 13512
rect 23339 13481 23351 13484
rect 23293 13475 23351 13481
rect 23385 13481 23397 13484
rect 23431 13512 23443 13515
rect 24026 13512 24032 13524
rect 23431 13484 24032 13512
rect 23431 13481 23443 13484
rect 23385 13475 23443 13481
rect 24026 13472 24032 13484
rect 24084 13472 24090 13524
rect 24489 13515 24547 13521
rect 24489 13481 24501 13515
rect 24535 13512 24547 13515
rect 24578 13512 24584 13524
rect 24535 13484 24584 13512
rect 24535 13481 24547 13484
rect 24489 13475 24547 13481
rect 1673 13447 1731 13453
rect 1673 13413 1685 13447
rect 1719 13444 1731 13447
rect 2038 13444 2044 13456
rect 1719 13416 2044 13444
rect 1719 13413 1731 13416
rect 1673 13407 1731 13413
rect 2038 13404 2044 13416
rect 2096 13404 2102 13456
rect 2958 13404 2964 13456
rect 3016 13444 3022 13456
rect 3237 13447 3295 13453
rect 3237 13444 3249 13447
rect 3016 13416 3249 13444
rect 3016 13404 3022 13416
rect 3237 13413 3249 13416
rect 3283 13413 3295 13447
rect 4338 13444 4344 13456
rect 4251 13416 4344 13444
rect 3237 13407 3295 13413
rect 4338 13404 4344 13416
rect 4396 13444 4402 13456
rect 6270 13444 6276 13456
rect 4396 13416 6276 13444
rect 4396 13404 4402 13416
rect 6270 13404 6276 13416
rect 6328 13404 6334 13456
rect 11149 13447 11207 13453
rect 11149 13413 11161 13447
rect 11195 13444 11207 13447
rect 11514 13444 11520 13456
rect 11195 13416 11520 13444
rect 11195 13413 11207 13416
rect 11149 13407 11207 13413
rect 11514 13404 11520 13416
rect 11572 13404 11578 13456
rect 13814 13404 13820 13456
rect 13872 13444 13878 13456
rect 17310 13444 17316 13456
rect 13872 13416 16620 13444
rect 17271 13416 17316 13444
rect 13872 13404 13878 13416
rect 2682 13336 2688 13388
rect 2740 13376 2746 13388
rect 2869 13379 2927 13385
rect 2869 13376 2881 13379
rect 2740 13348 2881 13376
rect 2740 13336 2746 13348
rect 2869 13345 2881 13348
rect 2915 13345 2927 13379
rect 2869 13339 2927 13345
rect 5169 13379 5227 13385
rect 5169 13345 5181 13379
rect 5215 13376 5227 13379
rect 5442 13376 5448 13388
rect 5215 13348 5448 13376
rect 5215 13345 5227 13348
rect 5169 13339 5227 13345
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 6178 13336 6184 13388
rect 6236 13376 6242 13388
rect 6621 13379 6679 13385
rect 6621 13376 6633 13379
rect 6236 13348 6633 13376
rect 6236 13336 6242 13348
rect 6621 13345 6633 13348
rect 6667 13345 6679 13379
rect 6621 13339 6679 13345
rect 7190 13336 7196 13388
rect 7248 13376 7254 13388
rect 9306 13376 9312 13388
rect 7248 13348 9312 13376
rect 7248 13336 7254 13348
rect 9306 13336 9312 13348
rect 9364 13376 9370 13388
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 9364 13348 10057 13376
rect 9364 13336 9370 13348
rect 10045 13345 10057 13348
rect 10091 13376 10103 13379
rect 10870 13376 10876 13388
rect 10091 13348 10876 13376
rect 10091 13345 10103 13348
rect 10045 13339 10103 13345
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 11701 13379 11759 13385
rect 11701 13345 11713 13379
rect 11747 13376 11759 13379
rect 11882 13376 11888 13388
rect 11747 13348 11888 13376
rect 11747 13345 11759 13348
rect 11701 13339 11759 13345
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 14090 13336 14096 13388
rect 14148 13376 14154 13388
rect 14734 13376 14740 13388
rect 14148 13348 14740 13376
rect 14148 13336 14154 13348
rect 14734 13336 14740 13348
rect 14792 13336 14798 13388
rect 16298 13376 16304 13388
rect 16259 13348 16304 13376
rect 16298 13336 16304 13348
rect 16356 13336 16362 13388
rect 16592 13376 16620 13416
rect 17310 13404 17316 13416
rect 17368 13404 17374 13456
rect 18874 13404 18880 13456
rect 18932 13444 18938 13456
rect 19794 13444 19800 13456
rect 18932 13416 19800 13444
rect 18932 13404 18938 13416
rect 19794 13404 19800 13416
rect 19852 13444 19858 13456
rect 20073 13447 20131 13453
rect 20073 13444 20085 13447
rect 19852 13416 20085 13444
rect 19852 13404 19858 13416
rect 20073 13413 20085 13416
rect 20119 13444 20131 13447
rect 22646 13444 22652 13456
rect 20119 13416 22652 13444
rect 20119 13413 20131 13416
rect 20073 13407 20131 13413
rect 17862 13376 17868 13388
rect 16592 13348 17868 13376
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 18414 13336 18420 13388
rect 18472 13376 18478 13388
rect 19426 13376 19432 13388
rect 18472 13348 19432 13376
rect 18472 13336 18478 13348
rect 19426 13336 19432 13348
rect 19484 13336 19490 13388
rect 20622 13336 20628 13388
rect 20680 13336 20686 13388
rect 1854 13268 1860 13320
rect 1912 13308 1918 13320
rect 2130 13308 2136 13320
rect 1912 13280 2136 13308
rect 1912 13268 1918 13280
rect 2130 13268 2136 13280
rect 2188 13308 2194 13320
rect 2409 13311 2467 13317
rect 2409 13308 2421 13311
rect 2188 13280 2421 13308
rect 2188 13268 2194 13280
rect 2409 13277 2421 13280
rect 2455 13277 2467 13311
rect 2409 13271 2467 13277
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 4982 13308 4988 13320
rect 4120 13280 4988 13308
rect 4120 13268 4126 13280
rect 4982 13268 4988 13280
rect 5040 13268 5046 13320
rect 5350 13308 5356 13320
rect 5311 13280 5356 13308
rect 5350 13268 5356 13280
rect 5408 13268 5414 13320
rect 6270 13268 6276 13320
rect 6328 13308 6334 13320
rect 6365 13311 6423 13317
rect 6365 13308 6377 13311
rect 6328 13280 6377 13308
rect 6328 13268 6334 13280
rect 6365 13277 6377 13280
rect 6411 13277 6423 13311
rect 6365 13271 6423 13277
rect 9490 13268 9496 13320
rect 9548 13308 9554 13320
rect 10137 13311 10195 13317
rect 10137 13308 10149 13311
rect 9548 13280 10149 13308
rect 9548 13268 9554 13280
rect 10137 13277 10149 13280
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13308 10287 13311
rect 10594 13308 10600 13320
rect 10275 13280 10600 13308
rect 10275 13277 10287 13280
rect 10229 13271 10287 13277
rect 4154 13200 4160 13252
rect 4212 13240 4218 13252
rect 4617 13243 4675 13249
rect 4617 13240 4629 13243
rect 4212 13212 4629 13240
rect 4212 13200 4218 13212
rect 4617 13209 4629 13212
rect 4663 13209 4675 13243
rect 4617 13203 4675 13209
rect 5074 13200 5080 13252
rect 5132 13240 5138 13252
rect 5132 13212 6408 13240
rect 5132 13200 5138 13212
rect 1670 13132 1676 13184
rect 1728 13172 1734 13184
rect 1857 13175 1915 13181
rect 1857 13172 1869 13175
rect 1728 13144 1869 13172
rect 1728 13132 1734 13144
rect 1857 13141 1869 13144
rect 1903 13141 1915 13175
rect 1857 13135 1915 13141
rect 5905 13175 5963 13181
rect 5905 13141 5917 13175
rect 5951 13172 5963 13175
rect 5994 13172 6000 13184
rect 5951 13144 6000 13172
rect 5951 13141 5963 13144
rect 5905 13135 5963 13141
rect 5994 13132 6000 13144
rect 6052 13132 6058 13184
rect 6178 13172 6184 13184
rect 6139 13144 6184 13172
rect 6178 13132 6184 13144
rect 6236 13132 6242 13184
rect 6380 13172 6408 13212
rect 10042 13200 10048 13252
rect 10100 13240 10106 13252
rect 10244 13240 10272 13271
rect 10594 13268 10600 13280
rect 10652 13308 10658 13320
rect 10689 13311 10747 13317
rect 10689 13308 10701 13311
rect 10652 13280 10701 13308
rect 10652 13268 10658 13280
rect 10689 13277 10701 13280
rect 10735 13308 10747 13311
rect 11422 13308 11428 13320
rect 10735 13280 11428 13308
rect 10735 13277 10747 13280
rect 10689 13271 10747 13277
rect 11422 13268 11428 13280
rect 11480 13308 11486 13320
rect 11793 13311 11851 13317
rect 11793 13308 11805 13311
rect 11480 13280 11805 13308
rect 11480 13268 11486 13280
rect 11793 13277 11805 13280
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 10100 13212 10272 13240
rect 11808 13240 11836 13271
rect 12250 13268 12256 13320
rect 12308 13308 12314 13320
rect 12345 13311 12403 13317
rect 12345 13308 12357 13311
rect 12308 13280 12357 13308
rect 12308 13268 12314 13280
rect 12345 13277 12357 13280
rect 12391 13308 12403 13311
rect 13262 13308 13268 13320
rect 12391 13280 13124 13308
rect 13223 13280 13268 13308
rect 12391 13277 12403 13280
rect 12345 13271 12403 13277
rect 13096 13240 13124 13280
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 13449 13311 13507 13317
rect 13449 13277 13461 13311
rect 13495 13308 13507 13311
rect 13722 13308 13728 13320
rect 13495 13280 13728 13308
rect 13495 13277 13507 13280
rect 13449 13271 13507 13277
rect 13464 13240 13492 13271
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 14918 13308 14924 13320
rect 14879 13280 14924 13308
rect 14918 13268 14924 13280
rect 14976 13268 14982 13320
rect 15286 13268 15292 13320
rect 15344 13308 15350 13320
rect 16393 13311 16451 13317
rect 16393 13308 16405 13311
rect 15344 13280 16405 13308
rect 15344 13268 15350 13280
rect 16393 13277 16405 13280
rect 16439 13277 16451 13311
rect 16393 13271 16451 13277
rect 16485 13311 16543 13317
rect 16485 13277 16497 13311
rect 16531 13277 16543 13311
rect 16485 13271 16543 13277
rect 16500 13240 16528 13271
rect 17586 13268 17592 13320
rect 17644 13308 17650 13320
rect 17957 13311 18015 13317
rect 17957 13308 17969 13311
rect 17644 13280 17969 13308
rect 17644 13268 17650 13280
rect 17957 13277 17969 13280
rect 18003 13277 18015 13311
rect 17957 13271 18015 13277
rect 18141 13311 18199 13317
rect 18141 13277 18153 13311
rect 18187 13308 18199 13311
rect 18969 13311 19027 13317
rect 18187 13280 18644 13308
rect 18187 13277 18199 13280
rect 18141 13271 18199 13277
rect 16758 13240 16764 13252
rect 11808 13212 13032 13240
rect 13096 13212 13492 13240
rect 15764 13212 16764 13240
rect 10100 13200 10106 13212
rect 7282 13172 7288 13184
rect 6380 13144 7288 13172
rect 7282 13132 7288 13144
rect 7340 13172 7346 13184
rect 11146 13172 11152 13184
rect 7340 13144 11152 13172
rect 7340 13132 7346 13144
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 12802 13172 12808 13184
rect 12763 13144 12808 13172
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 13004 13172 13032 13212
rect 15764 13184 15792 13212
rect 16758 13200 16764 13212
rect 16816 13200 16822 13252
rect 17494 13240 17500 13252
rect 17455 13212 17500 13240
rect 17494 13200 17500 13212
rect 17552 13200 17558 13252
rect 18616 13249 18644 13280
rect 18969 13277 18981 13311
rect 19015 13308 19027 13311
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19015 13280 19717 13308
rect 19015 13277 19027 13280
rect 18969 13271 19027 13277
rect 19705 13277 19717 13280
rect 19751 13308 19763 13311
rect 20640 13308 20668 13336
rect 20916 13317 20944 13416
rect 22646 13404 22652 13416
rect 22704 13404 22710 13456
rect 21168 13379 21226 13385
rect 21168 13345 21180 13379
rect 21214 13376 21226 13379
rect 21450 13376 21456 13388
rect 21214 13348 21456 13376
rect 21214 13345 21226 13348
rect 21168 13339 21226 13345
rect 21450 13336 21456 13348
rect 21508 13336 21514 13388
rect 22738 13336 22744 13388
rect 22796 13376 22802 13388
rect 23753 13379 23811 13385
rect 23753 13376 23765 13379
rect 22796 13348 23765 13376
rect 22796 13336 22802 13348
rect 23753 13345 23765 13348
rect 23799 13345 23811 13379
rect 23753 13339 23811 13345
rect 23845 13379 23903 13385
rect 23845 13345 23857 13379
rect 23891 13376 23903 13379
rect 24302 13376 24308 13388
rect 23891 13348 24308 13376
rect 23891 13345 23903 13348
rect 23845 13339 23903 13345
rect 19751 13280 20668 13308
rect 20901 13311 20959 13317
rect 19751 13277 19763 13280
rect 19705 13271 19763 13277
rect 20901 13277 20913 13311
rect 20947 13277 20959 13311
rect 20901 13271 20959 13277
rect 22278 13268 22284 13320
rect 22336 13308 22342 13320
rect 22554 13308 22560 13320
rect 22336 13280 22560 13308
rect 22336 13268 22342 13280
rect 22554 13268 22560 13280
rect 22612 13268 22618 13320
rect 23382 13268 23388 13320
rect 23440 13308 23446 13320
rect 23860 13308 23888 13339
rect 24302 13336 24308 13348
rect 24360 13336 24366 13388
rect 23440 13280 23888 13308
rect 24029 13311 24087 13317
rect 23440 13268 23446 13280
rect 24029 13277 24041 13311
rect 24075 13308 24087 13311
rect 24504 13308 24532 13475
rect 24578 13472 24584 13484
rect 24636 13472 24642 13524
rect 24854 13472 24860 13524
rect 24912 13512 24918 13524
rect 25133 13515 25191 13521
rect 24912 13484 24992 13512
rect 24912 13472 24918 13484
rect 24964 13444 24992 13484
rect 25133 13481 25145 13515
rect 25179 13512 25191 13515
rect 25314 13512 25320 13524
rect 25179 13484 25320 13512
rect 25179 13481 25191 13484
rect 25133 13475 25191 13481
rect 25314 13472 25320 13484
rect 25372 13472 25378 13524
rect 25866 13512 25872 13524
rect 25827 13484 25872 13512
rect 25866 13472 25872 13484
rect 25924 13472 25930 13524
rect 26234 13512 26240 13524
rect 26195 13484 26240 13512
rect 26234 13472 26240 13484
rect 26292 13472 26298 13524
rect 24964 13416 25360 13444
rect 24854 13336 24860 13388
rect 24912 13376 24918 13388
rect 24949 13379 25007 13385
rect 24949 13376 24961 13379
rect 24912 13348 24961 13376
rect 24912 13336 24918 13348
rect 24949 13345 24961 13348
rect 24995 13376 25007 13379
rect 25038 13376 25044 13388
rect 24995 13348 25044 13376
rect 24995 13345 25007 13348
rect 24949 13339 25007 13345
rect 25038 13336 25044 13348
rect 25096 13336 25102 13388
rect 25332 13320 25360 13416
rect 24075 13280 24532 13308
rect 24075 13277 24087 13280
rect 24029 13271 24087 13277
rect 18601 13243 18659 13249
rect 18601 13209 18613 13243
rect 18647 13240 18659 13243
rect 19150 13240 19156 13252
rect 18647 13212 19156 13240
rect 18647 13209 18659 13212
rect 18601 13203 18659 13209
rect 19150 13200 19156 13212
rect 19208 13200 19214 13252
rect 23474 13200 23480 13252
rect 23532 13240 23538 13252
rect 24044 13240 24072 13271
rect 25314 13268 25320 13320
rect 25372 13268 25378 13320
rect 23532 13212 24072 13240
rect 23532 13200 23538 13212
rect 13906 13172 13912 13184
rect 13004 13144 13912 13172
rect 13906 13132 13912 13144
rect 13964 13132 13970 13184
rect 14642 13172 14648 13184
rect 14603 13144 14648 13172
rect 14642 13132 14648 13144
rect 14700 13132 14706 13184
rect 15746 13172 15752 13184
rect 15707 13144 15752 13172
rect 15746 13132 15752 13144
rect 15804 13132 15810 13184
rect 15930 13172 15936 13184
rect 15891 13144 15936 13172
rect 15930 13132 15936 13144
rect 15988 13132 15994 13184
rect 20717 13175 20775 13181
rect 20717 13141 20729 13175
rect 20763 13172 20775 13175
rect 20806 13172 20812 13184
rect 20763 13144 20812 13172
rect 20763 13141 20775 13144
rect 20717 13135 20775 13141
rect 20806 13132 20812 13144
rect 20864 13132 20870 13184
rect 22278 13172 22284 13184
rect 22239 13144 22284 13172
rect 22278 13132 22284 13144
rect 22336 13132 22342 13184
rect 23842 13132 23848 13184
rect 23900 13172 23906 13184
rect 24026 13172 24032 13184
rect 23900 13144 24032 13172
rect 23900 13132 23906 13144
rect 24026 13132 24032 13144
rect 24084 13132 24090 13184
rect 24857 13175 24915 13181
rect 24857 13141 24869 13175
rect 24903 13172 24915 13175
rect 24946 13172 24952 13184
rect 24903 13144 24952 13172
rect 24903 13141 24915 13144
rect 24857 13135 24915 13141
rect 24946 13132 24952 13144
rect 25004 13132 25010 13184
rect 25498 13172 25504 13184
rect 25459 13144 25504 13172
rect 25498 13132 25504 13144
rect 25556 13132 25562 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1854 12968 1860 12980
rect 1815 12940 1860 12968
rect 1854 12928 1860 12940
rect 1912 12928 1918 12980
rect 2038 12968 2044 12980
rect 1999 12940 2044 12968
rect 2038 12928 2044 12940
rect 2096 12928 2102 12980
rect 2774 12928 2780 12980
rect 2832 12968 2838 12980
rect 3053 12971 3111 12977
rect 3053 12968 3065 12971
rect 2832 12940 3065 12968
rect 2832 12928 2838 12940
rect 3053 12937 3065 12940
rect 3099 12937 3111 12971
rect 3053 12931 3111 12937
rect 4709 12971 4767 12977
rect 4709 12937 4721 12971
rect 4755 12968 4767 12971
rect 5350 12968 5356 12980
rect 4755 12940 5356 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 8938 12928 8944 12980
rect 8996 12968 9002 12980
rect 9490 12968 9496 12980
rect 8996 12940 9496 12968
rect 8996 12928 9002 12940
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 9953 12971 10011 12977
rect 9953 12937 9965 12971
rect 9999 12968 10011 12971
rect 10226 12968 10232 12980
rect 9999 12940 10232 12968
rect 9999 12937 10011 12940
rect 9953 12931 10011 12937
rect 10226 12928 10232 12940
rect 10284 12928 10290 12980
rect 10686 12928 10692 12980
rect 10744 12968 10750 12980
rect 11238 12968 11244 12980
rect 10744 12940 11244 12968
rect 10744 12928 10750 12940
rect 11238 12928 11244 12940
rect 11296 12928 11302 12980
rect 11606 12968 11612 12980
rect 11567 12940 11612 12968
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 12526 12928 12532 12980
rect 12584 12968 12590 12980
rect 12897 12971 12955 12977
rect 12897 12968 12909 12971
rect 12584 12940 12909 12968
rect 12584 12928 12590 12940
rect 12897 12937 12909 12940
rect 12943 12968 12955 12971
rect 13262 12968 13268 12980
rect 12943 12940 13268 12968
rect 12943 12937 12955 12940
rect 12897 12931 12955 12937
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 14366 12968 14372 12980
rect 14327 12940 14372 12968
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 16114 12968 16120 12980
rect 16075 12940 16120 12968
rect 16114 12928 16120 12940
rect 16172 12968 16178 12980
rect 16482 12968 16488 12980
rect 16172 12940 16488 12968
rect 16172 12928 16178 12940
rect 16482 12928 16488 12940
rect 16540 12968 16546 12980
rect 18414 12968 18420 12980
rect 16540 12940 16712 12968
rect 18375 12940 18420 12968
rect 16540 12928 16546 12940
rect 2130 12860 2136 12912
rect 2188 12900 2194 12912
rect 3421 12903 3479 12909
rect 3421 12900 3433 12903
rect 2188 12872 3433 12900
rect 2188 12860 2194 12872
rect 2608 12841 2636 12872
rect 3421 12869 3433 12872
rect 3467 12869 3479 12903
rect 3421 12863 3479 12869
rect 3605 12903 3663 12909
rect 3605 12869 3617 12903
rect 3651 12900 3663 12903
rect 5442 12900 5448 12912
rect 3651 12872 5448 12900
rect 3651 12869 3663 12872
rect 3605 12863 3663 12869
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12832 2651 12835
rect 3436 12832 3464 12863
rect 5442 12860 5448 12872
rect 5500 12860 5506 12912
rect 7006 12900 7012 12912
rect 5552 12872 7012 12900
rect 4062 12832 4068 12844
rect 2639 12804 2673 12832
rect 3436 12804 4068 12832
rect 2639 12801 2651 12804
rect 2593 12795 2651 12801
rect 4062 12792 4068 12804
rect 4120 12832 4126 12844
rect 4157 12835 4215 12841
rect 4157 12832 4169 12835
rect 4120 12804 4169 12832
rect 4120 12792 4126 12804
rect 4157 12801 4169 12804
rect 4203 12801 4215 12835
rect 5552 12832 5580 12872
rect 7006 12860 7012 12872
rect 7064 12860 7070 12912
rect 8386 12900 8392 12912
rect 8347 12872 8392 12900
rect 8386 12860 8392 12872
rect 8444 12860 8450 12912
rect 15657 12903 15715 12909
rect 15657 12900 15669 12903
rect 9416 12872 15669 12900
rect 4157 12795 4215 12801
rect 4264 12804 5580 12832
rect 5813 12835 5871 12841
rect 3786 12724 3792 12776
rect 3844 12764 3850 12776
rect 3973 12767 4031 12773
rect 3973 12764 3985 12767
rect 3844 12736 3985 12764
rect 3844 12724 3850 12736
rect 3973 12733 3985 12736
rect 4019 12733 4031 12767
rect 3973 12727 4031 12733
rect 4062 12696 4068 12708
rect 4023 12668 4068 12696
rect 4062 12656 4068 12668
rect 4120 12656 4126 12708
rect 2406 12628 2412 12640
rect 2367 12600 2412 12628
rect 2406 12588 2412 12600
rect 2464 12588 2470 12640
rect 2501 12631 2559 12637
rect 2501 12597 2513 12631
rect 2547 12628 2559 12631
rect 2682 12628 2688 12640
rect 2547 12600 2688 12628
rect 2547 12597 2559 12600
rect 2501 12591 2559 12597
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 3602 12588 3608 12640
rect 3660 12628 3666 12640
rect 4264 12628 4292 12804
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 5994 12832 6000 12844
rect 5859 12804 6000 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 5994 12792 6000 12804
rect 6052 12832 6058 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 6052 12804 7389 12832
rect 6052 12792 6058 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 8478 12792 8484 12844
rect 8536 12832 8542 12844
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 8536 12804 8953 12832
rect 8536 12792 8542 12804
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 5350 12724 5356 12776
rect 5408 12764 5414 12776
rect 5537 12767 5595 12773
rect 5537 12764 5549 12767
rect 5408 12736 5549 12764
rect 5408 12724 5414 12736
rect 5537 12733 5549 12736
rect 5583 12733 5595 12767
rect 5537 12727 5595 12733
rect 6086 12724 6092 12776
rect 6144 12764 6150 12776
rect 6546 12764 6552 12776
rect 6144 12736 6552 12764
rect 6144 12724 6150 12736
rect 6546 12724 6552 12736
rect 6604 12724 6610 12776
rect 7282 12764 7288 12776
rect 7208 12736 7288 12764
rect 7208 12705 7236 12736
rect 7282 12724 7288 12736
rect 7340 12764 7346 12776
rect 7837 12767 7895 12773
rect 7837 12764 7849 12767
rect 7340 12736 7849 12764
rect 7340 12724 7346 12736
rect 7837 12733 7849 12736
rect 7883 12733 7895 12767
rect 7837 12727 7895 12733
rect 8297 12767 8355 12773
rect 8297 12733 8309 12767
rect 8343 12764 8355 12767
rect 8386 12764 8392 12776
rect 8343 12736 8392 12764
rect 8343 12733 8355 12736
rect 8297 12727 8355 12733
rect 8386 12724 8392 12736
rect 8444 12764 8450 12776
rect 8757 12767 8815 12773
rect 8757 12764 8769 12767
rect 8444 12736 8769 12764
rect 8444 12724 8450 12736
rect 8757 12733 8769 12736
rect 8803 12764 8815 12767
rect 9416 12764 9444 12872
rect 15657 12869 15669 12872
rect 15703 12900 15715 12903
rect 16298 12900 16304 12912
rect 15703 12872 16304 12900
rect 15703 12869 15715 12872
rect 15657 12863 15715 12869
rect 16298 12860 16304 12872
rect 16356 12860 16362 12912
rect 10594 12832 10600 12844
rect 10555 12804 10600 12832
rect 10594 12792 10600 12804
rect 10652 12792 10658 12844
rect 12802 12792 12808 12844
rect 12860 12832 12866 12844
rect 13449 12835 13507 12841
rect 13449 12832 13461 12835
rect 12860 12804 13461 12832
rect 12860 12792 12866 12804
rect 13449 12801 13461 12804
rect 13495 12801 13507 12835
rect 13449 12795 13507 12801
rect 13633 12835 13691 12841
rect 13633 12801 13645 12835
rect 13679 12832 13691 12835
rect 13906 12832 13912 12844
rect 13679 12804 13912 12832
rect 13679 12801 13691 12804
rect 13633 12795 13691 12801
rect 8803 12736 9444 12764
rect 8803 12733 8815 12736
rect 8757 12727 8815 12733
rect 9950 12724 9956 12776
rect 10008 12724 10014 12776
rect 11238 12724 11244 12776
rect 11296 12764 11302 12776
rect 12161 12767 12219 12773
rect 12161 12764 12173 12767
rect 11296 12736 12173 12764
rect 11296 12724 11302 12736
rect 12161 12733 12173 12736
rect 12207 12764 12219 12767
rect 13262 12764 13268 12776
rect 12207 12736 13268 12764
rect 12207 12733 12219 12736
rect 12161 12727 12219 12733
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 13464 12764 13492 12795
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 14642 12792 14648 12844
rect 14700 12832 14706 12844
rect 16684 12841 16712 12940
rect 18414 12928 18420 12940
rect 18472 12928 18478 12980
rect 18785 12971 18843 12977
rect 18785 12937 18797 12971
rect 18831 12968 18843 12971
rect 18874 12968 18880 12980
rect 18831 12940 18880 12968
rect 18831 12937 18843 12940
rect 18785 12931 18843 12937
rect 18874 12928 18880 12940
rect 18932 12968 18938 12980
rect 19242 12968 19248 12980
rect 18932 12940 19248 12968
rect 18932 12928 18938 12940
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 19794 12928 19800 12980
rect 19852 12928 19858 12980
rect 20530 12928 20536 12980
rect 20588 12968 20594 12980
rect 20714 12968 20720 12980
rect 20588 12940 20720 12968
rect 20588 12928 20594 12940
rect 20714 12928 20720 12940
rect 20772 12928 20778 12980
rect 20898 12928 20904 12980
rect 20956 12968 20962 12980
rect 21361 12971 21419 12977
rect 21361 12968 21373 12971
rect 20956 12940 21373 12968
rect 20956 12928 20962 12940
rect 21361 12937 21373 12940
rect 21407 12937 21419 12971
rect 22738 12968 22744 12980
rect 22699 12940 22744 12968
rect 21361 12931 21419 12937
rect 22738 12928 22744 12940
rect 22796 12928 22802 12980
rect 23382 12928 23388 12980
rect 23440 12968 23446 12980
rect 23477 12971 23535 12977
rect 23477 12968 23489 12971
rect 23440 12940 23489 12968
rect 23440 12928 23446 12940
rect 23477 12937 23489 12940
rect 23523 12937 23535 12971
rect 23477 12931 23535 12937
rect 23661 12971 23719 12977
rect 23661 12937 23673 12971
rect 23707 12968 23719 12971
rect 24118 12968 24124 12980
rect 23707 12940 24124 12968
rect 23707 12937 23719 12940
rect 23661 12931 23719 12937
rect 24118 12928 24124 12940
rect 24176 12928 24182 12980
rect 24854 12928 24860 12980
rect 24912 12968 24918 12980
rect 25409 12971 25467 12977
rect 25409 12968 25421 12971
rect 24912 12940 25421 12968
rect 24912 12928 24918 12940
rect 25409 12937 25421 12940
rect 25455 12937 25467 12971
rect 25409 12931 25467 12937
rect 17494 12900 17500 12912
rect 17455 12872 17500 12900
rect 17494 12860 17500 12872
rect 17552 12860 17558 12912
rect 17586 12860 17592 12912
rect 17644 12900 17650 12912
rect 18322 12900 18328 12912
rect 17644 12872 18328 12900
rect 17644 12860 17650 12872
rect 18322 12860 18328 12872
rect 18380 12860 18386 12912
rect 19812 12900 19840 12928
rect 20993 12903 21051 12909
rect 20993 12900 21005 12903
rect 19812 12872 21005 12900
rect 20993 12869 21005 12872
rect 21039 12869 21051 12903
rect 20993 12863 21051 12869
rect 21542 12860 21548 12912
rect 21600 12900 21606 12912
rect 22002 12900 22008 12912
rect 21600 12872 22008 12900
rect 21600 12860 21606 12872
rect 22002 12860 22008 12872
rect 22060 12860 22066 12912
rect 22370 12860 22376 12912
rect 22428 12900 22434 12912
rect 23017 12903 23075 12909
rect 23017 12900 23029 12903
rect 22428 12872 23029 12900
rect 22428 12860 22434 12872
rect 23017 12869 23029 12872
rect 23063 12900 23075 12903
rect 23201 12903 23259 12909
rect 23201 12900 23213 12903
rect 23063 12872 23213 12900
rect 23063 12869 23075 12872
rect 23017 12863 23075 12869
rect 23201 12869 23213 12872
rect 23247 12869 23259 12903
rect 23201 12863 23259 12869
rect 23290 12860 23296 12912
rect 23348 12900 23354 12912
rect 23842 12900 23848 12912
rect 23348 12872 23848 12900
rect 23348 12860 23354 12872
rect 23842 12860 23848 12872
rect 23900 12860 23906 12912
rect 24486 12900 24492 12912
rect 24136 12872 24492 12900
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 14700 12804 15117 12832
rect 14700 12792 14706 12804
rect 15105 12801 15117 12804
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 16669 12835 16727 12841
rect 16669 12801 16681 12835
rect 16715 12801 16727 12835
rect 16669 12795 16727 12801
rect 16758 12792 16764 12844
rect 16816 12832 16822 12844
rect 16816 12804 16861 12832
rect 16816 12792 16822 12804
rect 19978 12792 19984 12844
rect 20036 12832 20042 12844
rect 20254 12832 20260 12844
rect 20036 12804 20260 12832
rect 20036 12792 20042 12804
rect 20254 12792 20260 12804
rect 20312 12792 20318 12844
rect 20806 12792 20812 12844
rect 20864 12832 20870 12844
rect 21821 12835 21879 12841
rect 21821 12832 21833 12835
rect 20864 12804 21833 12832
rect 20864 12792 20870 12804
rect 21821 12801 21833 12804
rect 21867 12801 21879 12835
rect 21821 12795 21879 12801
rect 21913 12835 21971 12841
rect 21913 12801 21925 12835
rect 21959 12801 21971 12835
rect 21913 12795 21971 12801
rect 14001 12767 14059 12773
rect 14001 12764 14013 12767
rect 13464 12736 14013 12764
rect 14001 12733 14013 12736
rect 14047 12733 14059 12767
rect 14001 12727 14059 12733
rect 14366 12724 14372 12776
rect 14424 12764 14430 12776
rect 15013 12767 15071 12773
rect 15013 12764 15025 12767
rect 14424 12736 15025 12764
rect 14424 12724 14430 12736
rect 15013 12733 15025 12736
rect 15059 12733 15071 12767
rect 16574 12764 16580 12776
rect 16535 12736 16580 12764
rect 15013 12727 15071 12733
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 18877 12767 18935 12773
rect 18877 12733 18889 12767
rect 18923 12764 18935 12767
rect 18966 12764 18972 12776
rect 18923 12736 18972 12764
rect 18923 12733 18935 12736
rect 18877 12727 18935 12733
rect 18966 12724 18972 12736
rect 19024 12724 19030 12776
rect 19426 12724 19432 12776
rect 19484 12764 19490 12776
rect 20162 12764 20168 12776
rect 19484 12736 20168 12764
rect 19484 12724 19490 12736
rect 20162 12724 20168 12736
rect 20220 12764 20226 12776
rect 20898 12764 20904 12776
rect 20220 12736 20904 12764
rect 20220 12724 20226 12736
rect 20898 12724 20904 12736
rect 20956 12724 20962 12776
rect 21174 12724 21180 12776
rect 21232 12764 21238 12776
rect 21928 12764 21956 12795
rect 22830 12792 22836 12844
rect 22888 12832 22894 12844
rect 24136 12841 24164 12872
rect 24486 12860 24492 12872
rect 24544 12860 24550 12912
rect 25038 12900 25044 12912
rect 24999 12872 25044 12900
rect 25038 12860 25044 12872
rect 25096 12860 25102 12912
rect 24121 12835 24179 12841
rect 24121 12832 24133 12835
rect 22888 12804 24133 12832
rect 22888 12792 22894 12804
rect 24121 12801 24133 12804
rect 24167 12801 24179 12835
rect 24121 12795 24179 12801
rect 24213 12835 24271 12841
rect 24213 12801 24225 12835
rect 24259 12801 24271 12835
rect 24213 12795 24271 12801
rect 21232 12736 21956 12764
rect 21232 12724 21238 12736
rect 23106 12724 23112 12776
rect 23164 12764 23170 12776
rect 23290 12764 23296 12776
rect 23164 12736 23296 12764
rect 23164 12724 23170 12736
rect 23290 12724 23296 12736
rect 23348 12724 23354 12776
rect 24026 12724 24032 12776
rect 24084 12724 24090 12776
rect 5077 12699 5135 12705
rect 5077 12665 5089 12699
rect 5123 12696 5135 12699
rect 7193 12699 7251 12705
rect 5123 12668 5672 12696
rect 5123 12665 5135 12668
rect 5077 12659 5135 12665
rect 3660 12600 4292 12628
rect 5169 12631 5227 12637
rect 3660 12588 3666 12600
rect 5169 12597 5181 12631
rect 5215 12628 5227 12631
rect 5442 12628 5448 12640
rect 5215 12600 5448 12628
rect 5215 12597 5227 12600
rect 5169 12591 5227 12597
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 5644 12637 5672 12668
rect 7193 12665 7205 12699
rect 7239 12665 7251 12699
rect 7193 12659 7251 12665
rect 9861 12699 9919 12705
rect 9861 12665 9873 12699
rect 9907 12696 9919 12699
rect 9968 12696 9996 12724
rect 10413 12699 10471 12705
rect 10413 12696 10425 12699
rect 9907 12668 10425 12696
rect 9907 12665 9919 12668
rect 9861 12659 9919 12665
rect 10413 12665 10425 12668
rect 10459 12665 10471 12699
rect 10413 12659 10471 12665
rect 11333 12699 11391 12705
rect 11333 12665 11345 12699
rect 11379 12696 11391 12699
rect 11882 12696 11888 12708
rect 11379 12668 11888 12696
rect 11379 12665 11391 12668
rect 11333 12659 11391 12665
rect 11882 12656 11888 12668
rect 11940 12656 11946 12708
rect 13446 12696 13452 12708
rect 13004 12668 13452 12696
rect 5629 12631 5687 12637
rect 5629 12597 5641 12631
rect 5675 12628 5687 12631
rect 5718 12628 5724 12640
rect 5675 12600 5724 12628
rect 5675 12597 5687 12600
rect 5629 12591 5687 12597
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 6270 12588 6276 12640
rect 6328 12628 6334 12640
rect 6365 12631 6423 12637
rect 6365 12628 6377 12631
rect 6328 12600 6377 12628
rect 6328 12588 6334 12600
rect 6365 12597 6377 12600
rect 6411 12597 6423 12631
rect 6822 12628 6828 12640
rect 6783 12600 6828 12628
rect 6365 12591 6423 12597
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 7282 12628 7288 12640
rect 7243 12600 7288 12628
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 8846 12588 8852 12640
rect 8904 12628 8910 12640
rect 8904 12600 8949 12628
rect 8904 12588 8910 12600
rect 10042 12588 10048 12640
rect 10100 12628 10106 12640
rect 13004 12637 13032 12668
rect 13446 12656 13452 12668
rect 13504 12656 13510 12708
rect 14918 12696 14924 12708
rect 14831 12668 14924 12696
rect 14918 12656 14924 12668
rect 14976 12696 14982 12708
rect 15562 12696 15568 12708
rect 14976 12668 15568 12696
rect 14976 12656 14982 12668
rect 15562 12656 15568 12668
rect 15620 12656 15626 12708
rect 19150 12705 19156 12708
rect 19144 12696 19156 12705
rect 19111 12668 19156 12696
rect 19144 12659 19156 12668
rect 19150 12656 19156 12659
rect 19208 12656 19214 12708
rect 19610 12656 19616 12708
rect 19668 12696 19674 12708
rect 21726 12696 21732 12708
rect 19668 12668 20208 12696
rect 21687 12668 21732 12696
rect 19668 12656 19674 12668
rect 20180 12640 20208 12668
rect 21726 12656 21732 12668
rect 21784 12696 21790 12708
rect 22094 12696 22100 12708
rect 21784 12668 22100 12696
rect 21784 12656 21790 12668
rect 22094 12656 22100 12668
rect 22152 12656 22158 12708
rect 23474 12656 23480 12708
rect 23532 12696 23538 12708
rect 24044 12696 24072 12724
rect 24228 12696 24256 12795
rect 24302 12724 24308 12776
rect 24360 12764 24366 12776
rect 25038 12764 25044 12776
rect 24360 12736 25044 12764
rect 24360 12724 24366 12736
rect 25038 12724 25044 12736
rect 25096 12764 25102 12776
rect 25225 12767 25283 12773
rect 25225 12764 25237 12767
rect 25096 12736 25237 12764
rect 25096 12724 25102 12736
rect 25225 12733 25237 12736
rect 25271 12764 25283 12767
rect 25777 12767 25835 12773
rect 25777 12764 25789 12767
rect 25271 12736 25789 12764
rect 25271 12733 25283 12736
rect 25225 12727 25283 12733
rect 25777 12733 25789 12736
rect 25823 12733 25835 12767
rect 25777 12727 25835 12733
rect 23532 12668 24256 12696
rect 23532 12656 23538 12668
rect 10321 12631 10379 12637
rect 10321 12628 10333 12631
rect 10100 12600 10333 12628
rect 10100 12588 10106 12600
rect 10321 12597 10333 12600
rect 10367 12597 10379 12631
rect 10321 12591 10379 12597
rect 12989 12631 13047 12637
rect 12989 12597 13001 12631
rect 13035 12597 13047 12631
rect 13354 12628 13360 12640
rect 13315 12600 13360 12628
rect 12989 12591 13047 12597
rect 13354 12588 13360 12600
rect 13412 12588 13418 12640
rect 14550 12628 14556 12640
rect 14511 12600 14556 12628
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 16206 12628 16212 12640
rect 16167 12600 16212 12628
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 16298 12588 16304 12640
rect 16356 12628 16362 12640
rect 16942 12628 16948 12640
rect 16356 12600 16948 12628
rect 16356 12588 16362 12600
rect 16942 12588 16948 12600
rect 17000 12628 17006 12640
rect 18414 12628 18420 12640
rect 17000 12600 18420 12628
rect 17000 12588 17006 12600
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 20162 12588 20168 12640
rect 20220 12588 20226 12640
rect 20257 12631 20315 12637
rect 20257 12597 20269 12631
rect 20303 12628 20315 12631
rect 20714 12628 20720 12640
rect 20303 12600 20720 12628
rect 20303 12597 20315 12600
rect 20257 12591 20315 12597
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 20806 12588 20812 12640
rect 20864 12628 20870 12640
rect 21082 12628 21088 12640
rect 20864 12600 21088 12628
rect 20864 12588 20870 12600
rect 21082 12588 21088 12600
rect 21140 12588 21146 12640
rect 23201 12631 23259 12637
rect 23201 12597 23213 12631
rect 23247 12628 23259 12631
rect 24029 12631 24087 12637
rect 24029 12628 24041 12631
rect 23247 12600 24041 12628
rect 23247 12597 23259 12600
rect 23201 12591 23259 12597
rect 24029 12597 24041 12600
rect 24075 12628 24087 12631
rect 25314 12628 25320 12640
rect 24075 12600 25320 12628
rect 24075 12597 24087 12600
rect 24029 12591 24087 12597
rect 25314 12588 25320 12600
rect 25372 12588 25378 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 2130 12424 2136 12436
rect 2091 12396 2136 12424
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 4246 12424 4252 12436
rect 4207 12396 4252 12424
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 5442 12384 5448 12436
rect 5500 12424 5506 12436
rect 5500 12396 5948 12424
rect 5500 12384 5506 12396
rect 842 12316 848 12368
rect 900 12356 906 12368
rect 2038 12356 2044 12368
rect 900 12328 2044 12356
rect 900 12316 906 12328
rect 2038 12316 2044 12328
rect 2096 12356 2102 12368
rect 2777 12359 2835 12365
rect 2777 12356 2789 12359
rect 2096 12328 2789 12356
rect 2096 12316 2102 12328
rect 2777 12325 2789 12328
rect 2823 12325 2835 12359
rect 2777 12319 2835 12325
rect 2869 12359 2927 12365
rect 2869 12325 2881 12359
rect 2915 12356 2927 12359
rect 3786 12356 3792 12368
rect 2915 12328 3792 12356
rect 2915 12325 2927 12328
rect 2869 12319 2927 12325
rect 1762 12248 1768 12300
rect 1820 12288 1826 12300
rect 2884 12288 2912 12319
rect 3786 12316 3792 12328
rect 3844 12316 3850 12368
rect 5534 12356 5540 12368
rect 3896 12328 5540 12356
rect 1820 12260 2912 12288
rect 1820 12248 1826 12260
rect 2608 12232 2636 12260
rect 3142 12248 3148 12300
rect 3200 12288 3206 12300
rect 3513 12291 3571 12297
rect 3513 12288 3525 12291
rect 3200 12260 3525 12288
rect 3200 12248 3206 12260
rect 3513 12257 3525 12260
rect 3559 12288 3571 12291
rect 3896 12288 3924 12328
rect 5534 12316 5540 12328
rect 5592 12316 5598 12368
rect 3559 12260 3924 12288
rect 3559 12257 3571 12260
rect 3513 12251 3571 12257
rect 4062 12248 4068 12300
rect 4120 12288 4126 12300
rect 5920 12297 5948 12396
rect 5994 12384 6000 12436
rect 6052 12424 6058 12436
rect 6457 12427 6515 12433
rect 6457 12424 6469 12427
rect 6052 12396 6469 12424
rect 6052 12384 6058 12396
rect 6457 12393 6469 12396
rect 6503 12424 6515 12427
rect 6730 12424 6736 12436
rect 6503 12396 6736 12424
rect 6503 12393 6515 12396
rect 6457 12387 6515 12393
rect 6730 12384 6736 12396
rect 6788 12384 6794 12436
rect 7006 12424 7012 12436
rect 6967 12396 7012 12424
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 8202 12424 8208 12436
rect 7116 12396 8208 12424
rect 6914 12316 6920 12368
rect 6972 12356 6978 12368
rect 7116 12356 7144 12396
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 9030 12424 9036 12436
rect 8991 12396 9036 12424
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 9306 12384 9312 12436
rect 9364 12424 9370 12436
rect 9401 12427 9459 12433
rect 9401 12424 9413 12427
rect 9364 12396 9413 12424
rect 9364 12384 9370 12396
rect 9401 12393 9413 12396
rect 9447 12393 9459 12427
rect 9401 12387 9459 12393
rect 9674 12384 9680 12436
rect 9732 12424 9738 12436
rect 10042 12424 10048 12436
rect 9732 12396 10048 12424
rect 9732 12384 9738 12396
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 10321 12427 10379 12433
rect 10321 12393 10333 12427
rect 10367 12424 10379 12427
rect 11054 12424 11060 12436
rect 10367 12396 11060 12424
rect 10367 12393 10379 12396
rect 10321 12387 10379 12393
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 11422 12424 11428 12436
rect 11383 12396 11428 12424
rect 11422 12384 11428 12396
rect 11480 12384 11486 12436
rect 11698 12424 11704 12436
rect 11659 12396 11704 12424
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 12250 12384 12256 12436
rect 12308 12424 12314 12436
rect 14645 12427 14703 12433
rect 14645 12424 14657 12427
rect 12308 12396 14657 12424
rect 12308 12384 12314 12396
rect 14645 12393 14657 12396
rect 14691 12424 14703 12427
rect 14918 12424 14924 12436
rect 14691 12396 14924 12424
rect 14691 12393 14703 12396
rect 14645 12387 14703 12393
rect 14918 12384 14924 12396
rect 14976 12384 14982 12436
rect 15105 12427 15163 12433
rect 15105 12393 15117 12427
rect 15151 12424 15163 12427
rect 15194 12424 15200 12436
rect 15151 12396 15200 12424
rect 15151 12393 15163 12396
rect 15105 12387 15163 12393
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 15746 12384 15752 12436
rect 15804 12424 15810 12436
rect 16025 12427 16083 12433
rect 16025 12424 16037 12427
rect 15804 12396 16037 12424
rect 15804 12384 15810 12396
rect 16025 12393 16037 12396
rect 16071 12393 16083 12427
rect 16025 12387 16083 12393
rect 17589 12427 17647 12433
rect 17589 12393 17601 12427
rect 17635 12424 17647 12427
rect 17862 12424 17868 12436
rect 17635 12396 17868 12424
rect 17635 12393 17647 12396
rect 17589 12387 17647 12393
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 18966 12424 18972 12436
rect 18927 12396 18972 12424
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 19061 12427 19119 12433
rect 19061 12393 19073 12427
rect 19107 12393 19119 12427
rect 19061 12387 19119 12393
rect 6972 12328 7144 12356
rect 7469 12359 7527 12365
rect 6972 12316 6978 12328
rect 7469 12325 7481 12359
rect 7515 12356 7527 12359
rect 7558 12356 7564 12368
rect 7515 12328 7564 12356
rect 7515 12325 7527 12328
rect 7469 12319 7527 12325
rect 7558 12316 7564 12328
rect 7616 12316 7622 12368
rect 19076 12300 19104 12387
rect 19334 12384 19340 12436
rect 19392 12384 19398 12436
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 19484 12396 19529 12424
rect 19484 12384 19490 12396
rect 21174 12384 21180 12436
rect 21232 12424 21238 12436
rect 21361 12427 21419 12433
rect 21361 12424 21373 12427
rect 21232 12396 21373 12424
rect 21232 12384 21238 12396
rect 21361 12393 21373 12396
rect 21407 12393 21419 12427
rect 21361 12387 21419 12393
rect 21821 12427 21879 12433
rect 21821 12393 21833 12427
rect 21867 12393 21879 12427
rect 21821 12387 21879 12393
rect 5813 12291 5871 12297
rect 4120 12260 4165 12288
rect 4120 12248 4126 12260
rect 5813 12257 5825 12291
rect 5859 12257 5871 12291
rect 5813 12251 5871 12257
rect 5905 12291 5963 12297
rect 5905 12257 5917 12291
rect 5951 12288 5963 12291
rect 6086 12288 6092 12300
rect 5951 12260 6092 12288
rect 5951 12257 5963 12260
rect 5905 12251 5963 12257
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12220 1455 12223
rect 2314 12220 2320 12232
rect 1443 12192 2320 12220
rect 1443 12189 1455 12192
rect 1397 12183 1455 12189
rect 2314 12180 2320 12192
rect 2372 12180 2378 12232
rect 2590 12180 2596 12232
rect 2648 12180 2654 12232
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 3418 12220 3424 12232
rect 3099 12192 3424 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 3418 12180 3424 12192
rect 3476 12220 3482 12232
rect 3878 12220 3884 12232
rect 3476 12192 3884 12220
rect 3476 12180 3482 12192
rect 3878 12180 3884 12192
rect 3936 12180 3942 12232
rect 4338 12180 4344 12232
rect 4396 12220 4402 12232
rect 4614 12220 4620 12232
rect 4396 12192 4620 12220
rect 4396 12180 4402 12192
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 5350 12220 5356 12232
rect 5184 12192 5356 12220
rect 2406 12152 2412 12164
rect 2367 12124 2412 12152
rect 2406 12112 2412 12124
rect 2464 12112 2470 12164
rect 5184 12161 5212 12192
rect 5350 12180 5356 12192
rect 5408 12180 5414 12232
rect 5169 12155 5227 12161
rect 5169 12152 5181 12155
rect 3712 12124 5181 12152
rect 1394 12044 1400 12096
rect 1452 12084 1458 12096
rect 3712 12084 3740 12124
rect 5169 12121 5181 12124
rect 5215 12121 5227 12155
rect 5442 12152 5448 12164
rect 5403 12124 5448 12152
rect 5169 12115 5227 12121
rect 5442 12112 5448 12124
rect 5500 12112 5506 12164
rect 5828 12152 5856 12251
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12288 6331 12291
rect 6822 12288 6828 12300
rect 6319 12260 6828 12288
rect 6319 12257 6331 12260
rect 6273 12251 6331 12257
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 7282 12288 7288 12300
rect 7064 12260 7288 12288
rect 7064 12248 7070 12260
rect 7282 12248 7288 12260
rect 7340 12248 7346 12300
rect 7377 12291 7435 12297
rect 7377 12257 7389 12291
rect 7423 12257 7435 12291
rect 7377 12251 7435 12257
rect 5997 12223 6055 12229
rect 5997 12189 6009 12223
rect 6043 12220 6055 12223
rect 6178 12220 6184 12232
rect 6043 12192 6184 12220
rect 6043 12189 6055 12192
rect 5997 12183 6055 12189
rect 6178 12180 6184 12192
rect 6236 12220 6242 12232
rect 6236 12192 7236 12220
rect 6236 12180 6242 12192
rect 6273 12155 6331 12161
rect 6273 12152 6285 12155
rect 5828 12124 6285 12152
rect 6273 12121 6285 12124
rect 6319 12121 6331 12155
rect 6273 12115 6331 12121
rect 3878 12084 3884 12096
rect 1452 12056 3740 12084
rect 3839 12056 3884 12084
rect 1452 12044 1458 12056
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 4614 12084 4620 12096
rect 4575 12056 4620 12084
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 6454 12044 6460 12096
rect 6512 12084 6518 12096
rect 6825 12087 6883 12093
rect 6825 12084 6837 12087
rect 6512 12056 6837 12084
rect 6512 12044 6518 12056
rect 6825 12053 6837 12056
rect 6871 12084 6883 12087
rect 7006 12084 7012 12096
rect 6871 12056 7012 12084
rect 6871 12053 6883 12056
rect 6825 12047 6883 12053
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 7208 12084 7236 12192
rect 7282 12112 7288 12164
rect 7340 12152 7346 12164
rect 7392 12152 7420 12251
rect 7742 12248 7748 12300
rect 7800 12288 7806 12300
rect 7926 12288 7932 12300
rect 7800 12260 7932 12288
rect 7800 12248 7806 12260
rect 7926 12248 7932 12260
rect 7984 12248 7990 12300
rect 8754 12248 8760 12300
rect 8812 12288 8818 12300
rect 9398 12288 9404 12300
rect 8812 12260 9404 12288
rect 8812 12248 8818 12260
rect 9398 12248 9404 12260
rect 9456 12248 9462 12300
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 9858 12288 9864 12300
rect 9640 12260 9864 12288
rect 9640 12248 9646 12260
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 10042 12248 10048 12300
rect 10100 12288 10106 12300
rect 10689 12291 10747 12297
rect 10689 12288 10701 12291
rect 10100 12260 10701 12288
rect 10100 12248 10106 12260
rect 10689 12257 10701 12260
rect 10735 12288 10747 12291
rect 10870 12288 10876 12300
rect 10735 12260 10876 12288
rect 10735 12257 10747 12260
rect 10689 12251 10747 12257
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 12158 12297 12164 12300
rect 12152 12288 12164 12297
rect 10980 12260 12164 12288
rect 7561 12223 7619 12229
rect 7561 12220 7573 12223
rect 7340 12124 7420 12152
rect 7484 12192 7573 12220
rect 7340 12112 7346 12124
rect 7484 12084 7512 12192
rect 7561 12189 7573 12192
rect 7607 12220 7619 12223
rect 8202 12220 8208 12232
rect 7607 12192 8208 12220
rect 7607 12189 7619 12192
rect 7561 12183 7619 12189
rect 8202 12180 8208 12192
rect 8260 12220 8266 12232
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 8260 12192 8401 12220
rect 8260 12180 8266 12192
rect 8389 12189 8401 12192
rect 8435 12220 8447 12223
rect 8478 12220 8484 12232
rect 8435 12192 8484 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12220 8631 12223
rect 9306 12220 9312 12232
rect 8619 12192 9312 12220
rect 8619 12189 8631 12192
rect 8573 12183 8631 12189
rect 9306 12180 9312 12192
rect 9364 12180 9370 12232
rect 10778 12220 10784 12232
rect 10739 12192 10784 12220
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 10980 12229 11008 12260
rect 12152 12251 12164 12260
rect 12216 12288 12222 12300
rect 16574 12288 16580 12300
rect 12216 12260 12252 12288
rect 16535 12260 16580 12288
rect 12158 12248 12164 12251
rect 12216 12248 12222 12260
rect 16574 12248 16580 12260
rect 16632 12248 16638 12300
rect 19058 12248 19064 12300
rect 19116 12248 19122 12300
rect 19352 12288 19380 12384
rect 20714 12356 20720 12368
rect 20675 12328 20720 12356
rect 20714 12316 20720 12328
rect 20772 12316 20778 12368
rect 21836 12356 21864 12387
rect 22094 12384 22100 12436
rect 22152 12424 22158 12436
rect 22833 12427 22891 12433
rect 22833 12424 22845 12427
rect 22152 12396 22845 12424
rect 22152 12384 22158 12396
rect 22833 12393 22845 12396
rect 22879 12393 22891 12427
rect 23382 12424 23388 12436
rect 23343 12396 23388 12424
rect 22833 12387 22891 12393
rect 23382 12384 23388 12396
rect 23440 12384 23446 12436
rect 23750 12424 23756 12436
rect 23711 12396 23756 12424
rect 23750 12384 23756 12396
rect 23808 12384 23814 12436
rect 23842 12384 23848 12436
rect 23900 12424 23906 12436
rect 24486 12424 24492 12436
rect 23900 12396 23945 12424
rect 24447 12396 24492 12424
rect 23900 12384 23906 12396
rect 24486 12384 24492 12396
rect 24544 12384 24550 12436
rect 24854 12384 24860 12436
rect 24912 12424 24918 12436
rect 25133 12427 25191 12433
rect 25133 12424 25145 12427
rect 24912 12396 25145 12424
rect 24912 12384 24918 12396
rect 25133 12393 25145 12396
rect 25179 12393 25191 12427
rect 25133 12387 25191 12393
rect 22646 12356 22652 12368
rect 21836 12328 22652 12356
rect 22646 12316 22652 12328
rect 22704 12316 22710 12368
rect 23293 12359 23351 12365
rect 23293 12325 23305 12359
rect 23339 12356 23351 12359
rect 23474 12356 23480 12368
rect 23339 12328 23480 12356
rect 23339 12325 23351 12328
rect 23293 12319 23351 12325
rect 23474 12316 23480 12328
rect 23532 12316 23538 12368
rect 19426 12288 19432 12300
rect 19352 12260 19432 12288
rect 19426 12248 19432 12260
rect 19484 12248 19490 12300
rect 21726 12248 21732 12300
rect 21784 12288 21790 12300
rect 22189 12291 22247 12297
rect 22189 12288 22201 12291
rect 21784 12260 22201 12288
rect 21784 12248 21790 12260
rect 22189 12257 22201 12260
rect 22235 12257 22247 12291
rect 24946 12288 24952 12300
rect 22189 12251 22247 12257
rect 23584 12260 24952 12288
rect 10965 12223 11023 12229
rect 10965 12189 10977 12223
rect 11011 12189 11023 12223
rect 11882 12220 11888 12232
rect 11843 12192 11888 12220
rect 10965 12183 11023 12189
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 16666 12220 16672 12232
rect 16627 12192 16672 12220
rect 16666 12180 16672 12192
rect 16724 12180 16730 12232
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12220 16911 12223
rect 17402 12220 17408 12232
rect 16899 12192 17408 12220
rect 16899 12189 16911 12192
rect 16853 12183 16911 12189
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 18046 12220 18052 12232
rect 18007 12192 18052 12220
rect 18046 12180 18052 12192
rect 18104 12180 18110 12232
rect 18414 12180 18420 12232
rect 18472 12220 18478 12232
rect 19242 12220 19248 12232
rect 18472 12192 19248 12220
rect 18472 12180 18478 12192
rect 19242 12180 19248 12192
rect 19300 12180 19306 12232
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12220 19579 12223
rect 19610 12220 19616 12232
rect 19567 12192 19616 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 19610 12180 19616 12192
rect 19668 12180 19674 12232
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12189 19763 12223
rect 22278 12220 22284 12232
rect 19705 12183 19763 12189
rect 20272 12192 22140 12220
rect 22239 12192 22284 12220
rect 9398 12112 9404 12164
rect 9456 12152 9462 12164
rect 9950 12152 9956 12164
rect 9456 12124 9956 12152
rect 9456 12112 9462 12124
rect 9950 12112 9956 12124
rect 10008 12112 10014 12164
rect 17957 12155 18015 12161
rect 17957 12121 17969 12155
rect 18003 12152 18015 12155
rect 18601 12155 18659 12161
rect 18601 12152 18613 12155
rect 18003 12124 18613 12152
rect 18003 12121 18015 12124
rect 17957 12115 18015 12121
rect 18601 12121 18613 12124
rect 18647 12152 18659 12155
rect 19150 12152 19156 12164
rect 18647 12124 19156 12152
rect 18647 12121 18659 12124
rect 18601 12115 18659 12121
rect 19150 12112 19156 12124
rect 19208 12152 19214 12164
rect 19720 12152 19748 12183
rect 19208 12124 19748 12152
rect 19208 12112 19214 12124
rect 8018 12084 8024 12096
rect 7208 12056 7512 12084
rect 7979 12056 8024 12084
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 13265 12087 13323 12093
rect 13265 12084 13277 12087
rect 13228 12056 13277 12084
rect 13228 12044 13234 12056
rect 13265 12053 13277 12056
rect 13311 12084 13323 12087
rect 13817 12087 13875 12093
rect 13817 12084 13829 12087
rect 13311 12056 13829 12084
rect 13311 12053 13323 12056
rect 13265 12047 13323 12053
rect 13817 12053 13829 12056
rect 13863 12053 13875 12087
rect 14182 12084 14188 12096
rect 14143 12056 14188 12084
rect 13817 12047 13875 12053
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 15562 12084 15568 12096
rect 15523 12056 15568 12084
rect 15562 12044 15568 12056
rect 15620 12044 15626 12096
rect 16206 12084 16212 12096
rect 16167 12056 16212 12084
rect 16206 12044 16212 12056
rect 16264 12044 16270 12096
rect 19242 12044 19248 12096
rect 19300 12084 19306 12096
rect 20272 12084 20300 12192
rect 21082 12112 21088 12164
rect 21140 12152 21146 12164
rect 21358 12152 21364 12164
rect 21140 12124 21364 12152
rect 21140 12112 21146 12124
rect 21358 12112 21364 12124
rect 21416 12112 21422 12164
rect 22112 12152 22140 12192
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 22465 12223 22523 12229
rect 22465 12189 22477 12223
rect 22511 12220 22523 12223
rect 23474 12220 23480 12232
rect 22511 12192 23480 12220
rect 22511 12189 22523 12192
rect 22465 12183 22523 12189
rect 23474 12180 23480 12192
rect 23532 12180 23538 12232
rect 23584 12152 23612 12260
rect 24946 12248 24952 12260
rect 25004 12248 25010 12300
rect 25590 12288 25596 12300
rect 25551 12260 25596 12288
rect 25590 12248 25596 12260
rect 25648 12248 25654 12300
rect 24026 12220 24032 12232
rect 23987 12192 24032 12220
rect 24026 12180 24032 12192
rect 24084 12180 24090 12232
rect 24857 12223 24915 12229
rect 24857 12189 24869 12223
rect 24903 12220 24915 12223
rect 25774 12220 25780 12232
rect 24903 12192 25780 12220
rect 24903 12189 24915 12192
rect 24857 12183 24915 12189
rect 25774 12180 25780 12192
rect 25832 12180 25838 12232
rect 22112 12124 23612 12152
rect 19300 12056 20300 12084
rect 20349 12087 20407 12093
rect 19300 12044 19306 12056
rect 20349 12053 20361 12087
rect 20395 12084 20407 12087
rect 21818 12084 21824 12096
rect 20395 12056 21824 12084
rect 20395 12053 20407 12056
rect 20349 12047 20407 12053
rect 21818 12044 21824 12056
rect 21876 12044 21882 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2590 11880 2596 11892
rect 2551 11852 2596 11880
rect 2590 11840 2596 11852
rect 2648 11840 2654 11892
rect 3142 11880 3148 11892
rect 2700 11852 3148 11880
rect 2700 11812 2728 11852
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 3568 11852 4559 11880
rect 3568 11840 3574 11852
rect 2240 11784 2728 11812
rect 2240 11753 2268 11784
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11713 2283 11747
rect 2225 11707 2283 11713
rect 1394 11636 1400 11688
rect 1452 11676 1458 11688
rect 1946 11676 1952 11688
rect 1452 11648 1952 11676
rect 1452 11636 1458 11648
rect 1946 11636 1952 11648
rect 2004 11636 2010 11688
rect 2041 11679 2099 11685
rect 2041 11645 2053 11679
rect 2087 11676 2099 11679
rect 2406 11676 2412 11688
rect 2087 11648 2412 11676
rect 2087 11645 2099 11648
rect 2041 11639 2099 11645
rect 2406 11636 2412 11648
rect 2464 11636 2470 11688
rect 3053 11679 3111 11685
rect 3053 11645 3065 11679
rect 3099 11676 3111 11679
rect 3145 11679 3203 11685
rect 3145 11676 3157 11679
rect 3099 11648 3157 11676
rect 3099 11645 3111 11648
rect 3053 11639 3111 11645
rect 3145 11645 3157 11648
rect 3191 11676 3203 11679
rect 4531 11676 4559 11852
rect 5534 11840 5540 11892
rect 5592 11880 5598 11892
rect 5813 11883 5871 11889
rect 5813 11880 5825 11883
rect 5592 11852 5825 11880
rect 5592 11840 5598 11852
rect 5813 11849 5825 11852
rect 5859 11849 5871 11883
rect 5813 11843 5871 11849
rect 6730 11840 6736 11892
rect 6788 11880 6794 11892
rect 7006 11880 7012 11892
rect 6788 11852 7012 11880
rect 6788 11840 6794 11852
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 8202 11880 8208 11892
rect 8163 11852 8208 11880
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 8570 11840 8576 11892
rect 8628 11880 8634 11892
rect 8757 11883 8815 11889
rect 8757 11880 8769 11883
rect 8628 11852 8769 11880
rect 8628 11840 8634 11852
rect 8757 11849 8769 11852
rect 8803 11849 8815 11883
rect 9122 11880 9128 11892
rect 9083 11852 9128 11880
rect 8757 11843 8815 11849
rect 9122 11840 9128 11852
rect 9180 11840 9186 11892
rect 13906 11840 13912 11892
rect 13964 11880 13970 11892
rect 14921 11883 14979 11889
rect 14921 11880 14933 11883
rect 13964 11852 14933 11880
rect 13964 11840 13970 11852
rect 14921 11849 14933 11852
rect 14967 11849 14979 11883
rect 15286 11880 15292 11892
rect 15247 11852 15292 11880
rect 14921 11843 14979 11849
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 17865 11883 17923 11889
rect 17865 11849 17877 11883
rect 17911 11880 17923 11883
rect 18966 11880 18972 11892
rect 17911 11852 18972 11880
rect 17911 11849 17923 11852
rect 17865 11843 17923 11849
rect 5350 11772 5356 11824
rect 5408 11812 5414 11824
rect 6086 11812 6092 11824
rect 5408 11784 6092 11812
rect 5408 11772 5414 11784
rect 6086 11772 6092 11784
rect 6144 11772 6150 11824
rect 6270 11772 6276 11824
rect 6328 11812 6334 11824
rect 6328 11784 6684 11812
rect 6328 11772 6334 11784
rect 5629 11679 5687 11685
rect 5629 11676 5641 11679
rect 3191 11648 4108 11676
rect 4531 11648 5641 11676
rect 3191 11645 3203 11648
rect 3145 11639 3203 11645
rect 3412 11611 3470 11617
rect 3412 11577 3424 11611
rect 3458 11608 3470 11611
rect 3878 11608 3884 11620
rect 3458 11580 3884 11608
rect 3458 11577 3470 11580
rect 3412 11571 3470 11577
rect 3878 11568 3884 11580
rect 3936 11568 3942 11620
rect 4080 11608 4108 11648
rect 5629 11645 5641 11648
rect 5675 11676 5687 11679
rect 6270 11676 6276 11688
rect 5675 11648 6276 11676
rect 5675 11645 5687 11648
rect 5629 11639 5687 11645
rect 6270 11636 6276 11648
rect 6328 11636 6334 11688
rect 6656 11685 6684 11784
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 15304 11744 15332 11840
rect 18064 11753 18092 11852
rect 18966 11840 18972 11852
rect 19024 11840 19030 11892
rect 20901 11883 20959 11889
rect 20901 11849 20913 11883
rect 20947 11880 20959 11883
rect 21634 11880 21640 11892
rect 20947 11852 21640 11880
rect 20947 11849 20959 11852
rect 20901 11843 20959 11849
rect 21634 11840 21640 11852
rect 21692 11840 21698 11892
rect 21818 11880 21824 11892
rect 21779 11852 21824 11880
rect 21818 11840 21824 11852
rect 21876 11880 21882 11892
rect 22278 11880 22284 11892
rect 21876 11852 22284 11880
rect 21876 11840 21882 11852
rect 22278 11840 22284 11852
rect 22336 11840 22342 11892
rect 22925 11883 22983 11889
rect 22925 11849 22937 11883
rect 22971 11880 22983 11883
rect 23477 11883 23535 11889
rect 23477 11880 23489 11883
rect 22971 11852 23489 11880
rect 22971 11849 22983 11852
rect 22925 11843 22983 11849
rect 23477 11849 23489 11852
rect 23523 11880 23535 11883
rect 24026 11880 24032 11892
rect 23523 11852 24032 11880
rect 23523 11849 23535 11852
rect 23477 11843 23535 11849
rect 24026 11840 24032 11852
rect 24084 11840 24090 11892
rect 24946 11880 24952 11892
rect 24907 11852 24952 11880
rect 24946 11840 24952 11852
rect 25004 11840 25010 11892
rect 25406 11880 25412 11892
rect 25367 11852 25412 11880
rect 25406 11840 25412 11852
rect 25464 11840 25470 11892
rect 25869 11883 25927 11889
rect 25869 11849 25881 11883
rect 25915 11880 25927 11883
rect 26050 11880 26056 11892
rect 25915 11852 26056 11880
rect 25915 11849 25927 11852
rect 25869 11843 25927 11849
rect 15473 11747 15531 11753
rect 15473 11744 15485 11747
rect 9548 11716 9996 11744
rect 9548 11704 9554 11716
rect 6641 11679 6699 11685
rect 6641 11645 6653 11679
rect 6687 11676 6699 11679
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6687 11648 6837 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 6825 11645 6837 11648
rect 6871 11676 6883 11679
rect 9861 11679 9919 11685
rect 9861 11676 9873 11679
rect 6871 11648 9873 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 9861 11645 9873 11648
rect 9907 11645 9919 11679
rect 9968 11676 9996 11716
rect 11072 11716 13124 11744
rect 15304 11716 15485 11744
rect 10128 11679 10186 11685
rect 10128 11676 10140 11679
rect 9968 11648 10140 11676
rect 9861 11639 9919 11645
rect 10128 11645 10140 11648
rect 10174 11676 10186 11679
rect 11072 11676 11100 11716
rect 10174 11648 11100 11676
rect 12989 11679 13047 11685
rect 10174 11645 10186 11648
rect 10128 11639 10186 11645
rect 12989 11645 13001 11679
rect 13035 11645 13047 11679
rect 13096 11676 13124 11716
rect 15473 11713 15485 11716
rect 15519 11713 15531 11747
rect 15473 11707 15531 11713
rect 18049 11747 18107 11753
rect 18049 11713 18061 11747
rect 18095 11713 18107 11747
rect 18049 11707 18107 11713
rect 14642 11676 14648 11688
rect 13096 11648 14648 11676
rect 12989 11639 13047 11645
rect 4246 11608 4252 11620
rect 4080 11580 4252 11608
rect 4246 11568 4252 11580
rect 4304 11568 4310 11620
rect 4798 11568 4804 11620
rect 4856 11608 4862 11620
rect 5077 11611 5135 11617
rect 5077 11608 5089 11611
rect 4856 11580 5089 11608
rect 4856 11568 4862 11580
rect 5077 11577 5089 11580
rect 5123 11577 5135 11611
rect 5077 11571 5135 11577
rect 7006 11568 7012 11620
rect 7064 11617 7070 11620
rect 7064 11611 7128 11617
rect 7064 11577 7082 11611
rect 7116 11577 7128 11611
rect 7064 11571 7128 11577
rect 9769 11611 9827 11617
rect 9769 11577 9781 11611
rect 9815 11608 9827 11611
rect 9876 11608 9904 11639
rect 9815 11580 11928 11608
rect 9815 11577 9827 11580
rect 9769 11571 9827 11577
rect 7064 11568 7070 11571
rect 11900 11552 11928 11580
rect 1581 11543 1639 11549
rect 1581 11509 1593 11543
rect 1627 11540 1639 11543
rect 1762 11540 1768 11552
rect 1627 11512 1768 11540
rect 1627 11509 1639 11512
rect 1581 11503 1639 11509
rect 1762 11500 1768 11512
rect 1820 11500 1826 11552
rect 4522 11540 4528 11552
rect 4483 11512 4528 11540
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 5537 11543 5595 11549
rect 5537 11509 5549 11543
rect 5583 11540 5595 11543
rect 6178 11540 6184 11552
rect 5583 11512 6184 11540
rect 5583 11509 5595 11512
rect 5537 11503 5595 11509
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 7190 11500 7196 11552
rect 7248 11540 7254 11552
rect 7742 11540 7748 11552
rect 7248 11512 7748 11540
rect 7248 11500 7254 11512
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11241 11543 11299 11549
rect 11241 11540 11253 11543
rect 10928 11512 11253 11540
rect 10928 11500 10934 11512
rect 11241 11509 11253 11512
rect 11287 11509 11299 11543
rect 11241 11503 11299 11509
rect 11882 11500 11888 11552
rect 11940 11540 11946 11552
rect 11977 11543 12035 11549
rect 11977 11540 11989 11543
rect 11940 11512 11989 11540
rect 11940 11500 11946 11512
rect 11977 11509 11989 11512
rect 12023 11540 12035 11543
rect 12897 11543 12955 11549
rect 12897 11540 12909 11543
rect 12023 11512 12909 11540
rect 12023 11509 12035 11512
rect 11977 11503 12035 11509
rect 12897 11509 12909 11512
rect 12943 11540 12955 11543
rect 13004 11540 13032 11639
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 15488 11676 15516 11707
rect 19518 11704 19524 11756
rect 19576 11744 19582 11756
rect 19978 11744 19984 11756
rect 19576 11716 19984 11744
rect 19576 11704 19582 11716
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 20441 11747 20499 11753
rect 20441 11713 20453 11747
rect 20487 11744 20499 11747
rect 20898 11744 20904 11756
rect 20487 11716 20904 11744
rect 20487 11713 20499 11716
rect 20441 11707 20499 11713
rect 20898 11704 20904 11716
rect 20956 11704 20962 11756
rect 21266 11744 21272 11756
rect 21227 11716 21272 11744
rect 21266 11704 21272 11716
rect 21324 11704 21330 11756
rect 21450 11704 21456 11756
rect 21508 11744 21514 11756
rect 21637 11747 21695 11753
rect 21637 11744 21649 11747
rect 21508 11716 21649 11744
rect 21508 11704 21514 11716
rect 21637 11713 21649 11716
rect 21683 11713 21695 11747
rect 21637 11707 21695 11713
rect 16206 11676 16212 11688
rect 15488 11648 16212 11676
rect 16206 11636 16212 11648
rect 16264 11636 16270 11688
rect 20714 11676 20720 11688
rect 20675 11648 20720 11676
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 13170 11568 13176 11620
rect 13228 11617 13234 11620
rect 13228 11611 13292 11617
rect 13228 11577 13246 11611
rect 13280 11577 13292 11611
rect 13228 11571 13292 11577
rect 13228 11568 13234 11571
rect 15562 11568 15568 11620
rect 15620 11608 15626 11620
rect 15718 11611 15776 11617
rect 15718 11608 15730 11611
rect 15620 11580 15730 11608
rect 15620 11568 15626 11580
rect 15718 11577 15730 11580
rect 15764 11577 15776 11611
rect 18294 11611 18352 11617
rect 18294 11608 18306 11611
rect 15718 11571 15776 11577
rect 17420 11580 18306 11608
rect 17420 11552 17448 11580
rect 18294 11577 18306 11580
rect 18340 11577 18352 11611
rect 18294 11571 18352 11577
rect 19242 11568 19248 11620
rect 19300 11608 19306 11620
rect 19610 11608 19616 11620
rect 19300 11580 19616 11608
rect 19300 11568 19306 11580
rect 19610 11568 19616 11580
rect 19668 11608 19674 11620
rect 19981 11611 20039 11617
rect 19981 11608 19993 11611
rect 19668 11580 19993 11608
rect 19668 11568 19674 11580
rect 19981 11577 19993 11580
rect 20027 11577 20039 11611
rect 19981 11571 20039 11577
rect 13814 11540 13820 11552
rect 12943 11512 13820 11540
rect 12943 11509 12955 11512
rect 12897 11503 12955 11509
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 14182 11500 14188 11552
rect 14240 11540 14246 11552
rect 14369 11543 14427 11549
rect 14369 11540 14381 11543
rect 14240 11512 14381 11540
rect 14240 11500 14246 11512
rect 14369 11509 14381 11512
rect 14415 11509 14427 11543
rect 16850 11540 16856 11552
rect 16811 11512 16856 11540
rect 14369 11503 14427 11509
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 17402 11540 17408 11552
rect 17363 11512 17408 11540
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 19150 11500 19156 11552
rect 19208 11540 19214 11552
rect 19426 11540 19432 11552
rect 19208 11512 19432 11540
rect 19208 11500 19214 11512
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 21652 11540 21680 11707
rect 22094 11704 22100 11756
rect 22152 11704 22158 11756
rect 22370 11744 22376 11756
rect 22331 11716 22376 11744
rect 22370 11704 22376 11716
rect 22428 11704 22434 11756
rect 23474 11704 23480 11756
rect 23532 11744 23538 11756
rect 24213 11747 24271 11753
rect 24213 11744 24225 11747
rect 23532 11716 24225 11744
rect 23532 11704 23538 11716
rect 24213 11713 24225 11716
rect 24259 11713 24271 11747
rect 24213 11707 24271 11713
rect 22112 11676 22140 11704
rect 25225 11679 25283 11685
rect 22112 11648 22324 11676
rect 22296 11617 22324 11648
rect 25225 11645 25237 11679
rect 25271 11676 25283 11679
rect 25884 11676 25912 11843
rect 26050 11840 26056 11852
rect 26108 11840 26114 11892
rect 26234 11812 26240 11824
rect 26195 11784 26240 11812
rect 26234 11772 26240 11784
rect 26292 11772 26298 11824
rect 25271 11648 25912 11676
rect 25271 11645 25283 11648
rect 25225 11639 25283 11645
rect 22281 11611 22339 11617
rect 22281 11577 22293 11611
rect 22327 11577 22339 11611
rect 22281 11571 22339 11577
rect 22189 11543 22247 11549
rect 22189 11540 22201 11543
rect 21652 11512 22201 11540
rect 22189 11509 22201 11512
rect 22235 11509 22247 11543
rect 22189 11503 22247 11509
rect 23382 11500 23388 11552
rect 23440 11540 23446 11552
rect 23661 11543 23719 11549
rect 23661 11540 23673 11543
rect 23440 11512 23673 11540
rect 23440 11500 23446 11512
rect 23661 11509 23673 11512
rect 23707 11509 23719 11543
rect 24026 11540 24032 11552
rect 23987 11512 24032 11540
rect 23661 11503 23719 11509
rect 24026 11500 24032 11512
rect 24084 11500 24090 11552
rect 24121 11543 24179 11549
rect 24121 11509 24133 11543
rect 24167 11540 24179 11543
rect 24394 11540 24400 11552
rect 24167 11512 24400 11540
rect 24167 11509 24179 11512
rect 24121 11503 24179 11509
rect 24394 11500 24400 11512
rect 24452 11500 24458 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1946 11336 1952 11348
rect 1907 11308 1952 11336
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 2038 11296 2044 11348
rect 2096 11336 2102 11348
rect 2225 11339 2283 11345
rect 2225 11336 2237 11339
rect 2096 11308 2237 11336
rect 2096 11296 2102 11308
rect 2225 11305 2237 11308
rect 2271 11305 2283 11339
rect 2866 11336 2872 11348
rect 2827 11308 2872 11336
rect 2225 11299 2283 11305
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3418 11336 3424 11348
rect 3379 11308 3424 11336
rect 3418 11296 3424 11308
rect 3476 11296 3482 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4341 11339 4399 11345
rect 4341 11336 4353 11339
rect 4120 11308 4353 11336
rect 4120 11296 4126 11308
rect 4341 11305 4353 11308
rect 4387 11336 4399 11339
rect 5350 11336 5356 11348
rect 4387 11308 5356 11336
rect 4387 11305 4399 11308
rect 4341 11299 4399 11305
rect 5350 11296 5356 11308
rect 5408 11296 5414 11348
rect 6270 11296 6276 11348
rect 6328 11336 6334 11348
rect 6365 11339 6423 11345
rect 6365 11336 6377 11339
rect 6328 11308 6377 11336
rect 6328 11296 6334 11308
rect 6365 11305 6377 11308
rect 6411 11305 6423 11339
rect 6365 11299 6423 11305
rect 6822 11296 6828 11348
rect 6880 11336 6886 11348
rect 6917 11339 6975 11345
rect 6917 11336 6929 11339
rect 6880 11308 6929 11336
rect 6880 11296 6886 11308
rect 6917 11305 6929 11308
rect 6963 11336 6975 11339
rect 7006 11336 7012 11348
rect 6963 11308 7012 11336
rect 6963 11305 6975 11308
rect 6917 11299 6975 11305
rect 7006 11296 7012 11308
rect 7064 11336 7070 11348
rect 7193 11339 7251 11345
rect 7193 11336 7205 11339
rect 7064 11308 7205 11336
rect 7064 11296 7070 11308
rect 7193 11305 7205 11308
rect 7239 11305 7251 11339
rect 7193 11299 7251 11305
rect 7653 11339 7711 11345
rect 7653 11305 7665 11339
rect 7699 11336 7711 11339
rect 8202 11336 8208 11348
rect 7699 11308 8208 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 1302 11228 1308 11280
rect 1360 11268 1366 11280
rect 1854 11268 1860 11280
rect 1360 11240 1860 11268
rect 1360 11228 1366 11240
rect 1854 11228 1860 11240
rect 1912 11268 1918 11280
rect 2777 11271 2835 11277
rect 2777 11268 2789 11271
rect 1912 11240 2789 11268
rect 1912 11228 1918 11240
rect 2777 11237 2789 11240
rect 2823 11268 2835 11271
rect 6454 11268 6460 11280
rect 2823 11240 6460 11268
rect 2823 11237 2835 11240
rect 2777 11231 2835 11237
rect 4246 11160 4252 11212
rect 4304 11200 4310 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4304 11172 4445 11200
rect 4304 11160 4310 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 4522 11160 4528 11212
rect 4580 11200 4586 11212
rect 4689 11203 4747 11209
rect 4689 11200 4701 11203
rect 4580 11172 4701 11200
rect 4580 11160 4586 11172
rect 4689 11169 4701 11172
rect 4735 11200 4747 11203
rect 5442 11200 5448 11212
rect 4735 11172 5448 11200
rect 4735 11169 4747 11172
rect 4689 11163 4747 11169
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 6196 11144 6224 11240
rect 6454 11228 6460 11240
rect 6512 11228 6518 11280
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 3142 11132 3148 11144
rect 3099 11104 3148 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 6178 11092 6184 11144
rect 6236 11092 6242 11144
rect 7208 11132 7236 11299
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 8294 11296 8300 11348
rect 8352 11336 8358 11348
rect 9309 11339 9367 11345
rect 9309 11336 9321 11339
rect 8352 11308 9321 11336
rect 8352 11296 8358 11308
rect 9309 11305 9321 11308
rect 9355 11305 9367 11339
rect 9309 11299 9367 11305
rect 9490 11296 9496 11348
rect 9548 11336 9554 11348
rect 9861 11339 9919 11345
rect 9861 11336 9873 11339
rect 9548 11308 9873 11336
rect 9548 11296 9554 11308
rect 9861 11305 9873 11308
rect 9907 11305 9919 11339
rect 9861 11299 9919 11305
rect 10321 11339 10379 11345
rect 10321 11305 10333 11339
rect 10367 11336 10379 11339
rect 11606 11336 11612 11348
rect 10367 11308 11612 11336
rect 10367 11305 10379 11308
rect 10321 11299 10379 11305
rect 11606 11296 11612 11308
rect 11664 11336 11670 11348
rect 11793 11339 11851 11345
rect 11793 11336 11805 11339
rect 11664 11308 11805 11336
rect 11664 11296 11670 11308
rect 11793 11305 11805 11308
rect 11839 11336 11851 11339
rect 12158 11336 12164 11348
rect 11839 11308 12164 11336
rect 11839 11305 11851 11308
rect 11793 11299 11851 11305
rect 12158 11296 12164 11308
rect 12216 11336 12222 11348
rect 12345 11339 12403 11345
rect 12345 11336 12357 11339
rect 12216 11308 12357 11336
rect 12216 11296 12222 11308
rect 12345 11305 12357 11308
rect 12391 11305 12403 11339
rect 12710 11336 12716 11348
rect 12671 11308 12716 11336
rect 12345 11299 12403 11305
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 12989 11339 13047 11345
rect 12989 11305 13001 11339
rect 13035 11336 13047 11339
rect 13262 11336 13268 11348
rect 13035 11308 13268 11336
rect 13035 11305 13047 11308
rect 12989 11299 13047 11305
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 13357 11339 13415 11345
rect 13357 11305 13369 11339
rect 13403 11336 13415 11339
rect 13538 11336 13544 11348
rect 13403 11308 13544 11336
rect 13403 11305 13415 11308
rect 13357 11299 13415 11305
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 14274 11296 14280 11348
rect 14332 11336 14338 11348
rect 14369 11339 14427 11345
rect 14369 11336 14381 11339
rect 14332 11308 14381 11336
rect 14332 11296 14338 11308
rect 14369 11305 14381 11308
rect 14415 11305 14427 11339
rect 14369 11299 14427 11305
rect 15473 11339 15531 11345
rect 15473 11305 15485 11339
rect 15519 11336 15531 11339
rect 15654 11336 15660 11348
rect 15519 11308 15660 11336
rect 15519 11305 15531 11308
rect 15473 11299 15531 11305
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 16301 11339 16359 11345
rect 16301 11305 16313 11339
rect 16347 11336 16359 11339
rect 17402 11336 17408 11348
rect 16347 11308 17408 11336
rect 16347 11305 16359 11308
rect 16301 11299 16359 11305
rect 17402 11296 17408 11308
rect 17460 11336 17466 11348
rect 17865 11339 17923 11345
rect 17865 11336 17877 11339
rect 17460 11308 17877 11336
rect 17460 11296 17466 11308
rect 17865 11305 17877 11308
rect 17911 11305 17923 11339
rect 17865 11299 17923 11305
rect 18969 11339 19027 11345
rect 18969 11305 18981 11339
rect 19015 11336 19027 11339
rect 19150 11336 19156 11348
rect 19015 11308 19156 11336
rect 19015 11305 19027 11308
rect 18969 11299 19027 11305
rect 19150 11296 19156 11308
rect 19208 11336 19214 11348
rect 20714 11336 20720 11348
rect 19208 11308 20720 11336
rect 19208 11296 19214 11308
rect 20714 11296 20720 11308
rect 20772 11296 20778 11348
rect 20898 11336 20904 11348
rect 20859 11308 20904 11336
rect 20898 11296 20904 11308
rect 20956 11296 20962 11348
rect 21266 11336 21272 11348
rect 21227 11308 21272 11336
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 22002 11336 22008 11348
rect 21963 11308 22008 11336
rect 22002 11296 22008 11308
rect 22060 11296 22066 11348
rect 22462 11336 22468 11348
rect 22423 11308 22468 11336
rect 22462 11296 22468 11308
rect 22520 11296 22526 11348
rect 23842 11296 23848 11348
rect 23900 11336 23906 11348
rect 24029 11339 24087 11345
rect 24029 11336 24041 11339
rect 23900 11308 24041 11336
rect 23900 11296 23906 11308
rect 24029 11305 24041 11308
rect 24075 11305 24087 11339
rect 24029 11299 24087 11305
rect 24210 11296 24216 11348
rect 24268 11336 24274 11348
rect 24765 11339 24823 11345
rect 24765 11336 24777 11339
rect 24268 11308 24777 11336
rect 24268 11296 24274 11308
rect 24765 11305 24777 11308
rect 24811 11305 24823 11339
rect 24765 11299 24823 11305
rect 24854 11296 24860 11348
rect 24912 11336 24918 11348
rect 25133 11339 25191 11345
rect 25133 11336 25145 11339
rect 24912 11308 25145 11336
rect 24912 11296 24918 11308
rect 25133 11305 25145 11308
rect 25179 11305 25191 11339
rect 25133 11299 25191 11305
rect 10680 11271 10738 11277
rect 10680 11237 10692 11271
rect 10726 11268 10738 11271
rect 10870 11268 10876 11280
rect 10726 11240 10876 11268
rect 10726 11237 10738 11240
rect 10680 11231 10738 11237
rect 10870 11228 10876 11240
rect 10928 11228 10934 11280
rect 15930 11268 15936 11280
rect 15843 11240 15936 11268
rect 15930 11228 15936 11240
rect 15988 11268 15994 11280
rect 16752 11271 16810 11277
rect 16752 11268 16764 11271
rect 15988 11240 16764 11268
rect 15988 11228 15994 11240
rect 16752 11237 16764 11240
rect 16798 11268 16810 11271
rect 16850 11268 16856 11280
rect 16798 11240 16856 11268
rect 16798 11237 16810 11240
rect 16752 11231 16810 11237
rect 16850 11228 16856 11240
rect 16908 11228 16914 11280
rect 19426 11228 19432 11280
rect 19484 11268 19490 11280
rect 22370 11268 22376 11280
rect 19484 11240 20760 11268
rect 22331 11240 22376 11268
rect 19484 11228 19490 11240
rect 7374 11160 7380 11212
rect 7432 11200 7438 11212
rect 8113 11203 8171 11209
rect 8113 11200 8125 11203
rect 7432 11172 8125 11200
rect 7432 11160 7438 11172
rect 8113 11169 8125 11172
rect 8159 11200 8171 11203
rect 8202 11200 8208 11212
rect 8159 11172 8208 11200
rect 8159 11169 8171 11172
rect 8113 11163 8171 11169
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 10410 11200 10416 11212
rect 10323 11172 10416 11200
rect 10410 11160 10416 11172
rect 10468 11200 10474 11212
rect 11882 11200 11888 11212
rect 10468 11172 11888 11200
rect 10468 11160 10474 11172
rect 11882 11160 11888 11172
rect 11940 11160 11946 11212
rect 15286 11200 15292 11212
rect 15247 11172 15292 11200
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 15470 11160 15476 11212
rect 15528 11200 15534 11212
rect 16298 11200 16304 11212
rect 15528 11172 16304 11200
rect 15528 11160 15534 11172
rect 16298 11160 16304 11172
rect 16356 11160 16362 11212
rect 18966 11160 18972 11212
rect 19024 11200 19030 11212
rect 19337 11203 19395 11209
rect 19337 11200 19349 11203
rect 19024 11172 19349 11200
rect 19024 11160 19030 11172
rect 19337 11169 19349 11172
rect 19383 11169 19395 11203
rect 19702 11200 19708 11212
rect 19337 11163 19395 11169
rect 19444 11172 19708 11200
rect 19444 11144 19472 11172
rect 19702 11160 19708 11172
rect 19760 11160 19766 11212
rect 19886 11160 19892 11212
rect 19944 11200 19950 11212
rect 20346 11200 20352 11212
rect 19944 11172 20352 11200
rect 19944 11160 19950 11172
rect 20346 11160 20352 11172
rect 20404 11160 20410 11212
rect 20732 11209 20760 11240
rect 22370 11228 22376 11240
rect 22428 11228 22434 11280
rect 23566 11228 23572 11280
rect 23624 11268 23630 11280
rect 24397 11271 24455 11277
rect 24397 11268 24409 11271
rect 23624 11240 24409 11268
rect 23624 11228 23630 11240
rect 24397 11237 24409 11240
rect 24443 11237 24455 11271
rect 24397 11231 24455 11237
rect 20717 11203 20775 11209
rect 20717 11169 20729 11203
rect 20763 11200 20775 11203
rect 20763 11172 21588 11200
rect 20763 11169 20775 11172
rect 20717 11163 20775 11169
rect 8297 11135 8355 11141
rect 8297 11132 8309 11135
rect 7208 11104 8309 11132
rect 8297 11101 8309 11104
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 12986 11092 12992 11144
rect 13044 11132 13050 11144
rect 13449 11135 13507 11141
rect 13449 11132 13461 11135
rect 13044 11104 13461 11132
rect 13044 11092 13050 11104
rect 13449 11101 13461 11104
rect 13495 11101 13507 11135
rect 13449 11095 13507 11101
rect 13633 11135 13691 11141
rect 13633 11101 13645 11135
rect 13679 11132 13691 11135
rect 14734 11132 14740 11144
rect 13679 11104 14136 11132
rect 14695 11104 14740 11132
rect 13679 11101 13691 11104
rect 13633 11095 13691 11101
rect 2130 11024 2136 11076
rect 2188 11064 2194 11076
rect 2409 11067 2467 11073
rect 2409 11064 2421 11067
rect 2188 11036 2421 11064
rect 2188 11024 2194 11036
rect 2409 11033 2421 11036
rect 2455 11033 2467 11067
rect 2409 11027 2467 11033
rect 5813 11067 5871 11073
rect 5813 11033 5825 11067
rect 5859 11064 5871 11067
rect 6086 11064 6092 11076
rect 5859 11036 6092 11064
rect 5859 11033 5871 11036
rect 5813 11027 5871 11033
rect 6086 11024 6092 11036
rect 6144 11024 6150 11076
rect 7745 11067 7803 11073
rect 7745 11033 7757 11067
rect 7791 11064 7803 11067
rect 8110 11064 8116 11076
rect 7791 11036 8116 11064
rect 7791 11033 7803 11036
rect 7745 11027 7803 11033
rect 8110 11024 8116 11036
rect 8168 11024 8174 11076
rect 3786 10996 3792 11008
rect 3747 10968 3792 10996
rect 3786 10956 3792 10968
rect 3844 10956 3850 11008
rect 9030 10996 9036 11008
rect 8991 10968 9036 10996
rect 9030 10956 9036 10968
rect 9088 10956 9094 11008
rect 12158 10956 12164 11008
rect 12216 10996 12222 11008
rect 12434 10996 12440 11008
rect 12216 10968 12440 10996
rect 12216 10956 12222 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 14108 11005 14136 11104
rect 14734 11092 14740 11104
rect 14792 11092 14798 11144
rect 16206 11092 16212 11144
rect 16264 11132 16270 11144
rect 16390 11132 16396 11144
rect 16264 11104 16396 11132
rect 16264 11092 16270 11104
rect 16390 11092 16396 11104
rect 16448 11132 16454 11144
rect 16485 11135 16543 11141
rect 16485 11132 16497 11135
rect 16448 11104 16497 11132
rect 16448 11092 16454 11104
rect 16485 11101 16497 11104
rect 16531 11101 16543 11135
rect 19426 11132 19432 11144
rect 19339 11104 19432 11132
rect 16485 11095 16543 11101
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 19521 11135 19579 11141
rect 19521 11101 19533 11135
rect 19567 11101 19579 11135
rect 19521 11095 19579 11101
rect 18874 11064 18880 11076
rect 18787 11036 18880 11064
rect 18874 11024 18880 11036
rect 18932 11064 18938 11076
rect 19536 11064 19564 11095
rect 21082 11092 21088 11144
rect 21140 11132 21146 11144
rect 21560 11141 21588 11172
rect 22738 11160 22744 11212
rect 22796 11200 22802 11212
rect 22833 11203 22891 11209
rect 22833 11200 22845 11203
rect 22796 11172 22845 11200
rect 22796 11160 22802 11172
rect 22833 11169 22845 11172
rect 22879 11169 22891 11203
rect 22833 11163 22891 11169
rect 24210 11160 24216 11212
rect 24268 11200 24274 11212
rect 24581 11203 24639 11209
rect 24581 11200 24593 11203
rect 24268 11172 24593 11200
rect 24268 11160 24274 11172
rect 24581 11169 24593 11172
rect 24627 11169 24639 11203
rect 24581 11163 24639 11169
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 21140 11104 21373 11132
rect 21140 11092 21146 11104
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 21361 11095 21419 11101
rect 21545 11135 21603 11141
rect 21545 11101 21557 11135
rect 21591 11132 21603 11135
rect 22002 11132 22008 11144
rect 21591 11104 22008 11132
rect 21591 11101 21603 11104
rect 21545 11095 21603 11101
rect 22002 11092 22008 11104
rect 22060 11092 22066 11144
rect 22922 11132 22928 11144
rect 22883 11104 22928 11132
rect 22922 11092 22928 11104
rect 22980 11092 22986 11144
rect 23109 11135 23167 11141
rect 23109 11101 23121 11135
rect 23155 11132 23167 11135
rect 23198 11132 23204 11144
rect 23155 11104 23204 11132
rect 23155 11101 23167 11104
rect 23109 11095 23167 11101
rect 23198 11092 23204 11104
rect 23256 11092 23262 11144
rect 23474 11092 23480 11144
rect 23532 11132 23538 11144
rect 23661 11135 23719 11141
rect 23661 11132 23673 11135
rect 23532 11104 23673 11132
rect 23532 11092 23538 11104
rect 23661 11101 23673 11104
rect 23707 11101 23719 11135
rect 23661 11095 23719 11101
rect 24026 11092 24032 11144
rect 24084 11132 24090 11144
rect 25501 11135 25559 11141
rect 25501 11132 25513 11135
rect 24084 11104 25513 11132
rect 24084 11092 24090 11104
rect 25501 11101 25513 11104
rect 25547 11101 25559 11135
rect 25501 11095 25559 11101
rect 18932 11036 19564 11064
rect 18932 11024 18938 11036
rect 21818 11024 21824 11076
rect 21876 11064 21882 11076
rect 22940 11064 22968 11092
rect 24394 11064 24400 11076
rect 21876 11036 22968 11064
rect 24044 11036 24400 11064
rect 21876 11024 21882 11036
rect 24044 11008 24072 11036
rect 24394 11024 24400 11036
rect 24452 11024 24458 11076
rect 14093 10999 14151 11005
rect 14093 10965 14105 10999
rect 14139 10996 14151 10999
rect 14182 10996 14188 11008
rect 14139 10968 14188 10996
rect 14139 10965 14151 10968
rect 14093 10959 14151 10965
rect 14182 10956 14188 10968
rect 14240 10956 14246 11008
rect 18414 10996 18420 11008
rect 18375 10968 18420 10996
rect 18414 10956 18420 10968
rect 18472 10956 18478 11008
rect 19794 10956 19800 11008
rect 19852 10996 19858 11008
rect 20073 10999 20131 11005
rect 20073 10996 20085 10999
rect 19852 10968 20085 10996
rect 19852 10956 19858 10968
rect 20073 10965 20085 10968
rect 20119 10996 20131 10999
rect 20622 10996 20628 11008
rect 20119 10968 20628 10996
rect 20119 10965 20131 10968
rect 20073 10959 20131 10965
rect 20622 10956 20628 10968
rect 20680 10956 20686 11008
rect 23106 10956 23112 11008
rect 23164 10996 23170 11008
rect 23474 10996 23480 11008
rect 23164 10968 23480 10996
rect 23164 10956 23170 10968
rect 23474 10956 23480 10968
rect 23532 10956 23538 11008
rect 24026 10956 24032 11008
rect 24084 10956 24090 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1578 10792 1584 10804
rect 1539 10764 1584 10792
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 2501 10795 2559 10801
rect 2501 10761 2513 10795
rect 2547 10792 2559 10795
rect 4246 10792 4252 10804
rect 2547 10764 4252 10792
rect 2547 10761 2559 10764
rect 2501 10755 2559 10761
rect 2608 10665 2636 10764
rect 4246 10752 4252 10764
rect 4304 10792 4310 10804
rect 4525 10795 4583 10801
rect 4525 10792 4537 10795
rect 4304 10764 4537 10792
rect 4304 10752 4310 10764
rect 4525 10761 4537 10764
rect 4571 10761 4583 10795
rect 4982 10792 4988 10804
rect 4943 10764 4988 10792
rect 4525 10755 4583 10761
rect 4982 10752 4988 10764
rect 5040 10752 5046 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 6181 10795 6239 10801
rect 6181 10792 6193 10795
rect 5592 10764 6193 10792
rect 5592 10752 5598 10764
rect 6181 10761 6193 10764
rect 6227 10761 6239 10795
rect 6181 10755 6239 10761
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10792 6699 10795
rect 6822 10792 6828 10804
rect 6687 10764 6828 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 6822 10752 6828 10764
rect 6880 10792 6886 10804
rect 7282 10792 7288 10804
rect 6880 10764 7144 10792
rect 7243 10764 7288 10792
rect 6880 10752 6886 10764
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10625 2651 10659
rect 5000 10656 5028 10752
rect 5166 10724 5172 10736
rect 5127 10696 5172 10724
rect 5166 10684 5172 10696
rect 5224 10684 5230 10736
rect 5350 10684 5356 10736
rect 5408 10724 5414 10736
rect 7006 10724 7012 10736
rect 5408 10696 7012 10724
rect 5408 10684 5414 10696
rect 7006 10684 7012 10696
rect 7064 10684 7070 10736
rect 5629 10659 5687 10665
rect 5629 10656 5641 10659
rect 5000 10628 5641 10656
rect 2593 10619 2651 10625
rect 5629 10625 5641 10628
rect 5675 10625 5687 10659
rect 5810 10656 5816 10668
rect 5771 10628 5816 10656
rect 5629 10619 5687 10625
rect 5810 10616 5816 10628
rect 5868 10616 5874 10668
rect 7116 10656 7144 10764
rect 7282 10752 7288 10764
rect 7340 10752 7346 10804
rect 10410 10792 10416 10804
rect 10371 10764 10416 10792
rect 10410 10752 10416 10764
rect 10468 10752 10474 10804
rect 11606 10792 11612 10804
rect 11567 10764 11612 10792
rect 11606 10752 11612 10764
rect 11664 10752 11670 10804
rect 11882 10792 11888 10804
rect 11843 10764 11888 10792
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 12986 10792 12992 10804
rect 12947 10764 12992 10792
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 13449 10795 13507 10801
rect 13449 10761 13461 10795
rect 13495 10792 13507 10795
rect 13538 10792 13544 10804
rect 13495 10764 13544 10792
rect 13495 10761 13507 10764
rect 13449 10755 13507 10761
rect 13538 10752 13544 10764
rect 13596 10752 13602 10804
rect 18966 10752 18972 10804
rect 19024 10792 19030 10804
rect 19061 10795 19119 10801
rect 19061 10792 19073 10795
rect 19024 10764 19073 10792
rect 19024 10752 19030 10764
rect 19061 10761 19073 10764
rect 19107 10761 19119 10795
rect 19426 10792 19432 10804
rect 19387 10764 19432 10792
rect 19061 10755 19119 10761
rect 19426 10752 19432 10764
rect 19484 10752 19490 10804
rect 19613 10795 19671 10801
rect 19613 10761 19625 10795
rect 19659 10792 19671 10795
rect 20162 10792 20168 10804
rect 19659 10764 20168 10792
rect 19659 10761 19671 10764
rect 19613 10755 19671 10761
rect 20162 10752 20168 10764
rect 20220 10752 20226 10804
rect 22094 10792 22100 10804
rect 20272 10764 22100 10792
rect 8941 10727 8999 10733
rect 8941 10693 8953 10727
rect 8987 10724 8999 10727
rect 8987 10696 11008 10724
rect 8987 10693 8999 10696
rect 8941 10687 8999 10693
rect 10980 10668 11008 10696
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7116 10628 7849 10656
rect 7837 10625 7849 10628
rect 7883 10656 7895 10659
rect 8018 10656 8024 10668
rect 7883 10628 8024 10656
rect 7883 10625 7895 10628
rect 7837 10619 7895 10625
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 9030 10616 9036 10668
rect 9088 10656 9094 10668
rect 9585 10659 9643 10665
rect 9585 10656 9597 10659
rect 9088 10628 9597 10656
rect 9088 10616 9094 10628
rect 9585 10625 9597 10628
rect 9631 10625 9643 10659
rect 10962 10656 10968 10668
rect 10923 10628 10968 10656
rect 9585 10619 9643 10625
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10557 1455 10591
rect 2860 10591 2918 10597
rect 2860 10588 2872 10591
rect 1397 10551 1455 10557
rect 2792 10560 2872 10588
rect 1412 10520 1440 10551
rect 2792 10532 2820 10560
rect 2860 10557 2872 10560
rect 2906 10588 2918 10591
rect 3786 10588 3792 10600
rect 2906 10560 3792 10588
rect 2906 10557 2918 10560
rect 2860 10551 2918 10557
rect 3786 10548 3792 10560
rect 3844 10548 3850 10600
rect 4706 10548 4712 10600
rect 4764 10588 4770 10600
rect 5537 10591 5595 10597
rect 5537 10588 5549 10591
rect 4764 10560 5549 10588
rect 4764 10548 4770 10560
rect 5537 10557 5549 10560
rect 5583 10557 5595 10591
rect 5537 10551 5595 10557
rect 7193 10591 7251 10597
rect 7193 10557 7205 10591
rect 7239 10588 7251 10591
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 7239 10560 7757 10588
rect 7239 10557 7251 10560
rect 7193 10551 7251 10557
rect 7745 10557 7757 10560
rect 7791 10588 7803 10591
rect 7926 10588 7932 10600
rect 7791 10560 7932 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 9600 10588 9628 10619
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 11149 10659 11207 10665
rect 11149 10625 11161 10659
rect 11195 10656 11207 10659
rect 11624 10656 11652 10752
rect 17862 10684 17868 10736
rect 17920 10724 17926 10736
rect 20272 10724 20300 10764
rect 22094 10752 22100 10764
rect 22152 10752 22158 10804
rect 22465 10795 22523 10801
rect 22465 10761 22477 10795
rect 22511 10792 22523 10795
rect 22554 10792 22560 10804
rect 22511 10764 22560 10792
rect 22511 10761 22523 10764
rect 22465 10755 22523 10761
rect 22554 10752 22560 10764
rect 22612 10752 22618 10804
rect 22646 10752 22652 10804
rect 22704 10792 22710 10804
rect 23198 10792 23204 10804
rect 22704 10764 23204 10792
rect 22704 10752 22710 10764
rect 23198 10752 23204 10764
rect 23256 10792 23262 10804
rect 23293 10795 23351 10801
rect 23293 10792 23305 10795
rect 23256 10764 23305 10792
rect 23256 10752 23262 10764
rect 23293 10761 23305 10764
rect 23339 10761 23351 10795
rect 23293 10755 23351 10761
rect 23750 10752 23756 10804
rect 23808 10792 23814 10804
rect 23845 10795 23903 10801
rect 23845 10792 23857 10795
rect 23808 10764 23857 10792
rect 23808 10752 23814 10764
rect 23845 10761 23857 10764
rect 23891 10761 23903 10795
rect 24762 10792 24768 10804
rect 24723 10764 24768 10792
rect 23845 10755 23903 10761
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 25590 10792 25596 10804
rect 25551 10764 25596 10792
rect 25590 10752 25596 10764
rect 25648 10752 25654 10804
rect 17920 10696 20300 10724
rect 17920 10684 17926 10696
rect 20438 10684 20444 10736
rect 20496 10724 20502 10736
rect 24578 10724 24584 10736
rect 20496 10696 24584 10724
rect 20496 10684 20502 10696
rect 24578 10684 24584 10696
rect 24636 10684 24642 10736
rect 13814 10656 13820 10668
rect 11195 10628 11652 10656
rect 13727 10628 13820 10656
rect 11195 10625 11207 10628
rect 11149 10619 11207 10625
rect 13814 10616 13820 10628
rect 13872 10656 13878 10668
rect 13909 10659 13967 10665
rect 13909 10656 13921 10659
rect 13872 10628 13921 10656
rect 13872 10616 13878 10628
rect 13909 10625 13921 10628
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 15562 10616 15568 10668
rect 15620 10656 15626 10668
rect 16945 10659 17003 10665
rect 16945 10656 16957 10659
rect 15620 10628 16957 10656
rect 15620 10616 15626 10628
rect 16945 10625 16957 10628
rect 16991 10656 17003 10659
rect 17402 10656 17408 10668
rect 16991 10628 17408 10656
rect 16991 10625 17003 10628
rect 16945 10619 17003 10625
rect 17402 10616 17408 10628
rect 17460 10656 17466 10668
rect 18414 10656 18420 10668
rect 17460 10628 18420 10656
rect 17460 10616 17466 10628
rect 18414 10616 18420 10628
rect 18472 10656 18478 10668
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 18472 10628 18613 10656
rect 18472 10616 18478 10628
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 19886 10616 19892 10668
rect 19944 10656 19950 10668
rect 20073 10659 20131 10665
rect 20073 10656 20085 10659
rect 19944 10628 20085 10656
rect 19944 10616 19950 10628
rect 20073 10625 20085 10628
rect 20119 10656 20131 10659
rect 20162 10656 20168 10668
rect 20119 10628 20168 10656
rect 20119 10625 20131 10628
rect 20073 10619 20131 10625
rect 20162 10616 20168 10628
rect 20220 10616 20226 10668
rect 20257 10659 20315 10665
rect 20257 10625 20269 10659
rect 20303 10656 20315 10659
rect 20622 10656 20628 10668
rect 20303 10628 20628 10656
rect 20303 10625 20315 10628
rect 20257 10619 20315 10625
rect 20622 10616 20628 10628
rect 20680 10656 20686 10668
rect 21450 10656 21456 10668
rect 20680 10628 21456 10656
rect 20680 10616 20686 10628
rect 21450 10616 21456 10628
rect 21508 10616 21514 10668
rect 21542 10616 21548 10668
rect 21600 10656 21606 10668
rect 21637 10659 21695 10665
rect 21637 10656 21649 10659
rect 21600 10628 21649 10656
rect 21600 10616 21606 10628
rect 21637 10625 21649 10628
rect 21683 10625 21695 10659
rect 21637 10619 21695 10625
rect 21821 10659 21879 10665
rect 21821 10625 21833 10659
rect 21867 10656 21879 10659
rect 22002 10656 22008 10668
rect 21867 10628 22008 10656
rect 21867 10625 21879 10628
rect 21821 10619 21879 10625
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 22370 10616 22376 10668
rect 22428 10656 22434 10668
rect 22649 10659 22707 10665
rect 22649 10656 22661 10659
rect 22428 10628 22661 10656
rect 22428 10616 22434 10628
rect 22649 10625 22661 10628
rect 22695 10656 22707 10659
rect 22738 10656 22744 10668
rect 22695 10628 22744 10656
rect 22695 10625 22707 10628
rect 22649 10619 22707 10625
rect 22738 10616 22744 10628
rect 22796 10616 22802 10668
rect 10045 10591 10103 10597
rect 10045 10588 10057 10591
rect 9600 10560 10057 10588
rect 10045 10557 10057 10560
rect 10091 10588 10103 10591
rect 10870 10588 10876 10600
rect 10091 10560 10876 10588
rect 10091 10557 10103 10560
rect 10045 10551 10103 10557
rect 10870 10548 10876 10560
rect 10928 10548 10934 10600
rect 16206 10588 16212 10600
rect 16167 10560 16212 10588
rect 16206 10548 16212 10560
rect 16264 10588 16270 10600
rect 16853 10591 16911 10597
rect 16853 10588 16865 10591
rect 16264 10560 16865 10588
rect 16264 10548 16270 10560
rect 16853 10557 16865 10560
rect 16899 10588 16911 10591
rect 17770 10588 17776 10600
rect 16899 10560 17776 10588
rect 16899 10557 16911 10560
rect 16853 10551 16911 10557
rect 17770 10548 17776 10560
rect 17828 10588 17834 10600
rect 18230 10588 18236 10600
rect 17828 10560 18236 10588
rect 17828 10548 17834 10560
rect 18230 10548 18236 10560
rect 18288 10548 18294 10600
rect 21192 10560 22508 10588
rect 2038 10520 2044 10532
rect 1412 10492 2044 10520
rect 2038 10480 2044 10492
rect 2096 10480 2102 10532
rect 2774 10480 2780 10532
rect 2832 10480 2838 10532
rect 3234 10480 3240 10532
rect 3292 10520 3298 10532
rect 4798 10520 4804 10532
rect 3292 10492 4804 10520
rect 3292 10480 3298 10492
rect 4798 10480 4804 10492
rect 4856 10480 4862 10532
rect 9401 10523 9459 10529
rect 9401 10520 9413 10523
rect 8772 10492 9413 10520
rect 8772 10464 8800 10492
rect 9401 10489 9413 10492
rect 9447 10489 9459 10523
rect 12342 10520 12348 10532
rect 9401 10483 9459 10489
rect 10520 10492 12348 10520
rect 3878 10412 3884 10464
rect 3936 10452 3942 10464
rect 3973 10455 4031 10461
rect 3973 10452 3985 10455
rect 3936 10424 3985 10452
rect 3936 10412 3942 10424
rect 3973 10421 3985 10424
rect 4019 10421 4031 10455
rect 3973 10415 4031 10421
rect 5718 10412 5724 10464
rect 5776 10452 5782 10464
rect 6362 10452 6368 10464
rect 5776 10424 6368 10452
rect 5776 10412 5782 10424
rect 6362 10412 6368 10424
rect 6420 10412 6426 10464
rect 7282 10412 7288 10464
rect 7340 10452 7346 10464
rect 7653 10455 7711 10461
rect 7653 10452 7665 10455
rect 7340 10424 7665 10452
rect 7340 10412 7346 10424
rect 7653 10421 7665 10424
rect 7699 10421 7711 10455
rect 7653 10415 7711 10421
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 8389 10455 8447 10461
rect 8389 10452 8401 10455
rect 8260 10424 8401 10452
rect 8260 10412 8266 10424
rect 8389 10421 8401 10424
rect 8435 10452 8447 10455
rect 8478 10452 8484 10464
rect 8435 10424 8484 10452
rect 8435 10421 8447 10424
rect 8389 10415 8447 10421
rect 8478 10412 8484 10424
rect 8536 10412 8542 10464
rect 8754 10452 8760 10464
rect 8715 10424 8760 10452
rect 8754 10412 8760 10424
rect 8812 10412 8818 10464
rect 9309 10455 9367 10461
rect 9309 10421 9321 10455
rect 9355 10452 9367 10455
rect 9582 10452 9588 10464
rect 9355 10424 9588 10452
rect 9355 10421 9367 10424
rect 9309 10415 9367 10421
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 10520 10461 10548 10492
rect 12342 10480 12348 10492
rect 12400 10480 12406 10532
rect 14182 10529 14188 10532
rect 14176 10520 14188 10529
rect 14143 10492 14188 10520
rect 14176 10483 14188 10492
rect 14182 10480 14188 10483
rect 14240 10480 14246 10532
rect 15933 10523 15991 10529
rect 15933 10489 15945 10523
rect 15979 10520 15991 10523
rect 16758 10520 16764 10532
rect 15979 10492 16764 10520
rect 15979 10489 15991 10492
rect 15933 10483 15991 10489
rect 16758 10480 16764 10492
rect 16816 10480 16822 10532
rect 17865 10523 17923 10529
rect 17865 10489 17877 10523
rect 17911 10520 17923 10523
rect 18138 10520 18144 10532
rect 17911 10492 18144 10520
rect 17911 10489 17923 10492
rect 17865 10483 17923 10489
rect 18138 10480 18144 10492
rect 18196 10520 18202 10532
rect 18509 10523 18567 10529
rect 18509 10520 18521 10523
rect 18196 10492 18521 10520
rect 18196 10480 18202 10492
rect 18509 10489 18521 10492
rect 18555 10489 18567 10523
rect 18509 10483 18567 10489
rect 18782 10480 18788 10532
rect 18840 10520 18846 10532
rect 20898 10520 20904 10532
rect 18840 10492 20904 10520
rect 18840 10480 18846 10492
rect 20898 10480 20904 10492
rect 20956 10480 20962 10532
rect 20993 10523 21051 10529
rect 20993 10489 21005 10523
rect 21039 10520 21051 10523
rect 21082 10520 21088 10532
rect 21039 10492 21088 10520
rect 21039 10489 21051 10492
rect 20993 10483 21051 10489
rect 21082 10480 21088 10492
rect 21140 10480 21146 10532
rect 10505 10455 10563 10461
rect 10505 10421 10517 10455
rect 10551 10421 10563 10455
rect 10870 10452 10876 10464
rect 10831 10424 10876 10452
rect 10505 10415 10563 10421
rect 10870 10412 10876 10424
rect 10928 10412 10934 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12492 10424 12537 10452
rect 12492 10412 12498 10424
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 15289 10455 15347 10461
rect 15289 10452 15301 10455
rect 14792 10424 15301 10452
rect 14792 10412 14798 10424
rect 15289 10421 15301 10424
rect 15335 10452 15347 10455
rect 15562 10452 15568 10464
rect 15335 10424 15568 10452
rect 15335 10421 15347 10424
rect 15289 10415 15347 10421
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 16298 10412 16304 10464
rect 16356 10452 16362 10464
rect 16393 10455 16451 10461
rect 16393 10452 16405 10455
rect 16356 10424 16405 10452
rect 16356 10412 16362 10424
rect 16393 10421 16405 10424
rect 16439 10421 16451 10455
rect 18046 10452 18052 10464
rect 18007 10424 18052 10452
rect 16393 10415 16451 10421
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 18230 10412 18236 10464
rect 18288 10452 18294 10464
rect 18414 10452 18420 10464
rect 18288 10424 18420 10452
rect 18288 10412 18294 10424
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 19242 10412 19248 10464
rect 19300 10452 19306 10464
rect 19426 10452 19432 10464
rect 19300 10424 19432 10452
rect 19300 10412 19306 10424
rect 19426 10412 19432 10424
rect 19484 10412 19490 10464
rect 19978 10452 19984 10464
rect 19939 10424 19984 10452
rect 19978 10412 19984 10424
rect 20036 10412 20042 10464
rect 21192 10461 21220 10560
rect 21545 10523 21603 10529
rect 21545 10489 21557 10523
rect 21591 10520 21603 10523
rect 21634 10520 21640 10532
rect 21591 10492 21640 10520
rect 21591 10489 21603 10492
rect 21545 10483 21603 10489
rect 21634 10480 21640 10492
rect 21692 10520 21698 10532
rect 22189 10523 22247 10529
rect 22189 10520 22201 10523
rect 21692 10492 22201 10520
rect 21692 10480 21698 10492
rect 22189 10489 22201 10492
rect 22235 10489 22247 10523
rect 22480 10520 22508 10560
rect 22554 10548 22560 10600
rect 22612 10588 22618 10600
rect 22922 10588 22928 10600
rect 22612 10560 22928 10588
rect 22612 10548 22618 10560
rect 22922 10548 22928 10560
rect 22980 10548 22986 10600
rect 24581 10591 24639 10597
rect 24581 10557 24593 10591
rect 24627 10588 24639 10591
rect 24762 10588 24768 10600
rect 24627 10560 24768 10588
rect 24627 10557 24639 10560
rect 24581 10551 24639 10557
rect 24762 10548 24768 10560
rect 24820 10588 24826 10600
rect 25133 10591 25191 10597
rect 25133 10588 25145 10591
rect 24820 10560 25145 10588
rect 24820 10548 24826 10560
rect 25133 10557 25145 10560
rect 25179 10557 25191 10591
rect 25133 10551 25191 10557
rect 24026 10520 24032 10532
rect 22480 10492 24032 10520
rect 22189 10483 22247 10489
rect 24026 10480 24032 10492
rect 24084 10480 24090 10532
rect 21177 10455 21235 10461
rect 21177 10421 21189 10455
rect 21223 10421 21235 10455
rect 21177 10415 21235 10421
rect 22278 10412 22284 10464
rect 22336 10452 22342 10464
rect 22465 10455 22523 10461
rect 22465 10452 22477 10455
rect 22336 10424 22477 10452
rect 22336 10412 22342 10424
rect 22465 10421 22477 10424
rect 22511 10421 22523 10455
rect 22465 10415 22523 10421
rect 23842 10412 23848 10464
rect 23900 10452 23906 10464
rect 24210 10452 24216 10464
rect 23900 10424 24216 10452
rect 23900 10412 23906 10424
rect 24210 10412 24216 10424
rect 24268 10452 24274 10464
rect 24397 10455 24455 10461
rect 24397 10452 24409 10455
rect 24268 10424 24409 10452
rect 24268 10412 24274 10424
rect 24397 10421 24409 10424
rect 24443 10421 24455 10455
rect 24397 10415 24455 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1854 10248 1860 10260
rect 1815 10220 1860 10248
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 2317 10251 2375 10257
rect 2317 10217 2329 10251
rect 2363 10248 2375 10251
rect 2682 10248 2688 10260
rect 2363 10220 2688 10248
rect 2363 10217 2375 10220
rect 2317 10211 2375 10217
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 2866 10248 2872 10260
rect 2823 10220 2872 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 2866 10208 2872 10220
rect 2924 10248 2930 10260
rect 3326 10248 3332 10260
rect 2924 10220 3332 10248
rect 2924 10208 2930 10220
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 4706 10208 4712 10260
rect 4764 10248 4770 10260
rect 5169 10251 5227 10257
rect 5169 10248 5181 10251
rect 4764 10220 5181 10248
rect 4764 10208 4770 10220
rect 5169 10217 5181 10220
rect 5215 10217 5227 10251
rect 5902 10248 5908 10260
rect 5863 10220 5908 10248
rect 5169 10211 5227 10217
rect 5902 10208 5908 10220
rect 5960 10208 5966 10260
rect 6454 10248 6460 10260
rect 6415 10220 6460 10248
rect 6454 10208 6460 10220
rect 6512 10208 6518 10260
rect 9401 10251 9459 10257
rect 9401 10217 9413 10251
rect 9447 10248 9459 10251
rect 9490 10248 9496 10260
rect 9447 10220 9496 10248
rect 9447 10217 9459 10220
rect 9401 10211 9459 10217
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 9861 10251 9919 10257
rect 9861 10248 9873 10251
rect 9732 10220 9873 10248
rect 9732 10208 9738 10220
rect 9861 10217 9873 10220
rect 9907 10217 9919 10251
rect 9861 10211 9919 10217
rect 10321 10251 10379 10257
rect 10321 10217 10333 10251
rect 10367 10248 10379 10251
rect 10870 10248 10876 10260
rect 10367 10220 10876 10248
rect 10367 10217 10379 10220
rect 10321 10211 10379 10217
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 11146 10208 11152 10260
rect 11204 10248 11210 10260
rect 11701 10251 11759 10257
rect 11701 10248 11713 10251
rect 11204 10220 11713 10248
rect 11204 10208 11210 10220
rect 11701 10217 11713 10220
rect 11747 10217 11759 10251
rect 11701 10211 11759 10217
rect 11885 10251 11943 10257
rect 11885 10217 11897 10251
rect 11931 10248 11943 10251
rect 11974 10248 11980 10260
rect 11931 10220 11980 10248
rect 11931 10217 11943 10220
rect 11885 10211 11943 10217
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 13446 10248 13452 10260
rect 13407 10220 13452 10248
rect 13446 10208 13452 10220
rect 13504 10208 13510 10260
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14829 10251 14887 10257
rect 14829 10248 14841 10251
rect 13872 10220 14841 10248
rect 13872 10208 13878 10220
rect 14829 10217 14841 10220
rect 14875 10217 14887 10251
rect 14829 10211 14887 10217
rect 15289 10251 15347 10257
rect 15289 10217 15301 10251
rect 15335 10248 15347 10251
rect 15378 10248 15384 10260
rect 15335 10220 15384 10248
rect 15335 10217 15347 10220
rect 15289 10211 15347 10217
rect 15378 10208 15384 10220
rect 15436 10208 15442 10260
rect 15746 10248 15752 10260
rect 15707 10220 15752 10248
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 16390 10208 16396 10260
rect 16448 10248 16454 10260
rect 16485 10251 16543 10257
rect 16485 10248 16497 10251
rect 16448 10220 16497 10248
rect 16448 10208 16454 10220
rect 16485 10217 16497 10220
rect 16531 10248 16543 10251
rect 16574 10248 16580 10260
rect 16531 10220 16580 10248
rect 16531 10217 16543 10220
rect 16485 10211 16543 10217
rect 16574 10208 16580 10220
rect 16632 10208 16638 10260
rect 19426 10208 19432 10260
rect 19484 10248 19490 10260
rect 19978 10248 19984 10260
rect 19484 10220 19984 10248
rect 19484 10208 19490 10220
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 20806 10208 20812 10260
rect 20864 10248 20870 10260
rect 20901 10251 20959 10257
rect 20901 10248 20913 10251
rect 20864 10220 20913 10248
rect 20864 10208 20870 10220
rect 20901 10217 20913 10220
rect 20947 10217 20959 10251
rect 20901 10211 20959 10217
rect 21266 10208 21272 10260
rect 21324 10208 21330 10260
rect 21542 10208 21548 10260
rect 21600 10248 21606 10260
rect 21913 10251 21971 10257
rect 21913 10248 21925 10251
rect 21600 10220 21925 10248
rect 21600 10208 21606 10220
rect 21913 10217 21925 10220
rect 21959 10217 21971 10251
rect 21913 10211 21971 10217
rect 22002 10208 22008 10260
rect 22060 10248 22066 10260
rect 22281 10251 22339 10257
rect 22281 10248 22293 10251
rect 22060 10220 22293 10248
rect 22060 10208 22066 10220
rect 22281 10217 22293 10220
rect 22327 10217 22339 10251
rect 22462 10248 22468 10260
rect 22423 10220 22468 10248
rect 22281 10211 22339 10217
rect 22462 10208 22468 10220
rect 22520 10208 22526 10260
rect 23750 10248 23756 10260
rect 23711 10220 23756 10248
rect 23750 10208 23756 10220
rect 23808 10208 23814 10260
rect 24026 10208 24032 10260
rect 24084 10248 24090 10260
rect 24397 10251 24455 10257
rect 24397 10248 24409 10251
rect 24084 10220 24409 10248
rect 24084 10208 24090 10220
rect 24397 10217 24409 10220
rect 24443 10217 24455 10251
rect 24762 10248 24768 10260
rect 24723 10220 24768 10248
rect 24397 10211 24455 10217
rect 24762 10208 24768 10220
rect 24820 10208 24826 10260
rect 25038 10248 25044 10260
rect 24999 10220 25044 10248
rect 25038 10208 25044 10220
rect 25096 10208 25102 10260
rect 25774 10248 25780 10260
rect 25735 10220 25780 10248
rect 25774 10208 25780 10220
rect 25832 10208 25838 10260
rect 3142 10140 3148 10192
rect 3200 10180 3206 10192
rect 3421 10183 3479 10189
rect 3421 10180 3433 10183
rect 3200 10152 3433 10180
rect 3200 10140 3206 10152
rect 3421 10149 3433 10152
rect 3467 10180 3479 10183
rect 3789 10183 3847 10189
rect 3789 10180 3801 10183
rect 3467 10152 3801 10180
rect 3467 10149 3479 10152
rect 3421 10143 3479 10149
rect 3789 10149 3801 10152
rect 3835 10180 3847 10183
rect 4433 10183 4491 10189
rect 3835 10152 4200 10180
rect 3835 10149 3847 10152
rect 3789 10143 3847 10149
rect 2682 10072 2688 10124
rect 2740 10112 2746 10124
rect 2869 10115 2927 10121
rect 2869 10112 2881 10115
rect 2740 10084 2881 10112
rect 2740 10072 2746 10084
rect 2869 10081 2881 10084
rect 2915 10112 2927 10115
rect 2915 10084 4108 10112
rect 2915 10081 2927 10084
rect 2869 10075 2927 10081
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 3142 10044 3148 10056
rect 3099 10016 3148 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 2958 9936 2964 9988
rect 3016 9976 3022 9988
rect 3326 9976 3332 9988
rect 3016 9948 3332 9976
rect 3016 9936 3022 9948
rect 3326 9936 3332 9948
rect 3384 9936 3390 9988
rect 4080 9976 4108 10084
rect 4172 10044 4200 10152
rect 4433 10149 4445 10183
rect 4479 10180 4491 10183
rect 5074 10180 5080 10192
rect 4479 10152 5080 10180
rect 4479 10149 4491 10152
rect 4433 10143 4491 10149
rect 5074 10140 5080 10152
rect 5132 10140 5138 10192
rect 5534 10140 5540 10192
rect 5592 10180 5598 10192
rect 10781 10183 10839 10189
rect 10781 10180 10793 10183
rect 5592 10152 10793 10180
rect 5592 10140 5598 10152
rect 10781 10149 10793 10152
rect 10827 10180 10839 10183
rect 11054 10180 11060 10192
rect 10827 10152 11060 10180
rect 10827 10149 10839 10152
rect 10781 10143 10839 10149
rect 11054 10140 11060 10152
rect 11112 10140 11118 10192
rect 12345 10183 12403 10189
rect 12345 10149 12357 10183
rect 12391 10180 12403 10183
rect 12894 10180 12900 10192
rect 12391 10152 12900 10180
rect 12391 10149 12403 10152
rect 12345 10143 12403 10149
rect 12894 10140 12900 10152
rect 12952 10140 12958 10192
rect 13722 10140 13728 10192
rect 13780 10180 13786 10192
rect 13909 10183 13967 10189
rect 13909 10180 13921 10183
rect 13780 10152 13921 10180
rect 13780 10140 13786 10152
rect 13909 10149 13921 10152
rect 13955 10149 13967 10183
rect 13909 10143 13967 10149
rect 17954 10140 17960 10192
rect 18012 10180 18018 10192
rect 19705 10183 19763 10189
rect 18012 10152 18920 10180
rect 18012 10140 18018 10152
rect 4525 10115 4583 10121
rect 4525 10081 4537 10115
rect 4571 10112 4583 10115
rect 4706 10112 4712 10124
rect 4571 10084 4712 10112
rect 4571 10081 4583 10084
rect 4525 10075 4583 10081
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10112 5687 10115
rect 5810 10112 5816 10124
rect 5675 10084 5816 10112
rect 5675 10081 5687 10084
rect 5629 10075 5687 10081
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 7926 10072 7932 10124
rect 7984 10112 7990 10124
rect 8021 10115 8079 10121
rect 8021 10112 8033 10115
rect 7984 10084 8033 10112
rect 7984 10072 7990 10084
rect 8021 10081 8033 10084
rect 8067 10081 8079 10115
rect 8021 10075 8079 10081
rect 9214 10072 9220 10124
rect 9272 10112 9278 10124
rect 10318 10112 10324 10124
rect 9272 10084 10324 10112
rect 9272 10072 9278 10084
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 10594 10072 10600 10124
rect 10652 10112 10658 10124
rect 10689 10115 10747 10121
rect 10689 10112 10701 10115
rect 10652 10084 10701 10112
rect 10652 10072 10658 10084
rect 10689 10081 10701 10084
rect 10735 10081 10747 10115
rect 10689 10075 10747 10081
rect 12253 10115 12311 10121
rect 12253 10081 12265 10115
rect 12299 10081 12311 10115
rect 12253 10075 12311 10081
rect 4617 10047 4675 10053
rect 4617 10044 4629 10047
rect 4172 10016 4629 10044
rect 4617 10013 4629 10016
rect 4663 10013 4675 10047
rect 4617 10007 4675 10013
rect 6362 10004 6368 10056
rect 6420 10044 6426 10056
rect 6549 10047 6607 10053
rect 6549 10044 6561 10047
rect 6420 10016 6561 10044
rect 6420 10004 6426 10016
rect 6549 10013 6561 10016
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10013 6699 10047
rect 6641 10007 6699 10013
rect 4338 9976 4344 9988
rect 4080 9948 4344 9976
rect 4338 9936 4344 9948
rect 4396 9936 4402 9988
rect 5718 9936 5724 9988
rect 5776 9976 5782 9988
rect 6089 9979 6147 9985
rect 6089 9976 6101 9979
rect 5776 9948 6101 9976
rect 5776 9936 5782 9948
rect 6089 9945 6101 9948
rect 6135 9945 6147 9979
rect 6089 9939 6147 9945
rect 6270 9936 6276 9988
rect 6328 9976 6334 9988
rect 6656 9976 6684 10007
rect 7374 10004 7380 10056
rect 7432 10044 7438 10056
rect 8113 10047 8171 10053
rect 8113 10044 8125 10047
rect 7432 10016 8125 10044
rect 7432 10004 7438 10016
rect 8113 10013 8125 10016
rect 8159 10013 8171 10047
rect 8113 10007 8171 10013
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10044 8263 10047
rect 8570 10044 8576 10056
rect 8251 10016 8576 10044
rect 8251 10013 8263 10016
rect 8205 10007 8263 10013
rect 7650 9976 7656 9988
rect 6328 9948 6684 9976
rect 7611 9948 7656 9976
rect 6328 9936 6334 9948
rect 7650 9936 7656 9948
rect 7708 9936 7714 9988
rect 8018 9936 8024 9988
rect 8076 9976 8082 9988
rect 8220 9976 8248 10007
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 10962 10044 10968 10056
rect 10923 10016 10968 10044
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 12268 10044 12296 10075
rect 12986 10072 12992 10124
rect 13044 10112 13050 10124
rect 13814 10112 13820 10124
rect 13044 10084 13308 10112
rect 13775 10084 13820 10112
rect 13044 10072 13050 10084
rect 12342 10044 12348 10056
rect 12268 10016 12348 10044
rect 12342 10004 12348 10016
rect 12400 10004 12406 10056
rect 12526 10044 12532 10056
rect 12487 10016 12532 10044
rect 12526 10004 12532 10016
rect 12584 10044 12590 10056
rect 13170 10044 13176 10056
rect 12584 10016 13176 10044
rect 12584 10004 12590 10016
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 13280 10044 13308 10084
rect 13814 10072 13820 10084
rect 13872 10112 13878 10124
rect 14461 10115 14519 10121
rect 14461 10112 14473 10115
rect 13872 10084 14473 10112
rect 13872 10072 13878 10084
rect 14461 10081 14473 10084
rect 14507 10081 14519 10115
rect 14461 10075 14519 10081
rect 15657 10115 15715 10121
rect 15657 10081 15669 10115
rect 15703 10112 15715 10115
rect 16850 10112 16856 10124
rect 15703 10084 16856 10112
rect 15703 10081 15715 10084
rect 15657 10075 15715 10081
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 17218 10112 17224 10124
rect 17179 10084 17224 10112
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 18782 10112 18788 10124
rect 18743 10084 18788 10112
rect 18782 10072 18788 10084
rect 18840 10072 18846 10124
rect 18892 10121 18920 10152
rect 19705 10149 19717 10183
rect 19751 10180 19763 10183
rect 20162 10180 20168 10192
rect 19751 10152 20168 10180
rect 19751 10149 19763 10152
rect 19705 10143 19763 10149
rect 20162 10140 20168 10152
rect 20220 10140 20226 10192
rect 20717 10183 20775 10189
rect 20717 10149 20729 10183
rect 20763 10180 20775 10183
rect 21284 10180 21312 10208
rect 22922 10180 22928 10192
rect 20763 10152 21312 10180
rect 22883 10152 22928 10180
rect 20763 10149 20775 10152
rect 20717 10143 20775 10149
rect 22922 10140 22928 10152
rect 22980 10140 22986 10192
rect 24210 10140 24216 10192
rect 24268 10180 24274 10192
rect 24946 10180 24952 10192
rect 24268 10152 24952 10180
rect 24268 10140 24274 10152
rect 24946 10140 24952 10152
rect 25004 10140 25010 10192
rect 18877 10115 18935 10121
rect 18877 10081 18889 10115
rect 18923 10112 18935 10115
rect 18923 10084 19104 10112
rect 18923 10081 18935 10084
rect 18877 10075 18935 10081
rect 19076 10056 19104 10084
rect 20438 10072 20444 10124
rect 20496 10112 20502 10124
rect 21269 10115 21327 10121
rect 21269 10112 21281 10115
rect 20496 10084 21281 10112
rect 20496 10072 20502 10084
rect 21269 10081 21281 10084
rect 21315 10112 21327 10115
rect 22278 10112 22284 10124
rect 21315 10084 22284 10112
rect 21315 10081 21327 10084
rect 21269 10075 21327 10081
rect 22278 10072 22284 10084
rect 22336 10072 22342 10124
rect 23569 10115 23627 10121
rect 23569 10081 23581 10115
rect 23615 10112 23627 10115
rect 23658 10112 23664 10124
rect 23615 10084 23664 10112
rect 23615 10081 23627 10084
rect 23569 10075 23627 10081
rect 23658 10072 23664 10084
rect 23716 10072 23722 10124
rect 24578 10112 24584 10124
rect 24539 10084 24584 10112
rect 24578 10072 24584 10084
rect 24636 10112 24642 10124
rect 24762 10112 24768 10124
rect 24636 10084 24768 10112
rect 24636 10072 24642 10084
rect 24762 10072 24768 10084
rect 24820 10072 24826 10124
rect 14001 10047 14059 10053
rect 14001 10044 14013 10047
rect 13280 10016 14013 10044
rect 14001 10013 14013 10016
rect 14047 10013 14059 10047
rect 15930 10044 15936 10056
rect 15891 10016 15936 10044
rect 14001 10007 14059 10013
rect 15930 10004 15936 10016
rect 15988 10004 15994 10056
rect 17310 10044 17316 10056
rect 17271 10016 17316 10044
rect 17310 10004 17316 10016
rect 17368 10004 17374 10056
rect 17402 10004 17408 10056
rect 17460 10044 17466 10056
rect 18966 10044 18972 10056
rect 17460 10016 17505 10044
rect 18927 10016 18972 10044
rect 17460 10004 17466 10016
rect 18966 10004 18972 10016
rect 19024 10004 19030 10056
rect 19058 10004 19064 10056
rect 19116 10004 19122 10056
rect 20622 10004 20628 10056
rect 20680 10044 20686 10056
rect 21361 10047 21419 10053
rect 21361 10044 21373 10047
rect 20680 10016 21373 10044
rect 20680 10004 20686 10016
rect 21361 10013 21373 10016
rect 21407 10013 21419 10047
rect 21361 10007 21419 10013
rect 21450 10004 21456 10056
rect 21508 10044 21514 10056
rect 21545 10047 21603 10053
rect 21545 10044 21557 10047
rect 21508 10016 21557 10044
rect 21508 10004 21514 10016
rect 21545 10013 21557 10016
rect 21591 10044 21603 10047
rect 22646 10044 22652 10056
rect 21591 10016 22652 10044
rect 21591 10013 21603 10016
rect 21545 10007 21603 10013
rect 22646 10004 22652 10016
rect 22704 10004 22710 10056
rect 23290 10044 23296 10056
rect 23251 10016 23296 10044
rect 23290 10004 23296 10016
rect 23348 10004 23354 10056
rect 9490 9976 9496 9988
rect 8076 9948 8248 9976
rect 8956 9948 9496 9976
rect 8076 9936 8082 9948
rect 2409 9911 2467 9917
rect 2409 9877 2421 9911
rect 2455 9908 2467 9911
rect 2590 9908 2596 9920
rect 2455 9880 2596 9908
rect 2455 9877 2467 9880
rect 2409 9871 2467 9877
rect 2590 9868 2596 9880
rect 2648 9868 2654 9920
rect 4062 9908 4068 9920
rect 4023 9880 4068 9908
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 7282 9868 7288 9920
rect 7340 9908 7346 9920
rect 7377 9911 7435 9917
rect 7377 9908 7389 9911
rect 7340 9880 7389 9908
rect 7340 9868 7346 9880
rect 7377 9877 7389 9880
rect 7423 9908 7435 9911
rect 7558 9908 7564 9920
rect 7423 9880 7564 9908
rect 7423 9877 7435 9880
rect 7377 9871 7435 9877
rect 7558 9868 7564 9880
rect 7616 9868 7622 9920
rect 8202 9868 8208 9920
rect 8260 9908 8266 9920
rect 8956 9908 8984 9948
rect 9490 9936 9496 9948
rect 9548 9936 9554 9988
rect 11330 9976 11336 9988
rect 11291 9948 11336 9976
rect 11330 9936 11336 9948
rect 11388 9936 11394 9988
rect 13081 9979 13139 9985
rect 13081 9945 13093 9979
rect 13127 9976 13139 9979
rect 14182 9976 14188 9988
rect 13127 9948 14188 9976
rect 13127 9945 13139 9948
rect 13081 9939 13139 9945
rect 14182 9936 14188 9948
rect 14240 9936 14246 9988
rect 18874 9936 18880 9988
rect 18932 9976 18938 9988
rect 21634 9976 21640 9988
rect 18932 9948 21640 9976
rect 18932 9936 18938 9948
rect 21634 9936 21640 9948
rect 21692 9936 21698 9988
rect 23198 9936 23204 9988
rect 23256 9976 23262 9988
rect 25409 9979 25467 9985
rect 25409 9976 25421 9979
rect 23256 9948 25421 9976
rect 23256 9936 23262 9948
rect 25409 9945 25421 9948
rect 25455 9945 25467 9979
rect 25409 9939 25467 9945
rect 8260 9880 8984 9908
rect 9033 9911 9091 9917
rect 8260 9868 8266 9880
rect 9033 9877 9045 9911
rect 9079 9908 9091 9911
rect 9582 9908 9588 9920
rect 9079 9880 9588 9908
rect 9079 9877 9091 9880
rect 9033 9871 9091 9877
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 10318 9868 10324 9920
rect 10376 9908 10382 9920
rect 12250 9908 12256 9920
rect 10376 9880 12256 9908
rect 10376 9868 10382 9880
rect 12250 9868 12256 9880
rect 12308 9868 12314 9920
rect 16850 9908 16856 9920
rect 16811 9880 16856 9908
rect 16850 9868 16856 9880
rect 16908 9868 16914 9920
rect 17954 9868 17960 9920
rect 18012 9908 18018 9920
rect 18049 9911 18107 9917
rect 18049 9908 18061 9911
rect 18012 9880 18061 9908
rect 18012 9868 18018 9880
rect 18049 9877 18061 9880
rect 18095 9908 18107 9911
rect 18230 9908 18236 9920
rect 18095 9880 18236 9908
rect 18095 9877 18107 9880
rect 18049 9871 18107 9877
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 18414 9908 18420 9920
rect 18375 9880 18420 9908
rect 18414 9868 18420 9880
rect 18472 9868 18478 9920
rect 24026 9908 24032 9920
rect 23987 9880 24032 9908
rect 24026 9868 24032 9880
rect 24084 9868 24090 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2866 9704 2872 9716
rect 2827 9676 2872 9704
rect 2866 9664 2872 9676
rect 2924 9664 2930 9716
rect 3050 9704 3056 9716
rect 2963 9676 3056 9704
rect 1762 9636 1768 9648
rect 1723 9608 1768 9636
rect 1762 9596 1768 9608
rect 1820 9596 1826 9648
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9568 2467 9571
rect 2774 9568 2780 9580
rect 2455 9540 2780 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 2774 9528 2780 9540
rect 2832 9568 2838 9580
rect 2976 9568 3004 9676
rect 3050 9664 3056 9676
rect 3108 9704 3114 9716
rect 3108 9676 4292 9704
rect 3108 9664 3114 9676
rect 4264 9636 4292 9676
rect 5074 9664 5080 9716
rect 5132 9704 5138 9716
rect 5261 9707 5319 9713
rect 5261 9704 5273 9707
rect 5132 9676 5273 9704
rect 5132 9664 5138 9676
rect 5261 9673 5273 9676
rect 5307 9673 5319 9707
rect 5261 9667 5319 9673
rect 5813 9707 5871 9713
rect 5813 9673 5825 9707
rect 5859 9704 5871 9707
rect 6270 9704 6276 9716
rect 5859 9676 6276 9704
rect 5859 9673 5871 9676
rect 5813 9667 5871 9673
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 6454 9704 6460 9716
rect 6415 9676 6460 9704
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 9490 9664 9496 9716
rect 9548 9704 9554 9716
rect 10597 9707 10655 9713
rect 10597 9704 10609 9707
rect 9548 9676 10609 9704
rect 9548 9664 9554 9676
rect 10597 9673 10609 9676
rect 10643 9704 10655 9707
rect 10870 9704 10876 9716
rect 10643 9676 10876 9704
rect 10643 9673 10655 9676
rect 10597 9667 10655 9673
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 11054 9704 11060 9716
rect 10980 9676 11060 9704
rect 4709 9639 4767 9645
rect 4709 9636 4721 9639
rect 4264 9608 4721 9636
rect 4709 9605 4721 9608
rect 4755 9605 4767 9639
rect 8386 9636 8392 9648
rect 4709 9599 4767 9605
rect 4816 9608 8392 9636
rect 2832 9540 3004 9568
rect 2832 9528 2838 9540
rect 4338 9528 4344 9580
rect 4396 9568 4402 9580
rect 4816 9568 4844 9608
rect 8386 9596 8392 9608
rect 8444 9596 8450 9648
rect 10980 9636 11008 9676
rect 11054 9664 11060 9676
rect 11112 9664 11118 9716
rect 11977 9707 12035 9713
rect 11977 9673 11989 9707
rect 12023 9704 12035 9707
rect 12526 9704 12532 9716
rect 12023 9676 12532 9704
rect 12023 9673 12035 9676
rect 11977 9667 12035 9673
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 14182 9704 14188 9716
rect 12768 9676 14188 9704
rect 12768 9664 12774 9676
rect 14182 9664 14188 9676
rect 14240 9704 14246 9716
rect 17770 9704 17776 9716
rect 14240 9676 17632 9704
rect 17731 9676 17776 9704
rect 14240 9664 14246 9676
rect 11149 9639 11207 9645
rect 11149 9636 11161 9639
rect 10980 9608 11161 9636
rect 11149 9605 11161 9608
rect 11195 9636 11207 9639
rect 11330 9636 11336 9648
rect 11195 9608 11336 9636
rect 11195 9605 11207 9608
rect 11149 9599 11207 9605
rect 11330 9596 11336 9608
rect 11388 9596 11394 9648
rect 11514 9636 11520 9648
rect 11475 9608 11520 9636
rect 11514 9596 11520 9608
rect 11572 9596 11578 9648
rect 12894 9636 12900 9648
rect 12855 9608 12900 9636
rect 12894 9596 12900 9608
rect 12952 9596 12958 9648
rect 14550 9596 14556 9648
rect 14608 9596 14614 9648
rect 15841 9639 15899 9645
rect 15841 9605 15853 9639
rect 15887 9636 15899 9639
rect 16022 9636 16028 9648
rect 15887 9608 16028 9636
rect 15887 9605 15899 9608
rect 15841 9599 15899 9605
rect 16022 9596 16028 9608
rect 16080 9596 16086 9648
rect 17604 9636 17632 9676
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 19058 9704 19064 9716
rect 19019 9676 19064 9704
rect 19058 9664 19064 9676
rect 19116 9664 19122 9716
rect 20438 9704 20444 9716
rect 19159 9676 20444 9704
rect 19159 9636 19187 9676
rect 20438 9664 20444 9676
rect 20496 9704 20502 9716
rect 20622 9704 20628 9716
rect 20496 9676 20628 9704
rect 20496 9664 20502 9676
rect 20622 9664 20628 9676
rect 20680 9704 20686 9716
rect 20901 9707 20959 9713
rect 20901 9704 20913 9707
rect 20680 9676 20913 9704
rect 20680 9664 20686 9676
rect 20901 9673 20913 9676
rect 20947 9673 20959 9707
rect 22278 9704 22284 9716
rect 22239 9676 22284 9704
rect 20901 9667 20959 9673
rect 22278 9664 22284 9676
rect 22336 9664 22342 9716
rect 22646 9704 22652 9716
rect 22607 9676 22652 9704
rect 22646 9664 22652 9676
rect 22704 9664 22710 9716
rect 23477 9707 23535 9713
rect 23477 9673 23489 9707
rect 23523 9704 23535 9707
rect 23658 9704 23664 9716
rect 23523 9676 23664 9704
rect 23523 9673 23535 9676
rect 23477 9667 23535 9673
rect 23658 9664 23664 9676
rect 23716 9664 23722 9716
rect 23842 9704 23848 9716
rect 23803 9676 23848 9704
rect 23842 9664 23848 9676
rect 23900 9664 23906 9716
rect 24673 9707 24731 9713
rect 24673 9673 24685 9707
rect 24719 9704 24731 9707
rect 24762 9704 24768 9716
rect 24719 9676 24768 9704
rect 24719 9673 24731 9676
rect 24673 9667 24731 9673
rect 24762 9664 24768 9676
rect 24820 9664 24826 9716
rect 17604 9608 19187 9636
rect 19613 9639 19671 9645
rect 19613 9605 19625 9639
rect 19659 9636 19671 9639
rect 20530 9636 20536 9648
rect 19659 9608 20536 9636
rect 19659 9605 19671 9608
rect 19613 9599 19671 9605
rect 20530 9596 20536 9608
rect 20588 9596 20594 9648
rect 22922 9636 22928 9648
rect 22883 9608 22928 9636
rect 22922 9596 22928 9608
rect 22980 9596 22986 9648
rect 24949 9639 25007 9645
rect 24949 9636 24961 9639
rect 23032 9608 24961 9636
rect 4396 9540 4844 9568
rect 4396 9528 4402 9540
rect 6730 9528 6736 9580
rect 6788 9528 6794 9580
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 7064 9540 7205 9568
rect 7064 9528 7070 9540
rect 7193 9537 7205 9540
rect 7239 9568 7251 9571
rect 7926 9568 7932 9580
rect 7239 9540 7932 9568
rect 7239 9537 7251 9540
rect 7193 9531 7251 9537
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 8202 9568 8208 9580
rect 8163 9540 8208 9568
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 10244 9540 13575 9568
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9500 1731 9503
rect 2682 9500 2688 9512
rect 1719 9472 2688 9500
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 3237 9503 3295 9509
rect 3237 9469 3249 9503
rect 3283 9500 3295 9503
rect 3329 9503 3387 9509
rect 3329 9500 3341 9503
rect 3283 9472 3341 9500
rect 3283 9469 3295 9472
rect 3237 9463 3295 9469
rect 3329 9469 3341 9472
rect 3375 9500 3387 9503
rect 3375 9472 4292 9500
rect 3375 9469 3387 9472
rect 3329 9463 3387 9469
rect 4264 9444 4292 9472
rect 6748 9444 6776 9528
rect 8018 9500 8024 9512
rect 7931 9472 8024 9500
rect 8018 9460 8024 9472
rect 8076 9500 8082 9512
rect 8938 9500 8944 9512
rect 8076 9472 8944 9500
rect 8076 9460 8082 9472
rect 8938 9460 8944 9472
rect 8996 9460 9002 9512
rect 9030 9460 9036 9512
rect 9088 9500 9094 9512
rect 9490 9509 9496 9512
rect 9217 9503 9275 9509
rect 9217 9500 9229 9503
rect 9088 9472 9229 9500
rect 9088 9460 9094 9472
rect 9217 9469 9229 9472
rect 9263 9469 9275 9503
rect 9484 9500 9496 9509
rect 9451 9472 9496 9500
rect 9217 9463 9275 9469
rect 9484 9463 9496 9472
rect 9490 9460 9496 9463
rect 9548 9460 9554 9512
rect 2130 9432 2136 9444
rect 2091 9404 2136 9432
rect 2130 9392 2136 9404
rect 2188 9392 2194 9444
rect 3142 9392 3148 9444
rect 3200 9432 3206 9444
rect 3574 9435 3632 9441
rect 3574 9432 3586 9435
rect 3200 9404 3586 9432
rect 3200 9392 3206 9404
rect 3574 9401 3586 9404
rect 3620 9401 3632 9435
rect 3574 9395 3632 9401
rect 4246 9392 4252 9444
rect 4304 9392 4310 9444
rect 6730 9392 6736 9444
rect 6788 9392 6794 9444
rect 7742 9392 7748 9444
rect 7800 9432 7806 9444
rect 8113 9435 8171 9441
rect 8113 9432 8125 9435
rect 7800 9404 8125 9432
rect 7800 9392 7806 9404
rect 8113 9401 8125 9404
rect 8159 9432 8171 9435
rect 8665 9435 8723 9441
rect 8665 9432 8677 9435
rect 8159 9404 8677 9432
rect 8159 9401 8171 9404
rect 8113 9395 8171 9401
rect 8665 9401 8677 9404
rect 8711 9432 8723 9435
rect 9398 9432 9404 9444
rect 8711 9404 9404 9432
rect 8711 9401 8723 9404
rect 8665 9395 8723 9401
rect 9398 9392 9404 9404
rect 9456 9392 9462 9444
rect 9674 9392 9680 9444
rect 9732 9432 9738 9444
rect 10244 9432 10272 9540
rect 13449 9503 13507 9509
rect 13449 9500 13461 9503
rect 13280 9472 13461 9500
rect 9732 9404 10272 9432
rect 9732 9392 9738 9404
rect 10318 9392 10324 9444
rect 10376 9432 10382 9444
rect 11054 9432 11060 9444
rect 10376 9404 11060 9432
rect 10376 9392 10382 9404
rect 11054 9392 11060 9404
rect 11112 9392 11118 9444
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 2225 9367 2283 9373
rect 2225 9364 2237 9367
rect 1636 9336 2237 9364
rect 1636 9324 1642 9336
rect 2225 9333 2237 9336
rect 2271 9333 2283 9367
rect 2225 9327 2283 9333
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 6089 9367 6147 9373
rect 6089 9364 6101 9367
rect 5960 9336 6101 9364
rect 5960 9324 5966 9336
rect 6089 9333 6101 9336
rect 6135 9364 6147 9367
rect 6362 9364 6368 9376
rect 6135 9336 6368 9364
rect 6135 9333 6147 9336
rect 6089 9327 6147 9333
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 7374 9324 7380 9376
rect 7432 9364 7438 9376
rect 7469 9367 7527 9373
rect 7469 9364 7481 9367
rect 7432 9336 7481 9364
rect 7432 9324 7438 9336
rect 7469 9333 7481 9336
rect 7515 9333 7527 9367
rect 7650 9364 7656 9376
rect 7611 9336 7656 9364
rect 7469 9327 7527 9333
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 9030 9364 9036 9376
rect 8991 9336 9036 9364
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 12492 9336 12537 9364
rect 12492 9324 12498 9336
rect 12986 9324 12992 9376
rect 13044 9364 13050 9376
rect 13280 9373 13308 9472
rect 13449 9469 13461 9472
rect 13495 9469 13507 9503
rect 13547 9500 13575 9540
rect 14568 9500 14596 9596
rect 15102 9528 15108 9580
rect 15160 9568 15166 9580
rect 15473 9571 15531 9577
rect 15473 9568 15485 9571
rect 15160 9540 15485 9568
rect 15160 9528 15166 9540
rect 15473 9537 15485 9540
rect 15519 9568 15531 9571
rect 15930 9568 15936 9580
rect 15519 9540 15936 9568
rect 15519 9537 15531 9540
rect 15473 9531 15531 9537
rect 15930 9528 15936 9540
rect 15988 9568 15994 9580
rect 16485 9571 16543 9577
rect 16485 9568 16497 9571
rect 15988 9540 16497 9568
rect 15988 9528 15994 9540
rect 16485 9537 16497 9540
rect 16531 9537 16543 9571
rect 18598 9568 18604 9580
rect 18559 9540 18604 9568
rect 16485 9531 16543 9537
rect 18598 9528 18604 9540
rect 18656 9568 18662 9580
rect 18966 9568 18972 9580
rect 18656 9540 18972 9568
rect 18656 9528 18662 9540
rect 18966 9528 18972 9540
rect 19024 9568 19030 9580
rect 19429 9571 19487 9577
rect 19429 9568 19441 9571
rect 19024 9540 19441 9568
rect 19024 9528 19030 9540
rect 19429 9537 19441 9540
rect 19475 9537 19487 9571
rect 20254 9568 20260 9580
rect 20215 9540 20260 9568
rect 19429 9531 19487 9537
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 20622 9528 20628 9580
rect 20680 9568 20686 9580
rect 21174 9568 21180 9580
rect 20680 9540 21180 9568
rect 20680 9528 20686 9540
rect 21174 9528 21180 9540
rect 21232 9528 21238 9580
rect 21358 9528 21364 9580
rect 21416 9568 21422 9580
rect 21729 9571 21787 9577
rect 21729 9568 21741 9571
rect 21416 9540 21741 9568
rect 21416 9528 21422 9540
rect 21729 9537 21741 9540
rect 21775 9568 21787 9571
rect 21910 9568 21916 9580
rect 21775 9540 21916 9568
rect 21775 9537 21787 9540
rect 21729 9531 21787 9537
rect 21910 9528 21916 9540
rect 21968 9528 21974 9580
rect 22373 9571 22431 9577
rect 22373 9537 22385 9571
rect 22419 9568 22431 9571
rect 23032 9568 23060 9608
rect 24949 9605 24961 9608
rect 24995 9605 25007 9639
rect 24949 9599 25007 9605
rect 22419 9540 23060 9568
rect 22419 9537 22431 9540
rect 22373 9531 22431 9537
rect 23842 9528 23848 9580
rect 23900 9568 23906 9580
rect 25317 9571 25375 9577
rect 25317 9568 25329 9571
rect 23900 9540 25329 9568
rect 23900 9528 23906 9540
rect 25317 9537 25329 9540
rect 25363 9537 25375 9571
rect 25317 9531 25375 9537
rect 16390 9500 16396 9512
rect 13547 9472 14596 9500
rect 16351 9472 16396 9500
rect 13449 9463 13507 9469
rect 16390 9460 16396 9472
rect 16448 9460 16454 9512
rect 17770 9460 17776 9512
rect 17828 9500 17834 9512
rect 18417 9503 18475 9509
rect 18417 9500 18429 9503
rect 17828 9472 18429 9500
rect 17828 9460 17834 9472
rect 18417 9469 18429 9472
rect 18463 9469 18475 9503
rect 18417 9463 18475 9469
rect 19981 9503 20039 9509
rect 19981 9469 19993 9503
rect 20027 9500 20039 9503
rect 20530 9500 20536 9512
rect 20027 9472 20536 9500
rect 20027 9469 20039 9472
rect 19981 9463 20039 9469
rect 20530 9460 20536 9472
rect 20588 9460 20594 9512
rect 20806 9460 20812 9512
rect 20864 9500 20870 9512
rect 21634 9500 21640 9512
rect 20864 9472 21640 9500
rect 20864 9460 20870 9472
rect 21634 9460 21640 9472
rect 21692 9460 21698 9512
rect 23658 9500 23664 9512
rect 22020 9472 22416 9500
rect 23619 9472 23664 9500
rect 13694 9435 13752 9441
rect 13694 9432 13706 9435
rect 13464 9404 13706 9432
rect 13464 9376 13492 9404
rect 13694 9401 13706 9404
rect 13740 9401 13752 9435
rect 13694 9395 13752 9401
rect 15746 9392 15752 9444
rect 15804 9432 15810 9444
rect 17405 9435 17463 9441
rect 17405 9432 17417 9435
rect 15804 9404 17417 9432
rect 15804 9392 15810 9404
rect 17405 9401 17417 9404
rect 17451 9432 17463 9435
rect 17954 9432 17960 9444
rect 17451 9404 17960 9432
rect 17451 9401 17463 9404
rect 17405 9395 17463 9401
rect 17954 9392 17960 9404
rect 18012 9432 18018 9444
rect 18509 9435 18567 9441
rect 18509 9432 18521 9435
rect 18012 9404 18521 9432
rect 18012 9392 18018 9404
rect 18509 9401 18521 9404
rect 18555 9401 18567 9435
rect 18509 9395 18567 9401
rect 20073 9435 20131 9441
rect 20073 9401 20085 9435
rect 20119 9432 20131 9435
rect 21542 9432 21548 9444
rect 20119 9404 21220 9432
rect 21455 9404 21548 9432
rect 20119 9401 20131 9404
rect 20073 9395 20131 9401
rect 13265 9367 13323 9373
rect 13265 9364 13277 9367
rect 13044 9336 13277 9364
rect 13044 9324 13050 9336
rect 13265 9333 13277 9336
rect 13311 9333 13323 9367
rect 13265 9327 13323 9333
rect 13446 9324 13452 9376
rect 13504 9324 13510 9376
rect 14642 9324 14648 9376
rect 14700 9364 14706 9376
rect 14829 9367 14887 9373
rect 14829 9364 14841 9367
rect 14700 9336 14841 9364
rect 14700 9324 14706 9336
rect 14829 9333 14841 9336
rect 14875 9333 14887 9367
rect 14829 9327 14887 9333
rect 15933 9367 15991 9373
rect 15933 9333 15945 9367
rect 15979 9364 15991 9367
rect 16114 9364 16120 9376
rect 15979 9336 16120 9364
rect 15979 9333 15991 9336
rect 15933 9327 15991 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 16298 9364 16304 9376
rect 16259 9336 16304 9364
rect 16298 9324 16304 9336
rect 16356 9324 16362 9376
rect 17037 9367 17095 9373
rect 17037 9333 17049 9367
rect 17083 9364 17095 9367
rect 17218 9364 17224 9376
rect 17083 9336 17224 9364
rect 17083 9333 17095 9336
rect 17037 9327 17095 9333
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 18049 9367 18107 9373
rect 18049 9333 18061 9367
rect 18095 9364 18107 9367
rect 18322 9364 18328 9376
rect 18095 9336 18328 9364
rect 18095 9333 18107 9336
rect 18049 9327 18107 9333
rect 18322 9324 18328 9336
rect 18380 9324 18386 9376
rect 18966 9324 18972 9376
rect 19024 9364 19030 9376
rect 20806 9364 20812 9376
rect 19024 9336 20812 9364
rect 19024 9324 19030 9336
rect 20806 9324 20812 9336
rect 20864 9324 20870 9376
rect 21192 9373 21220 9404
rect 21542 9392 21548 9404
rect 21600 9432 21606 9444
rect 22020 9432 22048 9472
rect 21600 9404 22048 9432
rect 22388 9432 22416 9472
rect 23658 9460 23664 9472
rect 23716 9500 23722 9512
rect 24121 9503 24179 9509
rect 24121 9500 24133 9503
rect 23716 9472 24133 9500
rect 23716 9460 23722 9472
rect 24121 9469 24133 9472
rect 24167 9469 24179 9503
rect 24121 9463 24179 9469
rect 24854 9460 24860 9512
rect 24912 9500 24918 9512
rect 25685 9503 25743 9509
rect 25685 9500 25697 9503
rect 24912 9472 25697 9500
rect 24912 9460 24918 9472
rect 25685 9469 25697 9472
rect 25731 9469 25743 9503
rect 25685 9463 25743 9469
rect 24302 9432 24308 9444
rect 22388 9404 24308 9432
rect 21600 9392 21606 9404
rect 24302 9392 24308 9404
rect 24360 9392 24366 9444
rect 21177 9367 21235 9373
rect 21177 9333 21189 9367
rect 21223 9364 21235 9367
rect 22373 9367 22431 9373
rect 22373 9364 22385 9367
rect 21223 9336 22385 9364
rect 21223 9333 21235 9336
rect 21177 9327 21235 9333
rect 22373 9333 22385 9336
rect 22419 9333 22431 9367
rect 22373 9327 22431 9333
rect 23014 9324 23020 9376
rect 23072 9364 23078 9376
rect 23382 9364 23388 9376
rect 23072 9336 23388 9364
rect 23072 9324 23078 9336
rect 23382 9324 23388 9336
rect 23440 9324 23446 9376
rect 26050 9364 26056 9376
rect 26011 9336 26056 9364
rect 26050 9324 26056 9336
rect 26108 9324 26114 9376
rect 26418 9364 26424 9376
rect 26379 9336 26424 9364
rect 26418 9324 26424 9336
rect 26476 9324 26482 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2406 9160 2412 9172
rect 2367 9132 2412 9160
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 4341 9163 4399 9169
rect 4341 9129 4353 9163
rect 4387 9160 4399 9163
rect 4706 9160 4712 9172
rect 4387 9132 4712 9160
rect 4387 9129 4399 9132
rect 4341 9123 4399 9129
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 4890 9160 4896 9172
rect 4851 9132 4896 9160
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 7926 9160 7932 9172
rect 7800 9132 7932 9160
rect 7800 9120 7806 9132
rect 7926 9120 7932 9132
rect 7984 9120 7990 9172
rect 8481 9163 8539 9169
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 8938 9160 8944 9172
rect 8527 9132 8944 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 9309 9163 9367 9169
rect 9309 9129 9321 9163
rect 9355 9160 9367 9163
rect 9490 9160 9496 9172
rect 9355 9132 9496 9160
rect 9355 9129 9367 9132
rect 9309 9123 9367 9129
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 9861 9163 9919 9169
rect 9861 9160 9873 9163
rect 9824 9132 9873 9160
rect 9824 9120 9830 9132
rect 9861 9129 9873 9132
rect 9907 9129 9919 9163
rect 9861 9123 9919 9129
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10321 9163 10379 9169
rect 10321 9160 10333 9163
rect 10192 9132 10333 9160
rect 10192 9120 10198 9132
rect 10321 9129 10333 9132
rect 10367 9129 10379 9163
rect 10321 9123 10379 9129
rect 10781 9163 10839 9169
rect 10781 9129 10793 9163
rect 10827 9160 10839 9163
rect 10962 9160 10968 9172
rect 10827 9132 10968 9160
rect 10827 9129 10839 9132
rect 10781 9123 10839 9129
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 13170 9160 13176 9172
rect 13083 9132 13176 9160
rect 13170 9120 13176 9132
rect 13228 9160 13234 9172
rect 13722 9160 13728 9172
rect 13228 9132 13728 9160
rect 13228 9120 13234 9132
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 13998 9160 14004 9172
rect 13959 9132 14004 9160
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14093 9163 14151 9169
rect 14093 9129 14105 9163
rect 14139 9160 14151 9163
rect 14918 9160 14924 9172
rect 14139 9132 14924 9160
rect 14139 9129 14151 9132
rect 14093 9123 14151 9129
rect 4798 9092 4804 9104
rect 4759 9064 4804 9092
rect 4798 9052 4804 9064
rect 4856 9052 4862 9104
rect 5810 9092 5816 9104
rect 5771 9064 5816 9092
rect 5810 9052 5816 9064
rect 5868 9052 5874 9104
rect 7006 9092 7012 9104
rect 6288 9064 7012 9092
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2222 9024 2228 9036
rect 1443 8996 2228 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2222 8984 2228 8996
rect 2280 9024 2286 9036
rect 2777 9027 2835 9033
rect 2777 9024 2789 9027
rect 2280 8996 2789 9024
rect 2280 8984 2286 8996
rect 2777 8993 2789 8996
rect 2823 8993 2835 9027
rect 2777 8987 2835 8993
rect 4246 8984 4252 9036
rect 4304 9024 4310 9036
rect 6288 9024 6316 9064
rect 7006 9052 7012 9064
rect 7064 9052 7070 9104
rect 8570 9052 8576 9104
rect 8628 9092 8634 9104
rect 8757 9095 8815 9101
rect 8757 9092 8769 9095
rect 8628 9064 8769 9092
rect 8628 9052 8634 9064
rect 8757 9061 8769 9064
rect 8803 9061 8815 9095
rect 8757 9055 8815 9061
rect 11140 9095 11198 9101
rect 11140 9061 11152 9095
rect 11186 9092 11198 9095
rect 11790 9092 11796 9104
rect 11186 9064 11796 9092
rect 11186 9061 11198 9064
rect 11140 9055 11198 9061
rect 11790 9052 11796 9064
rect 11848 9052 11854 9104
rect 13354 9052 13360 9104
rect 13412 9092 13418 9104
rect 14108 9092 14136 9123
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 15102 9160 15108 9172
rect 15063 9132 15108 9160
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 17313 9163 17371 9169
rect 17313 9129 17325 9163
rect 17359 9160 17371 9163
rect 17402 9160 17408 9172
rect 17359 9132 17408 9160
rect 17359 9129 17371 9132
rect 17313 9123 17371 9129
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 18782 9160 18788 9172
rect 18743 9132 18788 9160
rect 18782 9120 18788 9132
rect 18840 9120 18846 9172
rect 20254 9160 20260 9172
rect 20215 9132 20260 9160
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 20714 9160 20720 9172
rect 20675 9132 20720 9160
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 20898 9120 20904 9172
rect 20956 9160 20962 9172
rect 21910 9160 21916 9172
rect 20956 9132 21588 9160
rect 21871 9132 21916 9160
rect 20956 9120 20962 9132
rect 13412 9064 14136 9092
rect 13412 9052 13418 9064
rect 15286 9052 15292 9104
rect 15344 9092 15350 9104
rect 15556 9095 15614 9101
rect 15556 9092 15568 9095
rect 15344 9064 15568 9092
rect 15344 9052 15350 9064
rect 15556 9061 15568 9064
rect 15602 9092 15614 9095
rect 15838 9092 15844 9104
rect 15602 9064 15844 9092
rect 15602 9061 15614 9064
rect 15556 9055 15614 9061
rect 15838 9052 15844 9064
rect 15896 9052 15902 9104
rect 19426 9052 19432 9104
rect 19484 9092 19490 9104
rect 21358 9092 21364 9104
rect 19484 9064 21364 9092
rect 19484 9052 19490 9064
rect 21358 9052 21364 9064
rect 21416 9052 21422 9104
rect 21560 9092 21588 9132
rect 21910 9120 21916 9132
rect 21968 9120 21974 9172
rect 23290 9160 23296 9172
rect 23251 9132 23296 9160
rect 23290 9120 23296 9132
rect 23348 9120 23354 9172
rect 23474 9120 23480 9172
rect 23532 9120 23538 9172
rect 24302 9160 24308 9172
rect 24263 9132 24308 9160
rect 24302 9120 24308 9132
rect 24360 9120 24366 9172
rect 25038 9160 25044 9172
rect 24999 9132 25044 9160
rect 25038 9120 25044 9132
rect 25096 9120 25102 9172
rect 25406 9160 25412 9172
rect 25367 9132 25412 9160
rect 25406 9120 25412 9132
rect 25464 9120 25470 9172
rect 25774 9160 25780 9172
rect 25735 9132 25780 9160
rect 25774 9120 25780 9132
rect 25832 9120 25838 9172
rect 26234 9160 26240 9172
rect 26195 9132 26240 9160
rect 26234 9120 26240 9132
rect 26292 9120 26298 9172
rect 23492 9092 23520 9120
rect 24673 9095 24731 9101
rect 24673 9092 24685 9095
rect 21560 9064 22048 9092
rect 23492 9064 24685 9092
rect 4304 8996 6316 9024
rect 4304 8984 4310 8996
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 3142 8956 3148 8968
rect 3099 8928 3148 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 1949 8891 2007 8897
rect 1949 8857 1961 8891
rect 1995 8888 2007 8891
rect 2317 8891 2375 8897
rect 2317 8888 2329 8891
rect 1995 8860 2329 8888
rect 1995 8857 2007 8860
rect 1949 8851 2007 8857
rect 2317 8857 2329 8860
rect 2363 8888 2375 8891
rect 3068 8888 3096 8919
rect 3142 8916 3148 8928
rect 3200 8956 3206 8968
rect 3513 8959 3571 8965
rect 3513 8956 3525 8959
rect 3200 8928 3525 8956
rect 3200 8916 3206 8928
rect 3513 8925 3525 8928
rect 3559 8956 3571 8959
rect 3694 8956 3700 8968
rect 3559 8928 3700 8956
rect 3559 8925 3571 8928
rect 3513 8919 3571 8925
rect 3694 8916 3700 8928
rect 3752 8956 3758 8968
rect 3881 8959 3939 8965
rect 3881 8956 3893 8959
rect 3752 8928 3893 8956
rect 3752 8916 3758 8928
rect 3881 8925 3893 8928
rect 3927 8956 3939 8959
rect 5077 8959 5135 8965
rect 5077 8956 5089 8959
rect 3927 8928 5089 8956
rect 3927 8925 3939 8928
rect 3881 8919 3939 8925
rect 5077 8925 5089 8928
rect 5123 8956 5135 8959
rect 5442 8956 5448 8968
rect 5123 8928 5448 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 6288 8956 6316 8996
rect 6362 8984 6368 9036
rect 6420 9024 6426 9036
rect 6713 9027 6771 9033
rect 6713 9024 6725 9027
rect 6420 8996 6725 9024
rect 6420 8984 6426 8996
rect 6713 8993 6725 8996
rect 6759 8993 6771 9027
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 6713 8987 6771 8993
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 11974 8984 11980 9036
rect 12032 9024 12038 9036
rect 17954 9024 17960 9036
rect 12032 8996 17960 9024
rect 12032 8984 12038 8996
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 18046 8984 18052 9036
rect 18104 9024 18110 9036
rect 18141 9027 18199 9033
rect 18141 9024 18153 9027
rect 18104 8996 18153 9024
rect 18104 8984 18110 8996
rect 18141 8993 18153 8996
rect 18187 9024 18199 9027
rect 19153 9027 19211 9033
rect 19153 9024 19165 9027
rect 18187 8996 19165 9024
rect 18187 8993 18199 8996
rect 18141 8987 18199 8993
rect 19153 8993 19165 8996
rect 19199 8993 19211 9027
rect 19153 8987 19211 8993
rect 19705 9027 19763 9033
rect 19705 8993 19717 9027
rect 19751 9024 19763 9027
rect 20162 9024 20168 9036
rect 19751 8996 20168 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 20162 8984 20168 8996
rect 20220 8984 20226 9036
rect 20806 8984 20812 9036
rect 20864 9024 20870 9036
rect 21269 9027 21327 9033
rect 21269 9024 21281 9027
rect 20864 8996 21281 9024
rect 20864 8984 20870 8996
rect 21269 8993 21281 8996
rect 21315 9024 21327 9027
rect 21726 9024 21732 9036
rect 21315 8996 21732 9024
rect 21315 8993 21327 8996
rect 21269 8987 21327 8993
rect 21726 8984 21732 8996
rect 21784 8984 21790 9036
rect 6457 8959 6515 8965
rect 6457 8956 6469 8959
rect 6288 8928 6469 8956
rect 6457 8925 6469 8928
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 9030 8916 9036 8968
rect 9088 8956 9094 8968
rect 9766 8956 9772 8968
rect 9088 8928 9772 8956
rect 9088 8916 9094 8928
rect 9766 8916 9772 8928
rect 9824 8956 9830 8968
rect 10873 8959 10931 8965
rect 10873 8956 10885 8959
rect 9824 8928 10885 8956
rect 9824 8916 9830 8928
rect 10873 8925 10885 8928
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 14182 8916 14188 8968
rect 14240 8956 14246 8968
rect 14734 8956 14740 8968
rect 14240 8928 14740 8956
rect 14240 8916 14246 8928
rect 14734 8916 14740 8928
rect 14792 8916 14798 8968
rect 15289 8959 15347 8965
rect 15289 8925 15301 8959
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 2363 8860 3096 8888
rect 2363 8857 2375 8860
rect 2317 8851 2375 8857
rect 13538 8848 13544 8900
rect 13596 8888 13602 8900
rect 13633 8891 13691 8897
rect 13633 8888 13645 8891
rect 13596 8860 13645 8888
rect 13596 8848 13602 8860
rect 13633 8857 13645 8860
rect 13679 8857 13691 8891
rect 13633 8851 13691 8857
rect 4433 8823 4491 8829
rect 4433 8789 4445 8823
rect 4479 8820 4491 8823
rect 5166 8820 5172 8832
rect 4479 8792 5172 8820
rect 4479 8789 4491 8792
rect 4433 8783 4491 8789
rect 5166 8780 5172 8792
rect 5224 8780 5230 8832
rect 5534 8820 5540 8832
rect 5495 8792 5540 8820
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 6273 8823 6331 8829
rect 6273 8789 6285 8823
rect 6319 8820 6331 8823
rect 6454 8820 6460 8832
rect 6319 8792 6460 8820
rect 6319 8789 6331 8792
rect 6273 8783 6331 8789
rect 6454 8780 6460 8792
rect 6512 8780 6518 8832
rect 7837 8823 7895 8829
rect 7837 8789 7849 8823
rect 7883 8820 7895 8823
rect 7926 8820 7932 8832
rect 7883 8792 7932 8820
rect 7883 8789 7895 8792
rect 7837 8783 7895 8789
rect 7926 8780 7932 8792
rect 7984 8780 7990 8832
rect 12158 8780 12164 8832
rect 12216 8820 12222 8832
rect 12253 8823 12311 8829
rect 12253 8820 12265 8823
rect 12216 8792 12265 8820
rect 12216 8780 12222 8792
rect 12253 8789 12265 8792
rect 12299 8789 12311 8823
rect 13446 8820 13452 8832
rect 13407 8792 13452 8820
rect 12253 8783 12311 8789
rect 13446 8780 13452 8792
rect 13504 8780 13510 8832
rect 14734 8820 14740 8832
rect 14695 8792 14740 8820
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 15304 8820 15332 8919
rect 16298 8916 16304 8968
rect 16356 8956 16362 8968
rect 17218 8956 17224 8968
rect 16356 8928 17224 8956
rect 16356 8916 16362 8928
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 18230 8956 18236 8968
rect 18191 8928 18236 8956
rect 18230 8916 18236 8928
rect 18288 8916 18294 8968
rect 18325 8959 18383 8965
rect 18325 8925 18337 8959
rect 18371 8956 18383 8959
rect 18598 8956 18604 8968
rect 18371 8928 18604 8956
rect 18371 8925 18383 8928
rect 18325 8919 18383 8925
rect 16574 8848 16580 8900
rect 16632 8888 16638 8900
rect 17773 8891 17831 8897
rect 17773 8888 17785 8891
rect 16632 8860 17785 8888
rect 16632 8848 16638 8860
rect 17773 8857 17785 8860
rect 17819 8857 17831 8891
rect 18340 8888 18368 8919
rect 18598 8916 18604 8928
rect 18656 8916 18662 8968
rect 19978 8916 19984 8968
rect 20036 8956 20042 8968
rect 20622 8956 20628 8968
rect 20036 8928 20628 8956
rect 20036 8916 20042 8928
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 21358 8956 21364 8968
rect 21319 8928 21364 8956
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 21450 8916 21456 8968
rect 21508 8956 21514 8968
rect 21508 8928 21553 8956
rect 21508 8916 21514 8928
rect 19610 8888 19616 8900
rect 17773 8851 17831 8857
rect 18248 8860 18368 8888
rect 19571 8860 19616 8888
rect 15562 8820 15568 8832
rect 15304 8792 15568 8820
rect 15562 8780 15568 8792
rect 15620 8780 15626 8832
rect 16669 8823 16727 8829
rect 16669 8789 16681 8823
rect 16715 8820 16727 8823
rect 17218 8820 17224 8832
rect 16715 8792 17224 8820
rect 16715 8789 16727 8792
rect 16669 8783 16727 8789
rect 17218 8780 17224 8792
rect 17276 8780 17282 8832
rect 17402 8780 17408 8832
rect 17460 8820 17466 8832
rect 17589 8823 17647 8829
rect 17589 8820 17601 8823
rect 17460 8792 17601 8820
rect 17460 8780 17466 8792
rect 17589 8789 17601 8792
rect 17635 8820 17647 8823
rect 18248 8820 18276 8860
rect 19610 8848 19616 8860
rect 19668 8848 19674 8900
rect 20990 8848 20996 8900
rect 21048 8888 21054 8900
rect 21910 8888 21916 8900
rect 21048 8860 21916 8888
rect 21048 8848 21054 8860
rect 21910 8848 21916 8860
rect 21968 8848 21974 8900
rect 22020 8888 22048 9064
rect 24673 9061 24685 9064
rect 24719 9061 24731 9095
rect 24673 9055 24731 9061
rect 22094 8984 22100 9036
rect 22152 9024 22158 9036
rect 22465 9027 22523 9033
rect 22465 9024 22477 9027
rect 22152 8996 22477 9024
rect 22152 8984 22158 8996
rect 22465 8993 22477 8996
rect 22511 9024 22523 9027
rect 23014 9024 23020 9036
rect 22511 8996 23020 9024
rect 22511 8993 22523 8996
rect 22465 8987 22523 8993
rect 23014 8984 23020 8996
rect 23072 8984 23078 9036
rect 23477 9027 23535 9033
rect 23477 8993 23489 9027
rect 23523 9024 23535 9027
rect 23934 9024 23940 9036
rect 23523 8996 23940 9024
rect 23523 8993 23535 8996
rect 23477 8987 23535 8993
rect 23934 8984 23940 8996
rect 23992 8984 23998 9036
rect 22189 8959 22247 8965
rect 22189 8925 22201 8959
rect 22235 8956 22247 8959
rect 26050 8956 26056 8968
rect 22235 8928 26056 8956
rect 22235 8925 22247 8928
rect 22189 8919 22247 8925
rect 26050 8916 26056 8928
rect 26108 8916 26114 8968
rect 23566 8888 23572 8900
rect 22020 8860 23572 8888
rect 23566 8848 23572 8860
rect 23624 8848 23630 8900
rect 17635 8792 18276 8820
rect 19889 8823 19947 8829
rect 17635 8789 17647 8792
rect 17589 8783 17647 8789
rect 19889 8789 19901 8823
rect 19935 8820 19947 8823
rect 20622 8820 20628 8832
rect 19935 8792 20628 8820
rect 19935 8789 19947 8792
rect 19889 8783 19947 8789
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 20898 8820 20904 8832
rect 20859 8792 20904 8820
rect 20898 8780 20904 8792
rect 20956 8780 20962 8832
rect 21358 8780 21364 8832
rect 21416 8820 21422 8832
rect 22097 8823 22155 8829
rect 22097 8820 22109 8823
rect 21416 8792 22109 8820
rect 21416 8780 21422 8792
rect 22097 8789 22109 8792
rect 22143 8789 22155 8823
rect 22278 8820 22284 8832
rect 22239 8792 22284 8820
rect 22097 8783 22155 8789
rect 22278 8780 22284 8792
rect 22336 8780 22342 8832
rect 22646 8820 22652 8832
rect 22607 8792 22652 8820
rect 22646 8780 22652 8792
rect 22704 8780 22710 8832
rect 22922 8820 22928 8832
rect 22883 8792 22928 8820
rect 22922 8780 22928 8792
rect 22980 8780 22986 8832
rect 23658 8820 23664 8832
rect 23619 8792 23664 8820
rect 23658 8780 23664 8792
rect 23716 8780 23722 8832
rect 23934 8820 23940 8832
rect 23895 8792 23940 8820
rect 23934 8780 23940 8792
rect 23992 8780 23998 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1489 8619 1547 8625
rect 1489 8585 1501 8619
rect 1535 8616 1547 8619
rect 2038 8616 2044 8628
rect 1535 8588 2044 8616
rect 1535 8585 1547 8588
rect 1489 8579 1547 8585
rect 2038 8576 2044 8588
rect 2096 8616 2102 8628
rect 2314 8616 2320 8628
rect 2096 8588 2320 8616
rect 2096 8576 2102 8588
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 4890 8616 4896 8628
rect 4203 8588 4896 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 5721 8619 5779 8625
rect 5721 8585 5733 8619
rect 5767 8616 5779 8619
rect 5997 8619 6055 8625
rect 5997 8616 6009 8619
rect 5767 8588 6009 8616
rect 5767 8585 5779 8588
rect 5721 8579 5779 8585
rect 5997 8585 6009 8588
rect 6043 8585 6055 8619
rect 5997 8579 6055 8585
rect 9125 8619 9183 8625
rect 9125 8585 9137 8619
rect 9171 8616 9183 8619
rect 9490 8616 9496 8628
rect 9171 8588 9496 8616
rect 9171 8585 9183 8588
rect 9125 8579 9183 8585
rect 2593 8551 2651 8557
rect 2593 8517 2605 8551
rect 2639 8548 2651 8551
rect 2866 8548 2872 8560
rect 2639 8520 2872 8548
rect 2639 8517 2651 8520
rect 2593 8511 2651 8517
rect 2866 8508 2872 8520
rect 2924 8548 2930 8560
rect 4617 8551 4675 8557
rect 2924 8520 3832 8548
rect 2924 8508 2930 8520
rect 1762 8440 1768 8492
rect 1820 8480 1826 8492
rect 1949 8483 2007 8489
rect 1949 8480 1961 8483
rect 1820 8452 1961 8480
rect 1820 8440 1826 8452
rect 1949 8449 1961 8452
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8449 2099 8483
rect 3694 8480 3700 8492
rect 3655 8452 3700 8480
rect 2041 8443 2099 8449
rect 1854 8412 1860 8424
rect 1815 8384 1860 8412
rect 1854 8372 1860 8384
rect 1912 8372 1918 8424
rect 2056 8276 2084 8443
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8412 3019 8415
rect 3326 8412 3332 8424
rect 3007 8384 3332 8412
rect 3007 8381 3019 8384
rect 2961 8375 3019 8381
rect 3326 8372 3332 8384
rect 3384 8412 3390 8424
rect 3421 8415 3479 8421
rect 3421 8412 3433 8415
rect 3384 8384 3433 8412
rect 3384 8372 3390 8384
rect 3421 8381 3433 8384
rect 3467 8381 3479 8415
rect 3421 8375 3479 8381
rect 3513 8415 3571 8421
rect 3513 8381 3525 8415
rect 3559 8412 3571 8415
rect 3559 8384 3740 8412
rect 3559 8381 3571 8384
rect 3513 8375 3571 8381
rect 3712 8356 3740 8384
rect 2884 8316 3188 8344
rect 2884 8276 2912 8316
rect 2056 8248 2912 8276
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 3053 8279 3111 8285
rect 3053 8276 3065 8279
rect 3016 8248 3065 8276
rect 3016 8236 3022 8248
rect 3053 8245 3065 8248
rect 3099 8245 3111 8279
rect 3160 8276 3188 8316
rect 3694 8304 3700 8356
rect 3752 8304 3758 8356
rect 3804 8344 3832 8520
rect 4617 8517 4629 8551
rect 4663 8548 4675 8551
rect 5258 8548 5264 8560
rect 4663 8520 5264 8548
rect 4663 8517 4675 8520
rect 4617 8511 4675 8517
rect 5258 8508 5264 8520
rect 5316 8508 5322 8560
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 4798 8480 4804 8492
rect 4571 8452 4804 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5442 8480 5448 8492
rect 5215 8452 5448 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 5442 8440 5448 8452
rect 5500 8480 5506 8492
rect 5736 8480 5764 8579
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 10042 8576 10048 8628
rect 10100 8616 10106 8628
rect 10229 8619 10287 8625
rect 10229 8616 10241 8619
rect 10100 8588 10241 8616
rect 10100 8576 10106 8588
rect 10229 8585 10241 8588
rect 10275 8585 10287 8619
rect 12066 8616 12072 8628
rect 12027 8588 12072 8616
rect 10229 8579 10287 8585
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 14645 8619 14703 8625
rect 14645 8616 14657 8619
rect 14516 8588 14657 8616
rect 14516 8576 14522 8588
rect 14645 8585 14657 8588
rect 14691 8585 14703 8619
rect 15746 8616 15752 8628
rect 15707 8588 15752 8616
rect 14645 8579 14703 8585
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 20073 8619 20131 8625
rect 20073 8585 20085 8619
rect 20119 8616 20131 8619
rect 20162 8616 20168 8628
rect 20119 8588 20168 8616
rect 20119 8585 20131 8588
rect 20073 8579 20131 8585
rect 20162 8576 20168 8588
rect 20220 8576 20226 8628
rect 20530 8616 20536 8628
rect 20491 8588 20536 8616
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 21450 8576 21456 8628
rect 21508 8616 21514 8628
rect 21545 8619 21603 8625
rect 21545 8616 21557 8619
rect 21508 8588 21557 8616
rect 21508 8576 21514 8588
rect 21545 8585 21557 8588
rect 21591 8585 21603 8619
rect 22741 8619 22799 8625
rect 22741 8616 22753 8619
rect 21545 8579 21603 8585
rect 22112 8588 22753 8616
rect 12084 8548 12112 8576
rect 10704 8520 12112 8548
rect 5500 8452 5764 8480
rect 5500 8440 5506 8452
rect 7006 8440 7012 8492
rect 7064 8440 7070 8492
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 10594 8480 10600 8492
rect 10100 8452 10600 8480
rect 10100 8440 10106 8452
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 10704 8489 10732 8520
rect 16022 8508 16028 8560
rect 16080 8548 16086 8560
rect 16080 8520 16344 8548
rect 16080 8508 16086 8520
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8480 10931 8483
rect 10962 8480 10968 8492
rect 10919 8452 10968 8480
rect 10919 8449 10931 8452
rect 10873 8443 10931 8449
rect 4706 8372 4712 8424
rect 4764 8412 4770 8424
rect 4985 8415 5043 8421
rect 4985 8412 4997 8415
rect 4764 8384 4997 8412
rect 4764 8372 4770 8384
rect 4985 8381 4997 8384
rect 5031 8412 5043 8415
rect 6178 8412 6184 8424
rect 5031 8384 6184 8412
rect 5031 8381 5043 8384
rect 4985 8375 5043 8381
rect 6178 8372 6184 8384
rect 6236 8372 6242 8424
rect 6549 8415 6607 8421
rect 6549 8412 6561 8415
rect 6288 8384 6561 8412
rect 5626 8344 5632 8356
rect 3804 8316 5632 8344
rect 5626 8304 5632 8316
rect 5684 8304 5690 8356
rect 3878 8276 3884 8288
rect 3160 8248 3884 8276
rect 3053 8239 3111 8245
rect 3878 8236 3884 8248
rect 3936 8236 3942 8288
rect 4982 8236 4988 8288
rect 5040 8276 5046 8288
rect 5077 8279 5135 8285
rect 5077 8276 5089 8279
rect 5040 8248 5089 8276
rect 5040 8236 5046 8248
rect 5077 8245 5089 8248
rect 5123 8245 5135 8279
rect 5077 8239 5135 8245
rect 6178 8236 6184 8288
rect 6236 8276 6242 8288
rect 6288 8276 6316 8384
rect 6549 8381 6561 8384
rect 6595 8412 6607 8415
rect 7024 8412 7052 8440
rect 7653 8415 7711 8421
rect 7653 8412 7665 8415
rect 6595 8384 7665 8412
rect 6595 8381 6607 8384
rect 6549 8375 6607 8381
rect 7653 8381 7665 8384
rect 7699 8412 7711 8415
rect 7745 8415 7803 8421
rect 7745 8412 7757 8415
rect 7699 8384 7757 8412
rect 7699 8381 7711 8384
rect 7653 8375 7711 8381
rect 7745 8381 7757 8384
rect 7791 8412 7803 8415
rect 9030 8412 9036 8424
rect 7791 8384 9036 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 9030 8372 9036 8384
rect 9088 8372 9094 8424
rect 9769 8415 9827 8421
rect 9769 8381 9781 8415
rect 9815 8412 9827 8415
rect 10888 8412 10916 8443
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 12986 8440 12992 8492
rect 13044 8480 13050 8492
rect 13081 8483 13139 8489
rect 13081 8480 13093 8483
rect 13044 8452 13093 8480
rect 13044 8440 13050 8452
rect 13081 8449 13093 8452
rect 13127 8480 13139 8483
rect 13265 8483 13323 8489
rect 13265 8480 13277 8483
rect 13127 8452 13277 8480
rect 13127 8449 13139 8452
rect 13081 8443 13139 8449
rect 13265 8449 13277 8452
rect 13311 8449 13323 8483
rect 13265 8443 13323 8449
rect 15657 8483 15715 8489
rect 15657 8449 15669 8483
rect 15703 8480 15715 8483
rect 16206 8480 16212 8492
rect 15703 8452 16212 8480
rect 15703 8449 15715 8452
rect 15657 8443 15715 8449
rect 16206 8440 16212 8452
rect 16264 8440 16270 8492
rect 16316 8489 16344 8520
rect 19058 8508 19064 8560
rect 19116 8548 19122 8560
rect 19429 8551 19487 8557
rect 19429 8548 19441 8551
rect 19116 8520 19441 8548
rect 19116 8508 19122 8520
rect 19429 8517 19441 8520
rect 19475 8548 19487 8551
rect 20441 8551 20499 8557
rect 20441 8548 20453 8551
rect 19475 8520 20453 8548
rect 19475 8517 19487 8520
rect 19429 8511 19487 8517
rect 20441 8517 20453 8520
rect 20487 8548 20499 8551
rect 20487 8520 21128 8548
rect 20487 8517 20499 8520
rect 20441 8511 20499 8517
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8449 16359 8483
rect 20990 8480 20996 8492
rect 20951 8452 20996 8480
rect 16301 8443 16359 8449
rect 20990 8440 20996 8452
rect 21048 8440 21054 8492
rect 21100 8489 21128 8520
rect 21085 8483 21143 8489
rect 21085 8449 21097 8483
rect 21131 8449 21143 8483
rect 21085 8443 21143 8449
rect 15838 8412 15844 8424
rect 9815 8384 10916 8412
rect 10980 8384 15844 8412
rect 9815 8381 9827 8384
rect 9769 8375 9827 8381
rect 7926 8304 7932 8356
rect 7984 8353 7990 8356
rect 7984 8347 8048 8353
rect 7984 8313 8002 8347
rect 8036 8313 8048 8347
rect 7984 8307 8048 8313
rect 10137 8347 10195 8353
rect 10137 8313 10149 8347
rect 10183 8344 10195 8347
rect 10597 8347 10655 8353
rect 10597 8344 10609 8347
rect 10183 8316 10609 8344
rect 10183 8313 10195 8316
rect 10137 8307 10195 8313
rect 10597 8313 10609 8316
rect 10643 8344 10655 8347
rect 10778 8344 10784 8356
rect 10643 8316 10784 8344
rect 10643 8313 10655 8316
rect 10597 8307 10655 8313
rect 7984 8304 7990 8307
rect 10778 8304 10784 8316
rect 10836 8344 10842 8356
rect 10980 8344 11008 8384
rect 15838 8372 15844 8384
rect 15896 8372 15902 8424
rect 16666 8372 16672 8424
rect 16724 8412 16730 8424
rect 17773 8415 17831 8421
rect 17773 8412 17785 8415
rect 16724 8384 17785 8412
rect 16724 8372 16730 8384
rect 10836 8316 11008 8344
rect 12805 8347 12863 8353
rect 10836 8304 10842 8316
rect 12805 8313 12817 8347
rect 12851 8344 12863 8347
rect 13532 8347 13590 8353
rect 13532 8344 13544 8347
rect 12851 8316 13544 8344
rect 12851 8313 12863 8316
rect 12805 8307 12863 8313
rect 13532 8313 13544 8316
rect 13578 8344 13590 8347
rect 13630 8344 13636 8356
rect 13578 8316 13636 8344
rect 13578 8313 13590 8316
rect 13532 8307 13590 8313
rect 13630 8304 13636 8316
rect 13688 8304 13694 8356
rect 15197 8347 15255 8353
rect 15197 8344 15209 8347
rect 14936 8316 15209 8344
rect 7006 8276 7012 8288
rect 6236 8248 6316 8276
rect 6967 8248 7012 8276
rect 6236 8236 6242 8248
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 9766 8236 9772 8288
rect 9824 8276 9830 8288
rect 11333 8279 11391 8285
rect 11333 8276 11345 8279
rect 9824 8248 11345 8276
rect 9824 8236 9830 8248
rect 11333 8245 11345 8248
rect 11379 8276 11391 8279
rect 11514 8276 11520 8288
rect 11379 8248 11520 8276
rect 11379 8245 11391 8248
rect 11333 8239 11391 8245
rect 11514 8236 11520 8248
rect 11572 8236 11578 8288
rect 11701 8279 11759 8285
rect 11701 8245 11713 8279
rect 11747 8276 11759 8279
rect 11790 8276 11796 8288
rect 11747 8248 11796 8276
rect 11747 8245 11759 8248
rect 11701 8239 11759 8245
rect 11790 8236 11796 8248
rect 11848 8236 11854 8288
rect 12434 8236 12440 8288
rect 12492 8276 12498 8288
rect 14936 8276 14964 8316
rect 15197 8313 15209 8316
rect 15243 8344 15255 8347
rect 15470 8344 15476 8356
rect 15243 8316 15476 8344
rect 15243 8313 15255 8316
rect 15197 8307 15255 8313
rect 15470 8304 15476 8316
rect 15528 8344 15534 8356
rect 16117 8347 16175 8353
rect 16117 8344 16129 8347
rect 15528 8316 16129 8344
rect 15528 8304 15534 8316
rect 16117 8313 16129 8316
rect 16163 8313 16175 8347
rect 16117 8307 16175 8313
rect 12492 8248 14964 8276
rect 12492 8236 12498 8248
rect 15286 8236 15292 8288
rect 15344 8276 15350 8288
rect 15562 8276 15568 8288
rect 15344 8248 15568 8276
rect 15344 8236 15350 8248
rect 15562 8236 15568 8248
rect 15620 8276 15626 8288
rect 16776 8285 16804 8384
rect 17773 8381 17785 8384
rect 17819 8412 17831 8415
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 17819 8384 18061 8412
rect 17819 8381 17831 8384
rect 17773 8375 17831 8381
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 20714 8372 20720 8424
rect 20772 8412 20778 8424
rect 20901 8415 20959 8421
rect 20901 8412 20913 8415
rect 20772 8384 20913 8412
rect 20772 8372 20778 8384
rect 20901 8381 20913 8384
rect 20947 8381 20959 8415
rect 21726 8412 21732 8424
rect 20901 8375 20959 8381
rect 21468 8384 21732 8412
rect 18294 8347 18352 8353
rect 18294 8344 18306 8347
rect 17420 8316 18306 8344
rect 17420 8288 17448 8316
rect 18294 8313 18306 8316
rect 18340 8313 18352 8347
rect 18294 8307 18352 8313
rect 20438 8304 20444 8356
rect 20496 8344 20502 8356
rect 21468 8344 21496 8384
rect 21726 8372 21732 8384
rect 21784 8372 21790 8424
rect 22112 8421 22140 8588
rect 22741 8585 22753 8588
rect 22787 8616 22799 8619
rect 22830 8616 22836 8628
rect 22787 8588 22836 8616
rect 22787 8585 22799 8588
rect 22741 8579 22799 8585
rect 22830 8576 22836 8588
rect 22888 8576 22894 8628
rect 23014 8616 23020 8628
rect 22975 8588 23020 8616
rect 23014 8576 23020 8588
rect 23072 8576 23078 8628
rect 23474 8616 23480 8628
rect 23435 8588 23480 8616
rect 23474 8576 23480 8588
rect 23532 8576 23538 8628
rect 24026 8576 24032 8628
rect 24084 8616 24090 8628
rect 24121 8619 24179 8625
rect 24121 8616 24133 8619
rect 24084 8588 24133 8616
rect 24084 8576 24090 8588
rect 24121 8585 24133 8588
rect 24167 8585 24179 8619
rect 24121 8579 24179 8585
rect 25130 8576 25136 8628
rect 25188 8616 25194 8628
rect 25225 8619 25283 8625
rect 25225 8616 25237 8619
rect 25188 8588 25237 8616
rect 25188 8576 25194 8588
rect 25225 8585 25237 8588
rect 25271 8585 25283 8619
rect 25682 8616 25688 8628
rect 25643 8588 25688 8616
rect 25225 8579 25283 8585
rect 25682 8576 25688 8588
rect 25740 8576 25746 8628
rect 25958 8616 25964 8628
rect 25919 8588 25964 8616
rect 25958 8576 25964 8588
rect 26016 8576 26022 8628
rect 26326 8616 26332 8628
rect 26287 8588 26332 8616
rect 26326 8576 26332 8588
rect 26384 8576 26390 8628
rect 22281 8551 22339 8557
rect 22281 8517 22293 8551
rect 22327 8548 22339 8551
rect 23198 8548 23204 8560
rect 22327 8520 23204 8548
rect 22327 8517 22339 8520
rect 22281 8511 22339 8517
rect 23198 8508 23204 8520
rect 23256 8508 23262 8560
rect 24949 8551 25007 8557
rect 24949 8517 24961 8551
rect 24995 8548 25007 8551
rect 26142 8548 26148 8560
rect 24995 8520 26148 8548
rect 24995 8517 25007 8520
rect 24949 8511 25007 8517
rect 26142 8508 26148 8520
rect 26200 8508 26206 8560
rect 22186 8440 22192 8492
rect 22244 8480 22250 8492
rect 23474 8480 23480 8492
rect 22244 8452 23480 8480
rect 22244 8440 22250 8452
rect 23474 8440 23480 8452
rect 23532 8440 23538 8492
rect 22097 8415 22155 8421
rect 22097 8381 22109 8415
rect 22143 8381 22155 8415
rect 23658 8412 23664 8424
rect 23619 8384 23664 8412
rect 22097 8375 22155 8381
rect 23658 8372 23664 8384
rect 23716 8412 23722 8424
rect 24489 8415 24547 8421
rect 24489 8412 24501 8415
rect 23716 8384 24501 8412
rect 23716 8372 23722 8384
rect 24489 8381 24501 8384
rect 24535 8381 24547 8415
rect 24489 8375 24547 8381
rect 20496 8316 21496 8344
rect 21560 8316 22048 8344
rect 20496 8304 20502 8316
rect 16761 8279 16819 8285
rect 16761 8276 16773 8279
rect 15620 8248 16773 8276
rect 15620 8236 15626 8248
rect 16761 8245 16773 8248
rect 16807 8245 16819 8279
rect 17402 8276 17408 8288
rect 17363 8248 17408 8276
rect 16761 8239 16819 8245
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 21266 8236 21272 8288
rect 21324 8276 21330 8288
rect 21560 8276 21588 8316
rect 21324 8248 21588 8276
rect 21324 8236 21330 8248
rect 21634 8236 21640 8288
rect 21692 8276 21698 8288
rect 21913 8279 21971 8285
rect 21913 8276 21925 8279
rect 21692 8248 21925 8276
rect 21692 8236 21698 8248
rect 21913 8245 21925 8248
rect 21959 8245 21971 8279
rect 22020 8276 22048 8316
rect 22738 8276 22744 8288
rect 22020 8248 22744 8276
rect 21913 8239 21971 8245
rect 22738 8236 22744 8248
rect 22796 8236 22802 8288
rect 23842 8276 23848 8288
rect 23803 8248 23848 8276
rect 23842 8236 23848 8248
rect 23900 8236 23906 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 2222 8072 2228 8084
rect 2183 8044 2228 8072
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 2406 8032 2412 8084
rect 2464 8072 2470 8084
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 2464 8044 2789 8072
rect 2464 8032 2470 8044
rect 2777 8041 2789 8044
rect 2823 8041 2835 8075
rect 2777 8035 2835 8041
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 4212 8044 4261 8072
rect 4212 8032 4218 8044
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 4706 8072 4712 8084
rect 4667 8044 4712 8072
rect 4249 8035 4307 8041
rect 4706 8032 4712 8044
rect 4764 8032 4770 8084
rect 4982 8032 4988 8084
rect 5040 8072 5046 8084
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 5040 8044 5089 8072
rect 5040 8032 5046 8044
rect 5077 8041 5089 8044
rect 5123 8072 5135 8075
rect 8662 8072 8668 8084
rect 5123 8044 8668 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 10505 8075 10563 8081
rect 10505 8041 10517 8075
rect 10551 8072 10563 8075
rect 10686 8072 10692 8084
rect 10551 8044 10692 8072
rect 10551 8041 10563 8044
rect 10505 8035 10563 8041
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 11146 8032 11152 8084
rect 11204 8072 11210 8084
rect 11609 8075 11667 8081
rect 11609 8072 11621 8075
rect 11204 8044 11621 8072
rect 11204 8032 11210 8044
rect 11609 8041 11621 8044
rect 11655 8072 11667 8075
rect 12342 8072 12348 8084
rect 11655 8044 12348 8072
rect 11655 8041 11667 8044
rect 11609 8035 11667 8041
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 14093 8075 14151 8081
rect 14093 8041 14105 8075
rect 14139 8072 14151 8075
rect 14182 8072 14188 8084
rect 14139 8044 14188 8072
rect 14139 8041 14151 8044
rect 14093 8035 14151 8041
rect 14182 8032 14188 8044
rect 14240 8032 14246 8084
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 17773 8075 17831 8081
rect 17773 8041 17785 8075
rect 17819 8072 17831 8075
rect 18230 8072 18236 8084
rect 17819 8044 18236 8072
rect 17819 8041 17831 8044
rect 17773 8035 17831 8041
rect 18230 8032 18236 8044
rect 18288 8072 18294 8084
rect 19153 8075 19211 8081
rect 19153 8072 19165 8075
rect 18288 8044 19165 8072
rect 18288 8032 18294 8044
rect 19153 8041 19165 8044
rect 19199 8041 19211 8075
rect 19153 8035 19211 8041
rect 20717 8075 20775 8081
rect 20717 8041 20729 8075
rect 20763 8072 20775 8075
rect 20990 8072 20996 8084
rect 20763 8044 20996 8072
rect 20763 8041 20775 8044
rect 20717 8035 20775 8041
rect 20990 8032 20996 8044
rect 21048 8032 21054 8084
rect 22830 8032 22836 8084
rect 22888 8072 22894 8084
rect 22925 8075 22983 8081
rect 22925 8072 22937 8075
rect 22888 8044 22937 8072
rect 22888 8032 22894 8044
rect 22925 8041 22937 8044
rect 22971 8041 22983 8075
rect 22925 8035 22983 8041
rect 24118 8032 24124 8084
rect 24176 8072 24182 8084
rect 24581 8075 24639 8081
rect 24581 8072 24593 8075
rect 24176 8044 24593 8072
rect 24176 8032 24182 8044
rect 24581 8041 24593 8044
rect 24627 8041 24639 8075
rect 25038 8072 25044 8084
rect 24999 8044 25044 8072
rect 24581 8035 24639 8041
rect 25038 8032 25044 8044
rect 25096 8032 25102 8084
rect 2869 8007 2927 8013
rect 2869 7973 2881 8007
rect 2915 8004 2927 8007
rect 2958 8004 2964 8016
rect 2915 7976 2964 8004
rect 2915 7973 2927 7976
rect 2869 7967 2927 7973
rect 2958 7964 2964 7976
rect 3016 7964 3022 8016
rect 5620 8007 5678 8013
rect 5620 7973 5632 8007
rect 5666 8004 5678 8007
rect 6086 8004 6092 8016
rect 5666 7976 6092 8004
rect 5666 7973 5678 7976
rect 5620 7967 5678 7973
rect 6086 7964 6092 7976
rect 6144 7964 6150 8016
rect 8481 8007 8539 8013
rect 8481 7973 8493 8007
rect 8527 8004 8539 8007
rect 8570 8004 8576 8016
rect 8527 7976 8576 8004
rect 8527 7973 8539 7976
rect 8481 7967 8539 7973
rect 8570 7964 8576 7976
rect 8628 7964 8634 8016
rect 10045 8007 10103 8013
rect 10045 7973 10057 8007
rect 10091 8004 10103 8007
rect 10778 8004 10784 8016
rect 10091 7976 10784 8004
rect 10091 7973 10103 7976
rect 10045 7967 10103 7973
rect 10778 7964 10784 7976
rect 10836 7964 10842 8016
rect 10873 8007 10931 8013
rect 10873 7973 10885 8007
rect 10919 8004 10931 8007
rect 10962 8004 10968 8016
rect 10919 7976 10968 8004
rect 10919 7973 10931 7976
rect 10873 7967 10931 7973
rect 10962 7964 10968 7976
rect 11020 7964 11026 8016
rect 14642 7964 14648 8016
rect 14700 8004 14706 8016
rect 15534 8007 15592 8013
rect 15534 8004 15546 8007
rect 14700 7976 15546 8004
rect 14700 7964 14706 7976
rect 15534 7973 15546 7976
rect 15580 8004 15592 8007
rect 16114 8004 16120 8016
rect 15580 7976 16120 8004
rect 15580 7973 15592 7976
rect 15534 7967 15592 7973
rect 16114 7964 16120 7976
rect 16172 8004 16178 8016
rect 17589 8007 17647 8013
rect 17589 8004 17601 8007
rect 16172 7976 17601 8004
rect 16172 7964 16178 7976
rect 17589 7973 17601 7976
rect 17635 8004 17647 8007
rect 17635 7976 18368 8004
rect 17635 7973 17647 7976
rect 17589 7967 17647 7973
rect 3602 7896 3608 7948
rect 3660 7936 3666 7948
rect 4065 7939 4123 7945
rect 4065 7936 4077 7939
rect 3660 7908 4077 7936
rect 3660 7896 3666 7908
rect 4065 7905 4077 7908
rect 4111 7905 4123 7939
rect 4065 7899 4123 7905
rect 5353 7939 5411 7945
rect 5353 7905 5365 7939
rect 5399 7936 5411 7939
rect 6178 7936 6184 7948
rect 5399 7908 6184 7936
rect 5399 7905 5411 7908
rect 5353 7899 5411 7905
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7936 7527 7939
rect 8386 7936 8392 7948
rect 7515 7908 8392 7936
rect 7515 7905 7527 7908
rect 7469 7899 7527 7905
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 10796 7936 10824 7964
rect 12158 7936 12164 7948
rect 10796 7908 11100 7936
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 3050 7868 3056 7880
rect 3007 7840 3056 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 1857 7803 1915 7809
rect 1857 7769 1869 7803
rect 1903 7800 1915 7803
rect 2976 7800 3004 7831
rect 3050 7828 3056 7840
rect 3108 7828 3114 7880
rect 3513 7871 3571 7877
rect 3513 7837 3525 7871
rect 3559 7868 3571 7871
rect 3694 7868 3700 7880
rect 3559 7840 3700 7868
rect 3559 7837 3571 7840
rect 3513 7831 3571 7837
rect 3694 7828 3700 7840
rect 3752 7828 3758 7880
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7868 7895 7871
rect 7926 7868 7932 7880
rect 7883 7840 7932 7868
rect 7883 7837 7895 7840
rect 7837 7831 7895 7837
rect 7926 7828 7932 7840
rect 7984 7828 7990 7880
rect 8202 7828 8208 7880
rect 8260 7868 8266 7880
rect 8573 7871 8631 7877
rect 8573 7868 8585 7871
rect 8260 7840 8585 7868
rect 8260 7828 8266 7840
rect 8573 7837 8585 7840
rect 8619 7837 8631 7871
rect 8573 7831 8631 7837
rect 1903 7772 3004 7800
rect 8588 7800 8616 7831
rect 9766 7828 9772 7880
rect 9824 7868 9830 7880
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 9824 7840 10333 7868
rect 9824 7828 9830 7840
rect 10321 7837 10333 7840
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 10870 7828 10876 7880
rect 10928 7868 10934 7880
rect 11072 7877 11100 7908
rect 11900 7908 12164 7936
rect 10965 7871 11023 7877
rect 10965 7868 10977 7871
rect 10928 7840 10977 7868
rect 10928 7828 10934 7840
rect 10965 7837 10977 7840
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7837 11115 7871
rect 11057 7831 11115 7837
rect 11900 7809 11928 7908
rect 12158 7896 12164 7908
rect 12216 7936 12222 7948
rect 12325 7939 12383 7945
rect 12325 7936 12337 7939
rect 12216 7908 12337 7936
rect 12216 7896 12222 7908
rect 12325 7905 12337 7908
rect 12371 7905 12383 7939
rect 18141 7939 18199 7945
rect 18141 7936 18153 7939
rect 12325 7899 12383 7905
rect 18064 7908 18153 7936
rect 12069 7871 12127 7877
rect 12069 7837 12081 7871
rect 12115 7837 12127 7871
rect 15286 7868 15292 7880
rect 15247 7840 15292 7868
rect 12069 7831 12127 7837
rect 11885 7803 11943 7809
rect 11885 7800 11897 7803
rect 8588 7772 11897 7800
rect 1903 7769 1915 7772
rect 1857 7763 1915 7769
rect 11885 7769 11897 7772
rect 11931 7769 11943 7803
rect 11885 7763 11943 7769
rect 2406 7732 2412 7744
rect 2367 7704 2412 7732
rect 2406 7692 2412 7704
rect 2464 7692 2470 7744
rect 3878 7732 3884 7744
rect 3791 7704 3884 7732
rect 3878 7692 3884 7704
rect 3936 7732 3942 7744
rect 4614 7732 4620 7744
rect 3936 7704 4620 7732
rect 3936 7692 3942 7704
rect 4614 7692 4620 7704
rect 4672 7692 4678 7744
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 6362 7732 6368 7744
rect 5592 7704 6368 7732
rect 5592 7692 5598 7704
rect 6362 7692 6368 7704
rect 6420 7732 6426 7744
rect 6733 7735 6791 7741
rect 6733 7732 6745 7735
rect 6420 7704 6745 7732
rect 6420 7692 6426 7704
rect 6733 7701 6745 7704
rect 6779 7732 6791 7735
rect 7006 7732 7012 7744
rect 6779 7704 7012 7732
rect 6779 7701 6791 7704
rect 6733 7695 6791 7701
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 8018 7732 8024 7744
rect 7979 7704 8024 7732
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 9309 7735 9367 7741
rect 9309 7701 9321 7735
rect 9355 7732 9367 7735
rect 9582 7732 9588 7744
rect 9355 7704 9588 7732
rect 9355 7701 9367 7704
rect 9309 7695 9367 7701
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 11514 7692 11520 7744
rect 11572 7732 11578 7744
rect 12084 7732 12112 7831
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 18064 7800 18092 7908
rect 18141 7905 18153 7908
rect 18187 7905 18199 7939
rect 18141 7899 18199 7905
rect 18230 7868 18236 7880
rect 18191 7840 18236 7868
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 18340 7877 18368 7976
rect 18506 7964 18512 8016
rect 18564 8004 18570 8016
rect 18601 8007 18659 8013
rect 18601 8004 18613 8007
rect 18564 7976 18613 8004
rect 18564 7964 18570 7976
rect 18601 7973 18613 7976
rect 18647 7973 18659 8007
rect 18601 7967 18659 7973
rect 21910 7964 21916 8016
rect 21968 8004 21974 8016
rect 21968 7976 22784 8004
rect 21968 7964 21974 7976
rect 22756 7948 22784 7976
rect 19334 7936 19340 7948
rect 19295 7908 19340 7936
rect 19334 7896 19340 7908
rect 19392 7896 19398 7948
rect 21269 7939 21327 7945
rect 21269 7905 21281 7939
rect 21315 7936 21327 7939
rect 22370 7936 22376 7948
rect 21315 7908 22376 7936
rect 21315 7905 21327 7908
rect 21269 7899 21327 7905
rect 22370 7896 22376 7908
rect 22428 7896 22434 7948
rect 22738 7896 22744 7948
rect 22796 7936 22802 7948
rect 22833 7939 22891 7945
rect 22833 7936 22845 7939
rect 22796 7908 22845 7936
rect 22796 7896 22802 7908
rect 22833 7905 22845 7908
rect 22879 7905 22891 7939
rect 22833 7899 22891 7905
rect 23474 7896 23480 7948
rect 23532 7936 23538 7948
rect 24026 7936 24032 7948
rect 23532 7908 24032 7936
rect 23532 7896 23538 7908
rect 24026 7896 24032 7908
rect 24084 7896 24090 7948
rect 25133 7939 25191 7945
rect 25133 7905 25145 7939
rect 25179 7936 25191 7939
rect 25222 7936 25228 7948
rect 25179 7908 25228 7936
rect 25179 7905 25191 7908
rect 25133 7899 25191 7905
rect 25222 7896 25228 7908
rect 25280 7896 25286 7948
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7868 18383 7871
rect 18598 7868 18604 7880
rect 18371 7840 18604 7868
rect 18371 7837 18383 7840
rect 18325 7831 18383 7837
rect 18598 7828 18604 7840
rect 18656 7868 18662 7880
rect 18785 7871 18843 7877
rect 18785 7868 18797 7871
rect 18656 7840 18797 7868
rect 18656 7828 18662 7840
rect 18785 7837 18797 7840
rect 18831 7837 18843 7871
rect 18785 7831 18843 7837
rect 19242 7828 19248 7880
rect 19300 7868 19306 7880
rect 20257 7871 20315 7877
rect 20257 7868 20269 7871
rect 19300 7840 20269 7868
rect 19300 7828 19306 7840
rect 20257 7837 20269 7840
rect 20303 7837 20315 7871
rect 20257 7831 20315 7837
rect 21361 7871 21419 7877
rect 21361 7837 21373 7871
rect 21407 7837 21419 7871
rect 21361 7831 21419 7837
rect 21545 7871 21603 7877
rect 21545 7837 21557 7871
rect 21591 7868 21603 7871
rect 21726 7868 21732 7880
rect 21591 7840 21732 7868
rect 21591 7837 21603 7840
rect 21545 7831 21603 7837
rect 18506 7800 18512 7812
rect 18064 7772 18512 7800
rect 18506 7760 18512 7772
rect 18564 7760 18570 7812
rect 19886 7800 19892 7812
rect 19847 7772 19892 7800
rect 19886 7760 19892 7772
rect 19944 7760 19950 7812
rect 20438 7800 20444 7812
rect 20180 7772 20444 7800
rect 12986 7732 12992 7744
rect 11572 7704 12992 7732
rect 11572 7692 11578 7704
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 13446 7732 13452 7744
rect 13407 7704 13452 7732
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 14458 7732 14464 7744
rect 14419 7704 14464 7732
rect 14458 7692 14464 7704
rect 14516 7692 14522 7744
rect 16022 7692 16028 7744
rect 16080 7732 16086 7744
rect 16669 7735 16727 7741
rect 16669 7732 16681 7735
rect 16080 7704 16681 7732
rect 16080 7692 16086 7704
rect 16669 7701 16681 7704
rect 16715 7732 16727 7735
rect 17221 7735 17279 7741
rect 17221 7732 17233 7735
rect 16715 7704 17233 7732
rect 16715 7701 16727 7704
rect 16669 7695 16727 7701
rect 17221 7701 17233 7704
rect 17267 7732 17279 7735
rect 17402 7732 17408 7744
rect 17267 7704 17408 7732
rect 17267 7701 17279 7704
rect 17221 7695 17279 7701
rect 17402 7692 17408 7704
rect 17460 7692 17466 7744
rect 18230 7692 18236 7744
rect 18288 7732 18294 7744
rect 18601 7735 18659 7741
rect 18601 7732 18613 7735
rect 18288 7704 18613 7732
rect 18288 7692 18294 7704
rect 18601 7701 18613 7704
rect 18647 7701 18659 7735
rect 18601 7695 18659 7701
rect 19521 7735 19579 7741
rect 19521 7701 19533 7735
rect 19567 7732 19579 7735
rect 20180 7732 20208 7772
rect 20438 7760 20444 7772
rect 20496 7760 20502 7812
rect 21376 7800 21404 7831
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 23014 7868 23020 7880
rect 22975 7840 23020 7868
rect 23014 7828 23020 7840
rect 23072 7828 23078 7880
rect 26050 7868 26056 7880
rect 26011 7840 26056 7868
rect 26050 7828 26056 7840
rect 26108 7828 26114 7880
rect 22465 7803 22523 7809
rect 21376 7772 21956 7800
rect 21928 7744 21956 7772
rect 22465 7769 22477 7803
rect 22511 7800 22523 7803
rect 23382 7800 23388 7812
rect 22511 7772 23388 7800
rect 22511 7769 22523 7772
rect 22465 7763 22523 7769
rect 23382 7760 23388 7772
rect 23440 7760 23446 7812
rect 19567 7704 20208 7732
rect 20901 7735 20959 7741
rect 19567 7701 19579 7704
rect 19521 7695 19579 7701
rect 20901 7701 20913 7735
rect 20947 7732 20959 7735
rect 21542 7732 21548 7744
rect 20947 7704 21548 7732
rect 20947 7701 20959 7704
rect 20901 7695 20959 7701
rect 21542 7692 21548 7704
rect 21600 7692 21606 7744
rect 21910 7732 21916 7744
rect 21871 7704 21916 7732
rect 21910 7692 21916 7704
rect 21968 7692 21974 7744
rect 22370 7732 22376 7744
rect 22331 7704 22376 7732
rect 22370 7692 22376 7704
rect 22428 7692 22434 7744
rect 23474 7732 23480 7744
rect 23435 7704 23480 7732
rect 23474 7692 23480 7704
rect 23532 7692 23538 7744
rect 23566 7692 23572 7744
rect 23624 7732 23630 7744
rect 23845 7735 23903 7741
rect 23845 7732 23857 7735
rect 23624 7704 23857 7732
rect 23624 7692 23630 7704
rect 23845 7701 23857 7704
rect 23891 7701 23903 7735
rect 23845 7695 23903 7701
rect 24213 7735 24271 7741
rect 24213 7701 24225 7735
rect 24259 7732 24271 7735
rect 25130 7732 25136 7744
rect 24259 7704 25136 7732
rect 24259 7701 24271 7704
rect 24213 7695 24271 7701
rect 25130 7692 25136 7704
rect 25188 7692 25194 7744
rect 25314 7732 25320 7744
rect 25275 7704 25320 7732
rect 25314 7692 25320 7704
rect 25372 7692 25378 7744
rect 25682 7732 25688 7744
rect 25643 7704 25688 7732
rect 25682 7692 25688 7704
rect 25740 7692 25746 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 3142 7528 3148 7540
rect 3103 7500 3148 7528
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 6086 7528 6092 7540
rect 6047 7500 6092 7528
rect 6086 7488 6092 7500
rect 6144 7488 6150 7540
rect 8202 7528 8208 7540
rect 8163 7500 8208 7528
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 8386 7488 8392 7540
rect 8444 7528 8450 7540
rect 10781 7531 10839 7537
rect 10781 7528 10793 7531
rect 8444 7500 10793 7528
rect 8444 7488 8450 7500
rect 10781 7497 10793 7500
rect 10827 7497 10839 7531
rect 10781 7491 10839 7497
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 11882 7528 11888 7540
rect 10928 7500 11888 7528
rect 10928 7488 10934 7500
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 18046 7528 18052 7540
rect 18007 7500 18052 7528
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 19334 7528 19340 7540
rect 19295 7500 19340 7528
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 19613 7531 19671 7537
rect 19613 7497 19625 7531
rect 19659 7528 19671 7531
rect 20806 7528 20812 7540
rect 19659 7500 20812 7528
rect 19659 7497 19671 7500
rect 19613 7491 19671 7497
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 21174 7528 21180 7540
rect 21135 7500 21180 7528
rect 21174 7488 21180 7500
rect 21232 7488 21238 7540
rect 22922 7528 22928 7540
rect 22883 7500 22928 7528
rect 22922 7488 22928 7500
rect 22980 7488 22986 7540
rect 24026 7488 24032 7540
rect 24084 7528 24090 7540
rect 24581 7531 24639 7537
rect 24581 7528 24593 7531
rect 24084 7500 24593 7528
rect 24084 7488 24090 7500
rect 24581 7497 24593 7500
rect 24627 7497 24639 7531
rect 24581 7491 24639 7497
rect 25222 7488 25228 7540
rect 25280 7528 25286 7540
rect 25317 7531 25375 7537
rect 25317 7528 25329 7531
rect 25280 7500 25329 7528
rect 25280 7488 25286 7500
rect 25317 7497 25329 7500
rect 25363 7497 25375 7531
rect 25317 7491 25375 7497
rect 25498 7488 25504 7540
rect 25556 7528 25562 7540
rect 25685 7531 25743 7537
rect 25685 7528 25697 7531
rect 25556 7500 25697 7528
rect 25556 7488 25562 7500
rect 25685 7497 25697 7500
rect 25731 7497 25743 7531
rect 25685 7491 25743 7497
rect 2685 7463 2743 7469
rect 2685 7429 2697 7463
rect 2731 7460 2743 7463
rect 3050 7460 3056 7472
rect 2731 7432 3056 7460
rect 2731 7429 2743 7432
rect 2685 7423 2743 7429
rect 3050 7420 3056 7432
rect 3108 7460 3114 7472
rect 4525 7463 4583 7469
rect 4525 7460 4537 7463
rect 3108 7432 4537 7460
rect 3108 7420 3114 7432
rect 2038 7392 2044 7404
rect 1999 7364 2044 7392
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 2222 7392 2228 7404
rect 2135 7364 2228 7392
rect 2222 7352 2228 7364
rect 2280 7392 2286 7404
rect 3712 7401 3740 7432
rect 4525 7429 4537 7432
rect 4571 7460 4583 7463
rect 7098 7460 7104 7472
rect 4571 7432 5304 7460
rect 7059 7432 7104 7460
rect 4571 7429 4583 7432
rect 4525 7423 4583 7429
rect 3697 7395 3755 7401
rect 2280 7364 3556 7392
rect 2280 7352 2286 7364
rect 1946 7324 1952 7336
rect 1907 7296 1952 7324
rect 1946 7284 1952 7296
rect 2004 7284 2010 7336
rect 3528 7256 3556 7364
rect 3697 7361 3709 7395
rect 3743 7361 3755 7395
rect 5166 7392 5172 7404
rect 5127 7364 5172 7392
rect 3697 7355 3755 7361
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 5276 7401 5304 7432
rect 7098 7420 7104 7432
rect 7156 7420 7162 7472
rect 8570 7460 8576 7472
rect 8531 7432 8576 7460
rect 8570 7420 8576 7432
rect 8628 7420 8634 7472
rect 12434 7420 12440 7472
rect 12492 7460 12498 7472
rect 17129 7463 17187 7469
rect 12492 7432 12537 7460
rect 12492 7420 12498 7432
rect 17129 7429 17141 7463
rect 17175 7460 17187 7463
rect 17586 7460 17592 7472
rect 17175 7432 17592 7460
rect 17175 7429 17187 7432
rect 17129 7423 17187 7429
rect 17586 7420 17592 7432
rect 17644 7460 17650 7472
rect 18506 7460 18512 7472
rect 17644 7432 18512 7460
rect 17644 7420 17650 7432
rect 18506 7420 18512 7432
rect 18564 7420 18570 7472
rect 19352 7460 19380 7488
rect 19352 7432 20668 7460
rect 5261 7395 5319 7401
rect 5261 7361 5273 7395
rect 5307 7361 5319 7395
rect 5261 7355 5319 7361
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7392 6699 7395
rect 7745 7395 7803 7401
rect 7745 7392 7757 7395
rect 6687 7364 7757 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 7745 7361 7757 7364
rect 7791 7392 7803 7395
rect 7926 7392 7932 7404
rect 7791 7364 7932 7392
rect 7791 7361 7803 7364
rect 7745 7355 7803 7361
rect 7926 7352 7932 7364
rect 7984 7352 7990 7404
rect 9766 7392 9772 7404
rect 9727 7364 9772 7392
rect 9766 7352 9772 7364
rect 9824 7392 9830 7404
rect 11333 7395 11391 7401
rect 11333 7392 11345 7395
rect 9824 7364 11345 7392
rect 9824 7352 9830 7364
rect 11333 7361 11345 7364
rect 11379 7392 11391 7395
rect 11790 7392 11796 7404
rect 11379 7364 11796 7392
rect 11379 7361 11391 7364
rect 11333 7355 11391 7361
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 13538 7392 13544 7404
rect 13127 7364 13544 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 13998 7352 14004 7404
rect 14056 7392 14062 7404
rect 14553 7395 14611 7401
rect 14553 7392 14565 7395
rect 14056 7364 14565 7392
rect 14056 7352 14062 7364
rect 14553 7361 14565 7364
rect 14599 7361 14611 7395
rect 16114 7392 16120 7404
rect 16075 7364 16120 7392
rect 14553 7355 14611 7361
rect 16114 7352 16120 7364
rect 16172 7392 16178 7404
rect 16577 7395 16635 7401
rect 16577 7392 16589 7395
rect 16172 7364 16589 7392
rect 16172 7352 16178 7364
rect 16577 7361 16589 7364
rect 16623 7361 16635 7395
rect 18598 7392 18604 7404
rect 18559 7364 18604 7392
rect 16577 7355 16635 7361
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 19886 7352 19892 7404
rect 19944 7392 19950 7404
rect 20165 7395 20223 7401
rect 20165 7392 20177 7395
rect 19944 7364 20177 7392
rect 19944 7352 19950 7364
rect 20165 7361 20177 7364
rect 20211 7361 20223 7395
rect 20165 7355 20223 7361
rect 20254 7352 20260 7404
rect 20312 7352 20318 7404
rect 20640 7392 20668 7432
rect 20714 7420 20720 7472
rect 20772 7460 20778 7472
rect 21085 7463 21143 7469
rect 21085 7460 21097 7463
rect 20772 7432 21097 7460
rect 20772 7420 20778 7432
rect 21085 7429 21097 7432
rect 21131 7460 21143 7463
rect 21131 7432 21772 7460
rect 21131 7429 21143 7432
rect 21085 7423 21143 7429
rect 20898 7392 20904 7404
rect 20640 7364 20904 7392
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 21634 7392 21640 7404
rect 21595 7364 21640 7392
rect 21634 7352 21640 7364
rect 21692 7352 21698 7404
rect 21744 7401 21772 7432
rect 21729 7395 21787 7401
rect 21729 7361 21741 7395
rect 21775 7361 21787 7395
rect 21729 7355 21787 7361
rect 22554 7352 22560 7404
rect 22612 7392 22618 7404
rect 24213 7395 24271 7401
rect 24213 7392 24225 7395
rect 22612 7364 24225 7392
rect 22612 7352 22618 7364
rect 3605 7327 3663 7333
rect 3605 7293 3617 7327
rect 3651 7324 3663 7327
rect 3786 7324 3792 7336
rect 3651 7296 3792 7324
rect 3651 7293 3663 7296
rect 3605 7287 3663 7293
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 5534 7324 5540 7336
rect 3896 7296 5540 7324
rect 3896 7256 3924 7296
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 5813 7327 5871 7333
rect 5813 7293 5825 7327
rect 5859 7324 5871 7327
rect 6178 7324 6184 7336
rect 5859 7296 6184 7324
rect 5859 7293 5871 7296
rect 5813 7287 5871 7293
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 7558 7324 7564 7336
rect 7519 7296 7564 7324
rect 7558 7284 7564 7296
rect 7616 7284 7622 7336
rect 11146 7324 11152 7336
rect 11107 7296 11152 7324
rect 11146 7284 11152 7296
rect 11204 7284 11210 7336
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 14458 7324 14464 7336
rect 13872 7296 14464 7324
rect 13872 7284 13878 7296
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 15105 7327 15163 7333
rect 15105 7293 15117 7327
rect 15151 7324 15163 7327
rect 15654 7324 15660 7336
rect 15151 7296 15660 7324
rect 15151 7293 15163 7296
rect 15105 7287 15163 7293
rect 15654 7284 15660 7296
rect 15712 7324 15718 7336
rect 16025 7327 16083 7333
rect 16025 7324 16037 7327
rect 15712 7296 16037 7324
rect 15712 7284 15718 7296
rect 16025 7293 16037 7296
rect 16071 7293 16083 7327
rect 16025 7287 16083 7293
rect 19978 7284 19984 7336
rect 20036 7324 20042 7336
rect 20073 7327 20131 7333
rect 20073 7324 20085 7327
rect 20036 7296 20085 7324
rect 20036 7284 20042 7296
rect 20073 7293 20085 7296
rect 20119 7324 20131 7327
rect 20272 7324 20300 7352
rect 21542 7324 21548 7336
rect 20119 7296 20300 7324
rect 21503 7296 21548 7324
rect 20119 7293 20131 7296
rect 20073 7287 20131 7293
rect 21542 7284 21548 7296
rect 21600 7284 21606 7336
rect 23676 7333 23704 7364
rect 24213 7361 24225 7364
rect 24259 7361 24271 7395
rect 24213 7355 24271 7361
rect 23661 7327 23719 7333
rect 23661 7293 23673 7327
rect 23707 7293 23719 7327
rect 23661 7287 23719 7293
rect 23842 7284 23848 7336
rect 23900 7324 23906 7336
rect 24762 7324 24768 7336
rect 23900 7296 24768 7324
rect 23900 7284 23906 7296
rect 24762 7284 24768 7296
rect 24820 7284 24826 7336
rect 3528 7228 3924 7256
rect 5077 7259 5135 7265
rect 5077 7225 5089 7259
rect 5123 7256 5135 7259
rect 5258 7256 5264 7268
rect 5123 7228 5264 7256
rect 5123 7225 5135 7228
rect 5077 7219 5135 7225
rect 5258 7216 5264 7228
rect 5316 7216 5322 7268
rect 7374 7216 7380 7268
rect 7432 7256 7438 7268
rect 7469 7259 7527 7265
rect 7469 7256 7481 7259
rect 7432 7228 7481 7256
rect 7432 7216 7438 7228
rect 7469 7225 7481 7228
rect 7515 7225 7527 7259
rect 7469 7219 7527 7225
rect 9125 7259 9183 7265
rect 9125 7225 9137 7259
rect 9171 7256 9183 7259
rect 9582 7256 9588 7268
rect 9171 7228 9588 7256
rect 9171 7225 9183 7228
rect 9125 7219 9183 7225
rect 9582 7216 9588 7228
rect 9640 7216 9646 7268
rect 10321 7259 10379 7265
rect 10321 7225 10333 7259
rect 10367 7256 10379 7259
rect 10962 7256 10968 7268
rect 10367 7228 10968 7256
rect 10367 7225 10379 7228
rect 10321 7219 10379 7225
rect 10962 7216 10968 7228
rect 11020 7216 11026 7268
rect 11054 7216 11060 7268
rect 11112 7256 11118 7268
rect 12253 7259 12311 7265
rect 12253 7256 12265 7259
rect 11112 7228 12265 7256
rect 11112 7216 11118 7228
rect 12253 7225 12265 7228
rect 12299 7256 12311 7259
rect 12805 7259 12863 7265
rect 12805 7256 12817 7259
rect 12299 7228 12817 7256
rect 12299 7225 12311 7228
rect 12253 7219 12311 7225
rect 12805 7225 12817 7228
rect 12851 7225 12863 7259
rect 12805 7219 12863 7225
rect 15473 7259 15531 7265
rect 15473 7225 15485 7259
rect 15519 7256 15531 7259
rect 15746 7256 15752 7268
rect 15519 7228 15752 7256
rect 15519 7225 15531 7228
rect 15473 7219 15531 7225
rect 15746 7216 15752 7228
rect 15804 7256 15810 7268
rect 15933 7259 15991 7265
rect 15933 7256 15945 7259
rect 15804 7228 15945 7256
rect 15804 7216 15810 7228
rect 15933 7225 15945 7228
rect 15979 7225 15991 7259
rect 15933 7219 15991 7225
rect 17865 7259 17923 7265
rect 17865 7225 17877 7259
rect 17911 7256 17923 7259
rect 17911 7228 18552 7256
rect 17911 7225 17923 7228
rect 17865 7219 17923 7225
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 3510 7188 3516 7200
rect 2832 7160 3516 7188
rect 2832 7148 2838 7160
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 4154 7188 4160 7200
rect 4115 7160 4160 7188
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 4706 7188 4712 7200
rect 4667 7160 4712 7188
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 7558 7148 7564 7200
rect 7616 7188 7622 7200
rect 7742 7188 7748 7200
rect 7616 7160 7748 7188
rect 7616 7148 7622 7160
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 9214 7188 9220 7200
rect 9175 7160 9220 7188
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 10689 7191 10747 7197
rect 9732 7160 9777 7188
rect 9732 7148 9738 7160
rect 10689 7157 10701 7191
rect 10735 7188 10747 7191
rect 11241 7191 11299 7197
rect 11241 7188 11253 7191
rect 10735 7160 11253 7188
rect 10735 7157 10747 7160
rect 10689 7151 10747 7157
rect 11241 7157 11253 7160
rect 11287 7188 11299 7191
rect 11330 7188 11336 7200
rect 11287 7160 11336 7188
rect 11287 7157 11299 7160
rect 11241 7151 11299 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 12897 7191 12955 7197
rect 12897 7188 12909 7191
rect 12584 7160 12909 7188
rect 12584 7148 12590 7160
rect 12897 7157 12909 7160
rect 12943 7157 12955 7191
rect 12897 7151 12955 7157
rect 12986 7148 12992 7200
rect 13044 7188 13050 7200
rect 13449 7191 13507 7197
rect 13449 7188 13461 7191
rect 13044 7160 13461 7188
rect 13044 7148 13050 7160
rect 13449 7157 13461 7160
rect 13495 7157 13507 7191
rect 13449 7151 13507 7157
rect 13538 7148 13544 7200
rect 13596 7188 13602 7200
rect 13817 7191 13875 7197
rect 13817 7188 13829 7191
rect 13596 7160 13829 7188
rect 13596 7148 13602 7160
rect 13817 7157 13829 7160
rect 13863 7157 13875 7191
rect 13817 7151 13875 7157
rect 13906 7148 13912 7200
rect 13964 7188 13970 7200
rect 14001 7191 14059 7197
rect 14001 7188 14013 7191
rect 13964 7160 14013 7188
rect 13964 7148 13970 7160
rect 14001 7157 14013 7160
rect 14047 7157 14059 7191
rect 14001 7151 14059 7157
rect 14274 7148 14280 7200
rect 14332 7188 14338 7200
rect 14369 7191 14427 7197
rect 14369 7188 14381 7191
rect 14332 7160 14381 7188
rect 14332 7148 14338 7160
rect 14369 7157 14381 7160
rect 14415 7157 14427 7191
rect 15562 7188 15568 7200
rect 15523 7160 15568 7188
rect 14369 7151 14427 7157
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 17497 7191 17555 7197
rect 17497 7157 17509 7191
rect 17543 7188 17555 7191
rect 18414 7188 18420 7200
rect 17543 7160 18420 7188
rect 17543 7157 17555 7160
rect 17497 7151 17555 7157
rect 18414 7148 18420 7160
rect 18472 7148 18478 7200
rect 18524 7197 18552 7228
rect 19334 7216 19340 7268
rect 19392 7256 19398 7268
rect 20162 7256 20168 7268
rect 19392 7228 20168 7256
rect 19392 7216 19398 7228
rect 20162 7216 20168 7228
rect 20220 7216 20226 7268
rect 22557 7259 22615 7265
rect 22557 7225 22569 7259
rect 22603 7256 22615 7259
rect 22738 7256 22744 7268
rect 22603 7228 22744 7256
rect 22603 7225 22615 7228
rect 22557 7219 22615 7225
rect 22738 7216 22744 7228
rect 22796 7256 22802 7268
rect 23934 7256 23940 7268
rect 22796 7228 23940 7256
rect 22796 7216 22802 7228
rect 23934 7216 23940 7228
rect 23992 7216 23998 7268
rect 18509 7191 18567 7197
rect 18509 7157 18521 7191
rect 18555 7188 18567 7191
rect 18782 7188 18788 7200
rect 18555 7160 18788 7188
rect 18555 7157 18567 7160
rect 18509 7151 18567 7157
rect 18782 7148 18788 7160
rect 18840 7148 18846 7200
rect 19426 7148 19432 7200
rect 19484 7188 19490 7200
rect 19981 7191 20039 7197
rect 19981 7188 19993 7191
rect 19484 7160 19993 7188
rect 19484 7148 19490 7160
rect 19981 7157 19993 7160
rect 20027 7157 20039 7191
rect 19981 7151 20039 7157
rect 20717 7191 20775 7197
rect 20717 7157 20729 7191
rect 20763 7188 20775 7191
rect 20806 7188 20812 7200
rect 20763 7160 20812 7188
rect 20763 7157 20775 7160
rect 20717 7151 20775 7157
rect 20806 7148 20812 7160
rect 20864 7188 20870 7200
rect 21726 7188 21732 7200
rect 20864 7160 21732 7188
rect 20864 7148 20870 7160
rect 21726 7148 21732 7160
rect 21784 7148 21790 7200
rect 22002 7148 22008 7200
rect 22060 7188 22066 7200
rect 22094 7188 22100 7200
rect 22060 7160 22100 7188
rect 22060 7148 22066 7160
rect 22094 7148 22100 7160
rect 22152 7148 22158 7200
rect 23014 7148 23020 7200
rect 23072 7188 23078 7200
rect 23290 7188 23296 7200
rect 23072 7160 23296 7188
rect 23072 7148 23078 7160
rect 23290 7148 23296 7160
rect 23348 7148 23354 7200
rect 23845 7191 23903 7197
rect 23845 7157 23857 7191
rect 23891 7188 23903 7191
rect 24118 7188 24124 7200
rect 23891 7160 24124 7188
rect 23891 7157 23903 7160
rect 23845 7151 23903 7157
rect 24118 7148 24124 7160
rect 24176 7148 24182 7200
rect 24949 7191 25007 7197
rect 24949 7157 24961 7191
rect 24995 7188 25007 7191
rect 25958 7188 25964 7200
rect 24995 7160 25964 7188
rect 24995 7157 25007 7160
rect 24949 7151 25007 7157
rect 25958 7148 25964 7160
rect 26016 7148 26022 7200
rect 26142 7188 26148 7200
rect 26103 7160 26148 7188
rect 26142 7148 26148 7160
rect 26200 7148 26206 7200
rect 26418 7188 26424 7200
rect 26379 7160 26424 7188
rect 26418 7148 26424 7160
rect 26476 7148 26482 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1673 6987 1731 6993
rect 1673 6953 1685 6987
rect 1719 6984 1731 6987
rect 1946 6984 1952 6996
rect 1719 6956 1952 6984
rect 1719 6953 1731 6956
rect 1673 6947 1731 6953
rect 1946 6944 1952 6956
rect 2004 6944 2010 6996
rect 2777 6987 2835 6993
rect 2777 6953 2789 6987
rect 2823 6984 2835 6987
rect 4062 6984 4068 6996
rect 2823 6956 4068 6984
rect 2823 6953 2835 6956
rect 2777 6947 2835 6953
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 4430 6984 4436 6996
rect 4391 6956 4436 6984
rect 4430 6944 4436 6956
rect 4488 6944 4494 6996
rect 6270 6944 6276 6996
rect 6328 6984 6334 6996
rect 6457 6987 6515 6993
rect 6457 6984 6469 6987
rect 6328 6956 6469 6984
rect 6328 6944 6334 6956
rect 6457 6953 6469 6956
rect 6503 6984 6515 6987
rect 7098 6984 7104 6996
rect 6503 6956 7104 6984
rect 6503 6953 6515 6956
rect 6457 6947 6515 6953
rect 7098 6944 7104 6956
rect 7156 6944 7162 6996
rect 9309 6987 9367 6993
rect 9309 6953 9321 6987
rect 9355 6984 9367 6987
rect 9766 6984 9772 6996
rect 9355 6956 9772 6984
rect 9355 6953 9367 6956
rect 9309 6947 9367 6953
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 11790 6984 11796 6996
rect 11751 6956 11796 6984
rect 11790 6944 11796 6956
rect 11848 6944 11854 6996
rect 12526 6984 12532 6996
rect 12487 6956 12532 6984
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 13998 6984 14004 6996
rect 13959 6956 14004 6984
rect 13998 6944 14004 6956
rect 14056 6944 14062 6996
rect 18690 6944 18696 6996
rect 18748 6984 18754 6996
rect 19334 6984 19340 6996
rect 18748 6956 19340 6984
rect 18748 6944 18754 6956
rect 19334 6944 19340 6956
rect 19392 6944 19398 6996
rect 21266 6984 21272 6996
rect 21227 6956 21272 6984
rect 21266 6944 21272 6956
rect 21324 6944 21330 6996
rect 22370 6944 22376 6996
rect 22428 6984 22434 6996
rect 22465 6987 22523 6993
rect 22465 6984 22477 6987
rect 22428 6956 22477 6984
rect 22428 6944 22434 6956
rect 22465 6953 22477 6956
rect 22511 6953 22523 6987
rect 22830 6984 22836 6996
rect 22791 6956 22836 6984
rect 22465 6947 22523 6953
rect 22830 6944 22836 6956
rect 22888 6944 22894 6996
rect 23658 6984 23664 6996
rect 22940 6956 23664 6984
rect 2314 6876 2320 6928
rect 2372 6916 2378 6928
rect 2869 6919 2927 6925
rect 2869 6916 2881 6919
rect 2372 6888 2881 6916
rect 2372 6876 2378 6888
rect 2869 6885 2881 6888
rect 2915 6885 2927 6919
rect 2869 6879 2927 6885
rect 3142 6876 3148 6928
rect 3200 6916 3206 6928
rect 3694 6916 3700 6928
rect 3200 6888 3700 6916
rect 3200 6876 3206 6888
rect 3694 6876 3700 6888
rect 3752 6876 3758 6928
rect 6178 6876 6184 6928
rect 6236 6916 6242 6928
rect 6236 6888 6592 6916
rect 6236 6876 6242 6888
rect 4525 6851 4583 6857
rect 4525 6817 4537 6851
rect 4571 6848 4583 6851
rect 4706 6848 4712 6860
rect 4571 6820 4712 6848
rect 4571 6817 4583 6820
rect 4525 6811 4583 6817
rect 4706 6808 4712 6820
rect 4764 6848 4770 6860
rect 6270 6848 6276 6860
rect 4764 6820 6276 6848
rect 4764 6808 4770 6820
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 6564 6848 6592 6888
rect 10410 6876 10416 6928
rect 10468 6916 10474 6928
rect 11606 6916 11612 6928
rect 10468 6888 11612 6916
rect 10468 6876 10474 6888
rect 11606 6876 11612 6888
rect 11664 6876 11670 6928
rect 13262 6916 13268 6928
rect 13223 6888 13268 6916
rect 13262 6876 13268 6888
rect 13320 6876 13326 6928
rect 18598 6876 18604 6928
rect 18656 6916 18662 6928
rect 18966 6916 18972 6928
rect 18656 6888 18972 6916
rect 18656 6876 18662 6888
rect 18966 6876 18972 6888
rect 19024 6876 19030 6928
rect 19429 6919 19487 6925
rect 19429 6916 19441 6919
rect 19260 6888 19441 6916
rect 7653 6851 7711 6857
rect 6564 6820 6684 6848
rect 2961 6783 3019 6789
rect 2961 6749 2973 6783
rect 3007 6780 3019 6783
rect 3234 6780 3240 6792
rect 3007 6752 3240 6780
rect 3007 6749 3019 6752
rect 2961 6743 3019 6749
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 4614 6780 4620 6792
rect 4575 6752 4620 6780
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 5258 6780 5264 6792
rect 5219 6752 5264 6780
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 5994 6740 6000 6792
rect 6052 6780 6058 6792
rect 6656 6789 6684 6820
rect 7653 6817 7665 6851
rect 7699 6848 7711 6851
rect 7742 6848 7748 6860
rect 7699 6820 7748 6848
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 7742 6808 7748 6820
rect 7800 6808 7806 6860
rect 8110 6848 8116 6860
rect 8071 6820 8116 6848
rect 8110 6808 8116 6820
rect 8168 6808 8174 6860
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 10321 6851 10379 6857
rect 8260 6820 8305 6848
rect 8260 6808 8266 6820
rect 10321 6817 10333 6851
rect 10367 6848 10379 6851
rect 10669 6851 10727 6857
rect 10669 6848 10681 6851
rect 10367 6820 10681 6848
rect 10367 6817 10379 6820
rect 10321 6811 10379 6817
rect 10669 6817 10681 6820
rect 10715 6848 10727 6851
rect 11146 6848 11152 6860
rect 10715 6820 11152 6848
rect 10715 6817 10727 6820
rect 10669 6811 10727 6817
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 13004 6820 13584 6848
rect 6549 6783 6607 6789
rect 6549 6780 6561 6783
rect 6052 6752 6561 6780
rect 6052 6740 6058 6752
rect 6549 6749 6561 6752
rect 6595 6749 6607 6783
rect 6549 6743 6607 6749
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6780 6699 6783
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 6687 6752 8309 6780
rect 6687 6749 6699 6752
rect 6641 6743 6699 6749
rect 8297 6749 8309 6752
rect 8343 6780 8355 6783
rect 8662 6780 8668 6792
rect 8343 6752 8668 6780
rect 8343 6749 8355 6752
rect 8297 6743 8355 6749
rect 8662 6740 8668 6752
rect 8720 6780 8726 6792
rect 8757 6783 8815 6789
rect 8757 6780 8769 6783
rect 8720 6752 8769 6780
rect 8720 6740 8726 6752
rect 8757 6749 8769 6752
rect 8803 6749 8815 6783
rect 8757 6743 8815 6749
rect 9030 6740 9036 6792
rect 9088 6780 9094 6792
rect 9214 6780 9220 6792
rect 9088 6752 9220 6780
rect 9088 6740 9094 6752
rect 9214 6740 9220 6752
rect 9272 6780 9278 6792
rect 10413 6783 10471 6789
rect 10413 6780 10425 6783
rect 9272 6752 10425 6780
rect 9272 6740 9278 6752
rect 10413 6749 10425 6752
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 2406 6712 2412 6724
rect 2367 6684 2412 6712
rect 2406 6672 2412 6684
rect 2464 6672 2470 6724
rect 3050 6672 3056 6724
rect 3108 6712 3114 6724
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 3108 6684 3801 6712
rect 3108 6672 3114 6684
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 5905 6715 5963 6721
rect 5905 6712 5917 6715
rect 3789 6675 3847 6681
rect 3896 6684 5917 6712
rect 2314 6644 2320 6656
rect 2275 6616 2320 6644
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 2832 6616 3433 6644
rect 2832 6604 2838 6616
rect 3421 6613 3433 6616
rect 3467 6613 3479 6647
rect 3421 6607 3479 6613
rect 3694 6604 3700 6656
rect 3752 6644 3758 6656
rect 3896 6644 3924 6684
rect 5905 6681 5917 6684
rect 5951 6681 5963 6715
rect 6086 6712 6092 6724
rect 6047 6684 6092 6712
rect 5905 6675 5963 6681
rect 6086 6672 6092 6684
rect 6144 6672 6150 6724
rect 7745 6715 7803 6721
rect 7745 6712 7757 6715
rect 6564 6684 7757 6712
rect 6564 6656 6592 6684
rect 7745 6681 7757 6684
rect 7791 6681 7803 6715
rect 7745 6675 7803 6681
rect 8938 6672 8944 6724
rect 8996 6712 9002 6724
rect 9490 6712 9496 6724
rect 8996 6684 9496 6712
rect 8996 6672 9002 6684
rect 9490 6672 9496 6684
rect 9548 6712 9554 6724
rect 9548 6684 10364 6712
rect 9548 6672 9554 6684
rect 3752 6616 3924 6644
rect 3752 6604 3758 6616
rect 4890 6604 4896 6656
rect 4948 6644 4954 6656
rect 5537 6647 5595 6653
rect 5537 6644 5549 6647
rect 4948 6616 5549 6644
rect 4948 6604 4954 6616
rect 5537 6613 5549 6616
rect 5583 6613 5595 6647
rect 5537 6607 5595 6613
rect 6546 6604 6552 6656
rect 6604 6604 6610 6656
rect 7285 6647 7343 6653
rect 7285 6613 7297 6647
rect 7331 6644 7343 6647
rect 7374 6644 7380 6656
rect 7331 6616 7380 6644
rect 7331 6613 7343 6616
rect 7285 6607 7343 6613
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 9766 6604 9772 6656
rect 9824 6644 9830 6656
rect 9861 6647 9919 6653
rect 9861 6644 9873 6647
rect 9824 6616 9873 6644
rect 9824 6604 9830 6616
rect 9861 6613 9873 6616
rect 9907 6613 9919 6647
rect 9861 6607 9919 6613
rect 9950 6604 9956 6656
rect 10008 6644 10014 6656
rect 10134 6644 10140 6656
rect 10008 6616 10140 6644
rect 10008 6604 10014 6616
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 10336 6644 10364 6684
rect 11790 6672 11796 6724
rect 11848 6712 11854 6724
rect 12710 6712 12716 6724
rect 11848 6684 12716 6712
rect 11848 6672 11854 6684
rect 12710 6672 12716 6684
rect 12768 6712 12774 6724
rect 13004 6712 13032 6820
rect 13556 6792 13584 6820
rect 14642 6808 14648 6860
rect 14700 6848 14706 6860
rect 15013 6851 15071 6857
rect 15013 6848 15025 6851
rect 14700 6820 15025 6848
rect 14700 6808 14706 6820
rect 15013 6817 15025 6820
rect 15059 6817 15071 6851
rect 15470 6848 15476 6860
rect 15431 6820 15476 6848
rect 15013 6811 15071 6817
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 16482 6848 16488 6860
rect 16443 6820 16488 6848
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 16666 6808 16672 6860
rect 16724 6848 16730 6860
rect 16844 6851 16902 6857
rect 16844 6848 16856 6851
rect 16724 6820 16856 6848
rect 16724 6808 16730 6820
rect 16844 6817 16856 6820
rect 16890 6848 16902 6851
rect 17862 6848 17868 6860
rect 16890 6820 17868 6848
rect 16890 6817 16902 6820
rect 16844 6811 16902 6817
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 17954 6808 17960 6860
rect 18012 6848 18018 6860
rect 19150 6848 19156 6860
rect 18012 6820 19156 6848
rect 18012 6808 18018 6820
rect 19150 6808 19156 6820
rect 19208 6848 19214 6860
rect 19260 6848 19288 6888
rect 19429 6885 19441 6888
rect 19475 6885 19487 6919
rect 19429 6879 19487 6885
rect 19889 6919 19947 6925
rect 19889 6885 19901 6919
rect 19935 6916 19947 6919
rect 22940 6916 22968 6956
rect 23658 6944 23664 6956
rect 23716 6944 23722 6996
rect 24026 6944 24032 6996
rect 24084 6944 24090 6996
rect 24762 6984 24768 6996
rect 24723 6956 24768 6984
rect 24762 6944 24768 6956
rect 24820 6944 24826 6996
rect 24044 6916 24072 6944
rect 19935 6888 22968 6916
rect 23400 6888 24072 6916
rect 19935 6885 19947 6888
rect 19889 6879 19947 6885
rect 22388 6860 22416 6888
rect 19208 6820 19288 6848
rect 19352 6820 19840 6848
rect 19208 6808 19214 6820
rect 13354 6780 13360 6792
rect 13315 6752 13360 6780
rect 13354 6740 13360 6752
rect 13412 6740 13418 6792
rect 13538 6780 13544 6792
rect 13499 6752 13544 6780
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 15286 6740 15292 6792
rect 15344 6780 15350 6792
rect 16114 6780 16120 6792
rect 15344 6752 16120 6780
rect 15344 6740 15350 6752
rect 16114 6740 16120 6752
rect 16172 6780 16178 6792
rect 16577 6783 16635 6789
rect 16577 6780 16589 6783
rect 16172 6752 16589 6780
rect 16172 6740 16178 6752
rect 16577 6749 16589 6752
rect 16623 6749 16635 6783
rect 16577 6743 16635 6749
rect 18230 6740 18236 6792
rect 18288 6780 18294 6792
rect 18601 6783 18659 6789
rect 18601 6780 18613 6783
rect 18288 6752 18613 6780
rect 18288 6740 18294 6752
rect 18601 6749 18613 6752
rect 18647 6780 18659 6783
rect 19352 6780 19380 6820
rect 18647 6752 19380 6780
rect 19521 6783 19579 6789
rect 18647 6749 18659 6752
rect 18601 6743 18659 6749
rect 19521 6749 19533 6783
rect 19567 6780 19579 6783
rect 19610 6780 19616 6792
rect 19567 6752 19616 6780
rect 19567 6749 19579 6752
rect 19521 6743 19579 6749
rect 19610 6740 19616 6752
rect 19668 6740 19674 6792
rect 19705 6783 19763 6789
rect 19705 6749 19717 6783
rect 19751 6749 19763 6783
rect 19812 6780 19840 6820
rect 22370 6808 22376 6860
rect 22428 6808 22434 6860
rect 22738 6808 22744 6860
rect 22796 6848 22802 6860
rect 23400 6848 23428 6888
rect 24026 6848 24032 6860
rect 22796 6820 23428 6848
rect 23987 6820 24032 6848
rect 22796 6808 22802 6820
rect 24026 6808 24032 6820
rect 24084 6808 24090 6860
rect 25133 6851 25191 6857
rect 25133 6817 25145 6851
rect 25179 6817 25191 6851
rect 25133 6811 25191 6817
rect 21174 6780 21180 6792
rect 19812 6752 21180 6780
rect 19705 6743 19763 6749
rect 12768 6684 13032 6712
rect 13372 6712 13400 6740
rect 14369 6715 14427 6721
rect 14369 6712 14381 6715
rect 13372 6684 14381 6712
rect 12768 6672 12774 6684
rect 14369 6681 14381 6684
rect 14415 6681 14427 6715
rect 14369 6675 14427 6681
rect 14734 6672 14740 6724
rect 14792 6712 14798 6724
rect 18877 6715 18935 6721
rect 18877 6712 18889 6715
rect 14792 6684 16436 6712
rect 14792 6672 14798 6684
rect 12526 6644 12532 6656
rect 10336 6616 12532 6644
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 12897 6647 12955 6653
rect 12897 6613 12909 6647
rect 12943 6644 12955 6647
rect 13722 6644 13728 6656
rect 12943 6616 13728 6644
rect 12943 6613 12955 6616
rect 12897 6607 12955 6613
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 15654 6644 15660 6656
rect 15615 6616 15660 6644
rect 15654 6604 15660 6616
rect 15712 6604 15718 6656
rect 16114 6644 16120 6656
rect 16075 6616 16120 6644
rect 16114 6604 16120 6616
rect 16172 6604 16178 6656
rect 16408 6644 16436 6684
rect 17604 6684 18889 6712
rect 17604 6644 17632 6684
rect 18877 6681 18889 6684
rect 18923 6712 18935 6715
rect 19720 6712 19748 6743
rect 21174 6740 21180 6752
rect 21232 6740 21238 6792
rect 21358 6780 21364 6792
rect 21319 6752 21364 6780
rect 21358 6740 21364 6752
rect 21416 6740 21422 6792
rect 21453 6783 21511 6789
rect 21453 6749 21465 6783
rect 21499 6749 21511 6783
rect 21453 6743 21511 6749
rect 20898 6712 20904 6724
rect 18923 6684 20208 6712
rect 20859 6684 20904 6712
rect 18923 6681 18935 6684
rect 18877 6675 18935 6681
rect 20180 6656 20208 6684
rect 20898 6672 20904 6684
rect 20956 6672 20962 6724
rect 21468 6712 21496 6743
rect 22554 6740 22560 6792
rect 22612 6780 22618 6792
rect 22925 6783 22983 6789
rect 22925 6780 22937 6783
rect 22612 6752 22937 6780
rect 22612 6740 22618 6752
rect 22925 6749 22937 6752
rect 22971 6749 22983 6783
rect 22925 6743 22983 6749
rect 23109 6783 23167 6789
rect 23109 6749 23121 6783
rect 23155 6780 23167 6783
rect 23290 6780 23296 6792
rect 23155 6752 23296 6780
rect 23155 6749 23167 6752
rect 23109 6743 23167 6749
rect 23290 6740 23296 6752
rect 23348 6780 23354 6792
rect 23750 6780 23756 6792
rect 23348 6752 23756 6780
rect 23348 6740 23354 6752
rect 23750 6740 23756 6752
rect 23808 6740 23814 6792
rect 21913 6715 21971 6721
rect 21913 6712 21925 6715
rect 21008 6684 21925 6712
rect 21008 6656 21036 6684
rect 21913 6681 21925 6684
rect 21959 6681 21971 6715
rect 21913 6675 21971 6681
rect 22002 6672 22008 6724
rect 22060 6712 22066 6724
rect 25148 6712 25176 6811
rect 25222 6740 25228 6792
rect 25280 6780 25286 6792
rect 25685 6783 25743 6789
rect 25685 6780 25697 6783
rect 25280 6752 25697 6780
rect 25280 6740 25286 6752
rect 25685 6749 25697 6752
rect 25731 6749 25743 6783
rect 25685 6743 25743 6749
rect 25774 6712 25780 6724
rect 22060 6684 25780 6712
rect 22060 6672 22066 6684
rect 25774 6672 25780 6684
rect 25832 6672 25838 6724
rect 17954 6644 17960 6656
rect 16408 6616 17632 6644
rect 17915 6616 17960 6644
rect 17954 6604 17960 6616
rect 18012 6604 18018 6656
rect 19058 6644 19064 6656
rect 19019 6616 19064 6644
rect 19058 6604 19064 6616
rect 19116 6604 19122 6656
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 19889 6647 19947 6653
rect 19889 6644 19901 6647
rect 19392 6616 19901 6644
rect 19392 6604 19398 6616
rect 19889 6613 19901 6616
rect 19935 6613 19947 6647
rect 20162 6644 20168 6656
rect 20123 6616 20168 6644
rect 19889 6607 19947 6613
rect 20162 6604 20168 6616
rect 20220 6604 20226 6656
rect 20717 6647 20775 6653
rect 20717 6613 20729 6647
rect 20763 6644 20775 6647
rect 20990 6644 20996 6656
rect 20763 6616 20996 6644
rect 20763 6613 20775 6616
rect 20717 6607 20775 6613
rect 20990 6604 20996 6616
rect 21048 6604 21054 6656
rect 22278 6644 22284 6656
rect 22239 6616 22284 6644
rect 22278 6604 22284 6616
rect 22336 6604 22342 6656
rect 23750 6644 23756 6656
rect 23711 6616 23756 6644
rect 23750 6604 23756 6616
rect 23808 6604 23814 6656
rect 23842 6604 23848 6656
rect 23900 6644 23906 6656
rect 24213 6647 24271 6653
rect 24213 6644 24225 6647
rect 23900 6616 24225 6644
rect 23900 6604 23906 6616
rect 24213 6613 24225 6616
rect 24259 6613 24271 6647
rect 24213 6607 24271 6613
rect 24854 6604 24860 6656
rect 24912 6644 24918 6656
rect 25317 6647 25375 6653
rect 25317 6644 25329 6647
rect 24912 6616 25329 6644
rect 24912 6604 24918 6616
rect 25317 6613 25329 6616
rect 25363 6613 25375 6647
rect 26050 6644 26056 6656
rect 26011 6616 26056 6644
rect 25317 6607 25375 6613
rect 26050 6604 26056 6616
rect 26108 6604 26114 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2225 6443 2283 6449
rect 2225 6409 2237 6443
rect 2271 6440 2283 6443
rect 2498 6440 2504 6452
rect 2271 6412 2504 6440
rect 2271 6409 2283 6412
rect 2225 6403 2283 6409
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 3234 6440 3240 6452
rect 3195 6412 3240 6440
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 5994 6400 6000 6452
rect 6052 6440 6058 6452
rect 6089 6443 6147 6449
rect 6089 6440 6101 6443
rect 6052 6412 6101 6440
rect 6052 6400 6058 6412
rect 6089 6409 6101 6412
rect 6135 6409 6147 6443
rect 6089 6403 6147 6409
rect 6549 6443 6607 6449
rect 6549 6409 6561 6443
rect 6595 6440 6607 6443
rect 7098 6440 7104 6452
rect 6595 6412 7104 6440
rect 6595 6409 6607 6412
rect 6549 6403 6607 6409
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 7745 6443 7803 6449
rect 7745 6409 7757 6443
rect 7791 6440 7803 6443
rect 8110 6440 8116 6452
rect 7791 6412 8116 6440
rect 7791 6409 7803 6412
rect 7745 6403 7803 6409
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 10008 6412 10057 6440
rect 10008 6400 10014 6412
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 10594 6440 10600 6452
rect 10555 6412 10600 6440
rect 10045 6403 10103 6409
rect 5813 6375 5871 6381
rect 5813 6341 5825 6375
rect 5859 6372 5871 6375
rect 6178 6372 6184 6384
rect 5859 6344 6184 6372
rect 5859 6341 5871 6344
rect 5813 6335 5871 6341
rect 6178 6332 6184 6344
rect 6236 6332 6242 6384
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6304 1731 6307
rect 2222 6304 2228 6316
rect 1719 6276 2228 6304
rect 1719 6273 1731 6276
rect 1673 6267 1731 6273
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 2314 6264 2320 6316
rect 2372 6304 2378 6316
rect 2869 6307 2927 6313
rect 2869 6304 2881 6307
rect 2372 6276 2881 6304
rect 2372 6264 2378 6276
rect 2869 6273 2881 6276
rect 2915 6304 2927 6307
rect 6822 6304 6828 6316
rect 2915 6276 3924 6304
rect 6783 6276 6828 6304
rect 2915 6273 2927 6276
rect 2869 6267 2927 6273
rect 2590 6236 2596 6248
rect 2551 6208 2596 6236
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 3234 6196 3240 6248
rect 3292 6236 3298 6248
rect 3697 6239 3755 6245
rect 3697 6236 3709 6239
rect 3292 6208 3709 6236
rect 3292 6196 3298 6208
rect 3697 6205 3709 6208
rect 3743 6236 3755 6239
rect 3789 6239 3847 6245
rect 3789 6236 3801 6239
rect 3743 6208 3801 6236
rect 3743 6205 3755 6208
rect 3697 6199 3755 6205
rect 3789 6205 3801 6208
rect 3835 6205 3847 6239
rect 3896 6236 3924 6276
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 4062 6245 4068 6248
rect 4056 6236 4068 6245
rect 3896 6208 4068 6236
rect 3789 6199 3847 6205
rect 4056 6199 4068 6208
rect 3804 6168 3832 6199
rect 4062 6196 4068 6199
rect 4120 6196 4126 6248
rect 7742 6196 7748 6248
rect 7800 6236 7806 6248
rect 7837 6239 7895 6245
rect 7837 6236 7849 6239
rect 7800 6208 7849 6236
rect 7800 6196 7806 6208
rect 7837 6205 7849 6208
rect 7883 6205 7895 6239
rect 7837 6199 7895 6205
rect 4246 6168 4252 6180
rect 3804 6140 4252 6168
rect 4246 6128 4252 6140
rect 4304 6128 4310 6180
rect 7374 6128 7380 6180
rect 7432 6168 7438 6180
rect 8104 6171 8162 6177
rect 8104 6168 8116 6171
rect 7432 6140 8116 6168
rect 7432 6128 7438 6140
rect 8104 6137 8116 6140
rect 8150 6168 8162 6171
rect 8294 6168 8300 6180
rect 8150 6140 8300 6168
rect 8150 6137 8162 6140
rect 8104 6131 8162 6137
rect 8294 6128 8300 6140
rect 8352 6128 8358 6180
rect 10060 6168 10088 6403
rect 10594 6400 10600 6412
rect 10652 6400 10658 6452
rect 13262 6400 13268 6452
rect 13320 6440 13326 6452
rect 15013 6443 15071 6449
rect 15013 6440 15025 6443
rect 13320 6412 15025 6440
rect 13320 6400 13326 6412
rect 15013 6409 15025 6412
rect 15059 6409 15071 6443
rect 15013 6403 15071 6409
rect 15562 6400 15568 6452
rect 15620 6440 15626 6452
rect 15841 6443 15899 6449
rect 15841 6440 15853 6443
rect 15620 6412 15853 6440
rect 15620 6400 15626 6412
rect 15841 6409 15853 6412
rect 15887 6409 15899 6443
rect 15841 6403 15899 6409
rect 15930 6400 15936 6452
rect 15988 6440 15994 6452
rect 16393 6443 16451 6449
rect 16393 6440 16405 6443
rect 15988 6412 16405 6440
rect 15988 6400 15994 6412
rect 16393 6409 16405 6412
rect 16439 6409 16451 6443
rect 16393 6403 16451 6409
rect 16850 6400 16856 6452
rect 16908 6440 16914 6452
rect 18049 6443 18107 6449
rect 18049 6440 18061 6443
rect 16908 6412 18061 6440
rect 16908 6400 16914 6412
rect 18049 6409 18061 6412
rect 18095 6409 18107 6443
rect 18049 6403 18107 6409
rect 21082 6400 21088 6452
rect 21140 6440 21146 6452
rect 22554 6440 22560 6452
rect 21140 6412 22560 6440
rect 21140 6400 21146 6412
rect 22554 6400 22560 6412
rect 22612 6400 22618 6452
rect 22830 6440 22836 6452
rect 22791 6412 22836 6440
rect 22830 6400 22836 6412
rect 22888 6400 22894 6452
rect 24026 6400 24032 6452
rect 24084 6440 24090 6452
rect 24673 6443 24731 6449
rect 24673 6440 24685 6443
rect 24084 6412 24685 6440
rect 24084 6400 24090 6412
rect 24673 6409 24685 6412
rect 24719 6409 24731 6443
rect 25038 6440 25044 6452
rect 24999 6412 25044 6440
rect 24673 6403 24731 6409
rect 25038 6400 25044 6412
rect 25096 6400 25102 6452
rect 25774 6440 25780 6452
rect 25735 6412 25780 6440
rect 25774 6400 25780 6412
rect 25832 6400 25838 6452
rect 10502 6372 10508 6384
rect 10463 6344 10508 6372
rect 10502 6332 10508 6344
rect 10560 6372 10566 6384
rect 14461 6375 14519 6381
rect 10560 6344 11008 6372
rect 10560 6332 10566 6344
rect 10980 6245 11008 6344
rect 14461 6341 14473 6375
rect 14507 6372 14519 6375
rect 14550 6372 14556 6384
rect 14507 6344 14556 6372
rect 14507 6341 14519 6344
rect 14461 6335 14519 6341
rect 14550 6332 14556 6344
rect 14608 6332 14614 6384
rect 17862 6372 17868 6384
rect 17775 6344 17868 6372
rect 17862 6332 17868 6344
rect 17920 6372 17926 6384
rect 19610 6372 19616 6384
rect 17920 6344 18736 6372
rect 17920 6332 17926 6344
rect 11146 6304 11152 6316
rect 11107 6276 11152 6304
rect 11146 6264 11152 6276
rect 11204 6304 11210 6316
rect 11977 6307 12035 6313
rect 11977 6304 11989 6307
rect 11204 6276 11989 6304
rect 11204 6264 11210 6276
rect 11977 6273 11989 6276
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6304 16359 6307
rect 17037 6307 17095 6313
rect 17037 6304 17049 6307
rect 16347 6276 17049 6304
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 17037 6273 17049 6276
rect 17083 6304 17095 6307
rect 17126 6304 17132 6316
rect 17083 6276 17132 6304
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 17126 6264 17132 6276
rect 17184 6304 17190 6316
rect 17954 6304 17960 6316
rect 17184 6276 17960 6304
rect 17184 6264 17190 6276
rect 17954 6264 17960 6276
rect 18012 6264 18018 6316
rect 18230 6264 18236 6316
rect 18288 6304 18294 6316
rect 18708 6313 18736 6344
rect 19352 6344 19616 6372
rect 18509 6307 18567 6313
rect 18509 6304 18521 6307
rect 18288 6276 18521 6304
rect 18288 6264 18294 6276
rect 18509 6273 18521 6276
rect 18555 6273 18567 6307
rect 18509 6267 18567 6273
rect 18693 6307 18751 6313
rect 18693 6273 18705 6307
rect 18739 6304 18751 6307
rect 18966 6304 18972 6316
rect 18739 6276 18972 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 18966 6264 18972 6276
rect 19024 6264 19030 6316
rect 19153 6307 19211 6313
rect 19153 6273 19165 6307
rect 19199 6304 19211 6307
rect 19352 6304 19380 6344
rect 19610 6332 19616 6344
rect 19668 6332 19674 6384
rect 20993 6375 21051 6381
rect 20993 6341 21005 6375
rect 21039 6372 21051 6375
rect 21266 6372 21272 6384
rect 21039 6344 21272 6372
rect 21039 6341 21051 6344
rect 20993 6335 21051 6341
rect 21266 6332 21272 6344
rect 21324 6332 21330 6384
rect 19199 6276 19380 6304
rect 19199 6273 19211 6276
rect 19153 6267 19211 6273
rect 10965 6239 11023 6245
rect 10965 6205 10977 6239
rect 11011 6205 11023 6239
rect 12986 6236 12992 6248
rect 12899 6208 12992 6236
rect 10965 6199 11023 6205
rect 11057 6171 11115 6177
rect 11057 6168 11069 6171
rect 10060 6140 11069 6168
rect 11057 6137 11069 6140
rect 11103 6137 11115 6171
rect 11057 6131 11115 6137
rect 2133 6103 2191 6109
rect 2133 6069 2145 6103
rect 2179 6100 2191 6103
rect 2685 6103 2743 6109
rect 2685 6100 2697 6103
rect 2179 6072 2697 6100
rect 2179 6069 2191 6072
rect 2133 6063 2191 6069
rect 2685 6069 2697 6072
rect 2731 6100 2743 6103
rect 3142 6100 3148 6112
rect 2731 6072 3148 6100
rect 2731 6069 2743 6072
rect 2685 6063 2743 6069
rect 3142 6060 3148 6072
rect 3200 6060 3206 6112
rect 5169 6103 5227 6109
rect 5169 6069 5181 6103
rect 5215 6100 5227 6103
rect 5442 6100 5448 6112
rect 5215 6072 5448 6100
rect 5215 6069 5227 6072
rect 5169 6063 5227 6069
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 7285 6103 7343 6109
rect 7285 6069 7297 6103
rect 7331 6100 7343 6103
rect 8202 6100 8208 6112
rect 7331 6072 8208 6100
rect 7331 6069 7343 6072
rect 7285 6063 7343 6069
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 9217 6103 9275 6109
rect 9217 6069 9229 6103
rect 9263 6100 9275 6103
rect 9950 6100 9956 6112
rect 9263 6072 9956 6100
rect 9263 6069 9275 6072
rect 9217 6063 9275 6069
rect 9950 6060 9956 6072
rect 10008 6060 10014 6112
rect 11701 6103 11759 6109
rect 11701 6069 11713 6103
rect 11747 6100 11759 6103
rect 11790 6100 11796 6112
rect 11747 6072 11796 6100
rect 11747 6069 11759 6072
rect 11701 6063 11759 6069
rect 11790 6060 11796 6072
rect 11848 6100 11854 6112
rect 12912 6109 12940 6208
rect 12986 6196 12992 6208
rect 13044 6236 13050 6248
rect 13081 6239 13139 6245
rect 13081 6236 13093 6239
rect 13044 6208 13093 6236
rect 13044 6196 13050 6208
rect 13081 6205 13093 6208
rect 13127 6205 13139 6239
rect 13081 6199 13139 6205
rect 13348 6239 13406 6245
rect 13348 6205 13360 6239
rect 13394 6236 13406 6239
rect 14090 6236 14096 6248
rect 13394 6208 14096 6236
rect 13394 6205 13406 6208
rect 13348 6199 13406 6205
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 16850 6236 16856 6248
rect 16811 6208 16856 6236
rect 16850 6196 16856 6208
rect 16908 6196 16914 6248
rect 18414 6236 18420 6248
rect 18327 6208 18420 6236
rect 18414 6196 18420 6208
rect 18472 6236 18478 6248
rect 19242 6236 19248 6248
rect 18472 6208 19248 6236
rect 18472 6196 18478 6208
rect 19242 6196 19248 6208
rect 19300 6196 19306 6248
rect 16758 6168 16764 6180
rect 16719 6140 16764 6168
rect 16758 6128 16764 6140
rect 16816 6128 16822 6180
rect 18046 6128 18052 6180
rect 18104 6168 18110 6180
rect 19352 6168 19380 6276
rect 19518 6264 19524 6316
rect 19576 6304 19582 6316
rect 19978 6304 19984 6316
rect 19576 6276 19984 6304
rect 19576 6264 19582 6276
rect 19978 6264 19984 6276
rect 20036 6304 20042 6316
rect 20073 6307 20131 6313
rect 20073 6304 20085 6307
rect 20036 6276 20085 6304
rect 20036 6264 20042 6276
rect 20073 6273 20085 6276
rect 20119 6273 20131 6307
rect 20073 6267 20131 6273
rect 20162 6264 20168 6316
rect 20220 6304 20226 6316
rect 20257 6307 20315 6313
rect 20257 6304 20269 6307
rect 20220 6276 20269 6304
rect 20220 6264 20226 6276
rect 20257 6273 20269 6276
rect 20303 6304 20315 6307
rect 20530 6304 20536 6316
rect 20303 6276 20536 6304
rect 20303 6273 20315 6276
rect 20257 6267 20315 6273
rect 20530 6264 20536 6276
rect 20588 6264 20594 6316
rect 21082 6264 21088 6316
rect 21140 6304 21146 6316
rect 21729 6307 21787 6313
rect 21729 6304 21741 6307
rect 21140 6276 21741 6304
rect 21140 6264 21146 6276
rect 21729 6273 21741 6276
rect 21775 6273 21787 6307
rect 21729 6267 21787 6273
rect 23750 6264 23756 6316
rect 23808 6304 23814 6316
rect 24026 6304 24032 6316
rect 23808 6276 24032 6304
rect 23808 6264 23814 6276
rect 24026 6264 24032 6276
rect 24084 6304 24090 6316
rect 24213 6307 24271 6313
rect 24213 6304 24225 6307
rect 24084 6276 24225 6304
rect 24084 6264 24090 6276
rect 24213 6273 24225 6276
rect 24259 6273 24271 6307
rect 24213 6267 24271 6273
rect 19426 6196 19432 6248
rect 19484 6236 19490 6248
rect 21542 6236 21548 6248
rect 19484 6208 20116 6236
rect 21503 6208 21548 6236
rect 19484 6196 19490 6208
rect 19981 6171 20039 6177
rect 19981 6168 19993 6171
rect 18104 6140 19380 6168
rect 19444 6140 19993 6168
rect 18104 6128 18110 6140
rect 19444 6112 19472 6140
rect 19981 6137 19993 6140
rect 20027 6137 20039 6171
rect 20088 6168 20116 6208
rect 21542 6196 21548 6208
rect 21600 6196 21606 6248
rect 22554 6196 22560 6248
rect 22612 6236 22618 6248
rect 23658 6236 23664 6248
rect 22612 6208 23664 6236
rect 22612 6196 22618 6208
rect 23658 6196 23664 6208
rect 23716 6196 23722 6248
rect 24121 6239 24179 6245
rect 24121 6205 24133 6239
rect 24167 6236 24179 6239
rect 24302 6236 24308 6248
rect 24167 6208 24308 6236
rect 24167 6205 24179 6208
rect 24121 6199 24179 6205
rect 24302 6196 24308 6208
rect 24360 6236 24366 6248
rect 24762 6236 24768 6248
rect 24360 6208 24768 6236
rect 24360 6196 24366 6208
rect 24762 6196 24768 6208
rect 24820 6196 24826 6248
rect 25038 6196 25044 6248
rect 25096 6236 25102 6248
rect 25225 6239 25283 6245
rect 25225 6236 25237 6239
rect 25096 6208 25237 6236
rect 25096 6196 25102 6208
rect 25225 6205 25237 6208
rect 25271 6205 25283 6239
rect 25225 6199 25283 6205
rect 23290 6168 23296 6180
rect 20088 6140 23296 6168
rect 19981 6131 20039 6137
rect 23290 6128 23296 6140
rect 23348 6128 23354 6180
rect 23477 6171 23535 6177
rect 23477 6137 23489 6171
rect 23523 6168 23535 6171
rect 23750 6168 23756 6180
rect 23523 6140 23756 6168
rect 23523 6137 23535 6140
rect 23477 6131 23535 6137
rect 23750 6128 23756 6140
rect 23808 6168 23814 6180
rect 24029 6171 24087 6177
rect 24029 6168 24041 6171
rect 23808 6140 24041 6168
rect 23808 6128 23814 6140
rect 24029 6137 24041 6140
rect 24075 6137 24087 6171
rect 24029 6131 24087 6137
rect 12897 6103 12955 6109
rect 12897 6100 12909 6103
rect 11848 6072 12909 6100
rect 11848 6060 11854 6072
rect 12897 6069 12909 6072
rect 12943 6069 12955 6103
rect 15470 6100 15476 6112
rect 15431 6072 15476 6100
rect 12897 6063 12955 6069
rect 15470 6060 15476 6072
rect 15528 6060 15534 6112
rect 17402 6100 17408 6112
rect 17363 6072 17408 6100
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 19426 6100 19432 6112
rect 19387 6072 19432 6100
rect 19426 6060 19432 6072
rect 19484 6060 19490 6112
rect 19518 6060 19524 6112
rect 19576 6100 19582 6112
rect 19613 6103 19671 6109
rect 19613 6100 19625 6103
rect 19576 6072 19625 6100
rect 19576 6060 19582 6072
rect 19613 6069 19625 6072
rect 19659 6069 19671 6103
rect 21174 6100 21180 6112
rect 21135 6072 21180 6100
rect 19613 6063 19671 6069
rect 21174 6060 21180 6072
rect 21232 6060 21238 6112
rect 21637 6103 21695 6109
rect 21637 6069 21649 6103
rect 21683 6100 21695 6103
rect 22462 6100 22468 6112
rect 21683 6072 22468 6100
rect 21683 6069 21695 6072
rect 21637 6063 21695 6069
rect 22462 6060 22468 6072
rect 22520 6060 22526 6112
rect 23658 6100 23664 6112
rect 23619 6072 23664 6100
rect 23658 6060 23664 6072
rect 23716 6060 23722 6112
rect 25409 6103 25467 6109
rect 25409 6069 25421 6103
rect 25455 6100 25467 6103
rect 25682 6100 25688 6112
rect 25455 6072 25688 6100
rect 25455 6069 25467 6072
rect 25409 6063 25467 6069
rect 25682 6060 25688 6072
rect 25740 6060 25746 6112
rect 26234 6100 26240 6112
rect 26195 6072 26240 6100
rect 26234 6060 26240 6072
rect 26292 6060 26298 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 2130 5856 2136 5908
rect 2188 5896 2194 5908
rect 2409 5899 2467 5905
rect 2409 5896 2421 5899
rect 2188 5868 2421 5896
rect 2188 5856 2194 5868
rect 2409 5865 2421 5868
rect 2455 5865 2467 5899
rect 2409 5859 2467 5865
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 2958 5896 2964 5908
rect 2915 5868 2964 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 2958 5856 2964 5868
rect 3016 5896 3022 5908
rect 3326 5896 3332 5908
rect 3016 5868 3332 5896
rect 3016 5856 3022 5868
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4249 5899 4307 5905
rect 4249 5896 4261 5899
rect 4028 5868 4261 5896
rect 4028 5856 4034 5868
rect 4249 5865 4261 5868
rect 4295 5865 4307 5899
rect 4614 5896 4620 5908
rect 4575 5868 4620 5896
rect 4249 5859 4307 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5350 5896 5356 5908
rect 5311 5868 5356 5896
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 5813 5899 5871 5905
rect 5813 5865 5825 5899
rect 5859 5896 5871 5899
rect 6086 5896 6092 5908
rect 5859 5868 6092 5896
rect 5859 5865 5871 5868
rect 5813 5859 5871 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 6825 5899 6883 5905
rect 6825 5865 6837 5899
rect 6871 5896 6883 5899
rect 7098 5896 7104 5908
rect 6871 5868 7104 5896
rect 6871 5865 6883 5868
rect 6825 5859 6883 5865
rect 7098 5856 7104 5868
rect 7156 5896 7162 5908
rect 8294 5896 8300 5908
rect 7156 5868 7420 5896
rect 8255 5868 8300 5896
rect 7156 5856 7162 5868
rect 1394 5788 1400 5840
rect 1452 5828 1458 5840
rect 5721 5831 5779 5837
rect 1452 5800 5672 5828
rect 1452 5788 1458 5800
rect 2777 5763 2835 5769
rect 2777 5729 2789 5763
rect 2823 5760 2835 5763
rect 3050 5760 3056 5772
rect 2823 5732 3056 5760
rect 2823 5729 2835 5732
rect 2777 5723 2835 5729
rect 3050 5720 3056 5732
rect 3108 5720 3114 5772
rect 3602 5720 3608 5772
rect 3660 5760 3666 5772
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 3660 5732 4077 5760
rect 3660 5720 3666 5732
rect 4065 5729 4077 5732
rect 4111 5729 4123 5763
rect 5644 5760 5672 5800
rect 5721 5797 5733 5831
rect 5767 5828 5779 5831
rect 6546 5828 6552 5840
rect 5767 5800 6552 5828
rect 5767 5797 5779 5800
rect 5721 5791 5779 5797
rect 6546 5788 6552 5800
rect 6604 5788 6610 5840
rect 6914 5788 6920 5840
rect 6972 5828 6978 5840
rect 7190 5837 7196 5840
rect 7184 5828 7196 5837
rect 6972 5800 7196 5828
rect 6972 5788 6978 5800
rect 7184 5791 7196 5800
rect 7190 5788 7196 5791
rect 7248 5788 7254 5840
rect 7392 5828 7420 5868
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 8846 5896 8852 5908
rect 8807 5868 8852 5896
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 11057 5899 11115 5905
rect 11057 5865 11069 5899
rect 11103 5896 11115 5899
rect 11146 5896 11152 5908
rect 11103 5868 11152 5896
rect 11103 5865 11115 5868
rect 11057 5859 11115 5865
rect 11146 5856 11152 5868
rect 11204 5856 11210 5908
rect 12621 5899 12679 5905
rect 12621 5865 12633 5899
rect 12667 5896 12679 5899
rect 12710 5896 12716 5908
rect 12667 5868 12716 5896
rect 12667 5865 12679 5868
rect 12621 5859 12679 5865
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 12802 5856 12808 5908
rect 12860 5896 12866 5908
rect 13354 5896 13360 5908
rect 12860 5868 13360 5896
rect 12860 5856 12866 5868
rect 13354 5856 13360 5868
rect 13412 5856 13418 5908
rect 14090 5896 14096 5908
rect 14051 5868 14096 5896
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 14274 5856 14280 5908
rect 14332 5896 14338 5908
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 14332 5868 14657 5896
rect 14332 5856 14338 5868
rect 14645 5865 14657 5868
rect 14691 5865 14703 5899
rect 15286 5896 15292 5908
rect 15247 5868 15292 5896
rect 14645 5859 14703 5865
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 15562 5856 15568 5908
rect 15620 5896 15626 5908
rect 15749 5899 15807 5905
rect 15749 5896 15761 5899
rect 15620 5868 15761 5896
rect 15620 5856 15626 5868
rect 15749 5865 15761 5868
rect 15795 5865 15807 5899
rect 16666 5896 16672 5908
rect 16627 5868 16672 5896
rect 15749 5859 15807 5865
rect 16666 5856 16672 5868
rect 16724 5856 16730 5908
rect 19150 5896 19156 5908
rect 19111 5868 19156 5896
rect 19150 5856 19156 5868
rect 19208 5856 19214 5908
rect 19518 5856 19524 5908
rect 19576 5896 19582 5908
rect 21358 5896 21364 5908
rect 19576 5868 21364 5896
rect 19576 5856 19582 5868
rect 21358 5856 21364 5868
rect 21416 5856 21422 5908
rect 21542 5856 21548 5908
rect 21600 5896 21606 5908
rect 21913 5899 21971 5905
rect 21913 5896 21925 5899
rect 21600 5868 21925 5896
rect 21600 5856 21606 5868
rect 21913 5865 21925 5868
rect 21959 5865 21971 5899
rect 22462 5896 22468 5908
rect 22375 5868 22468 5896
rect 21913 5859 21971 5865
rect 22462 5856 22468 5868
rect 22520 5856 22526 5908
rect 22922 5896 22928 5908
rect 22883 5868 22928 5896
rect 22922 5856 22928 5868
rect 22980 5856 22986 5908
rect 23658 5856 23664 5908
rect 23716 5896 23722 5908
rect 24397 5899 24455 5905
rect 24397 5896 24409 5899
rect 23716 5868 24409 5896
rect 23716 5856 23722 5868
rect 24397 5865 24409 5868
rect 24443 5896 24455 5899
rect 25041 5899 25099 5905
rect 25041 5896 25053 5899
rect 24443 5868 25053 5896
rect 24443 5865 24455 5868
rect 24397 5859 24455 5865
rect 25041 5865 25053 5868
rect 25087 5865 25099 5899
rect 25041 5859 25099 5865
rect 9950 5837 9956 5840
rect 9944 5828 9956 5837
rect 7392 5800 8340 5828
rect 9911 5800 9956 5828
rect 5644 5732 6040 5760
rect 4065 5723 4123 5729
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 3237 5695 3295 5701
rect 3237 5692 3249 5695
rect 3007 5664 3249 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 3237 5661 3249 5664
rect 3283 5661 3295 5695
rect 3510 5692 3516 5704
rect 3423 5664 3516 5692
rect 3237 5655 3295 5661
rect 3510 5652 3516 5664
rect 3568 5692 3574 5704
rect 5442 5692 5448 5704
rect 3568 5664 5448 5692
rect 3568 5652 3574 5664
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5661 5963 5695
rect 5905 5655 5963 5661
rect 2682 5584 2688 5636
rect 2740 5624 2746 5636
rect 4985 5627 5043 5633
rect 4985 5624 4997 5627
rect 2740 5596 4997 5624
rect 2740 5584 2746 5596
rect 4985 5593 4997 5596
rect 5031 5593 5043 5627
rect 4985 5587 5043 5593
rect 5350 5584 5356 5636
rect 5408 5624 5414 5636
rect 5534 5624 5540 5636
rect 5408 5596 5540 5624
rect 5408 5584 5414 5596
rect 5534 5584 5540 5596
rect 5592 5624 5598 5636
rect 5920 5624 5948 5655
rect 5592 5596 5948 5624
rect 6012 5624 6040 5732
rect 6086 5720 6092 5772
rect 6144 5760 6150 5772
rect 6822 5760 6828 5772
rect 6144 5732 6828 5760
rect 6144 5720 6150 5732
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 8312 5760 8340 5800
rect 9944 5791 9956 5800
rect 9950 5788 9956 5791
rect 10008 5788 10014 5840
rect 11882 5828 11888 5840
rect 11843 5800 11888 5828
rect 11882 5788 11888 5800
rect 11940 5788 11946 5840
rect 12253 5831 12311 5837
rect 12253 5797 12265 5831
rect 12299 5828 12311 5831
rect 14108 5828 14136 5856
rect 17126 5837 17132 5840
rect 17120 5828 17132 5837
rect 12299 5800 14136 5828
rect 17087 5800 17132 5828
rect 12299 5797 12311 5800
rect 12253 5791 12311 5797
rect 17120 5791 17132 5800
rect 17126 5788 17132 5791
rect 17184 5788 17190 5840
rect 19978 5828 19984 5840
rect 19939 5800 19984 5828
rect 19978 5788 19984 5800
rect 20036 5788 20042 5840
rect 21266 5828 21272 5840
rect 21227 5800 21272 5828
rect 21266 5788 21272 5800
rect 21324 5788 21330 5840
rect 22480 5828 22508 5856
rect 23566 5828 23572 5840
rect 22480 5800 23572 5828
rect 23566 5788 23572 5800
rect 23624 5788 23630 5840
rect 23753 5831 23811 5837
rect 23753 5797 23765 5831
rect 23799 5828 23811 5831
rect 24302 5828 24308 5840
rect 23799 5800 24308 5828
rect 23799 5797 23811 5800
rect 23753 5791 23811 5797
rect 24302 5788 24308 5800
rect 24360 5788 24366 5840
rect 26234 5828 26240 5840
rect 26195 5800 26240 5828
rect 26234 5788 26240 5800
rect 26292 5788 26298 5840
rect 11974 5760 11980 5772
rect 8312 5732 11980 5760
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 12986 5769 12992 5772
rect 12980 5760 12992 5769
rect 12947 5732 12992 5760
rect 12980 5723 12992 5732
rect 12986 5720 12992 5723
rect 13044 5720 13050 5772
rect 15470 5720 15476 5772
rect 15528 5760 15534 5772
rect 15657 5763 15715 5769
rect 15657 5760 15669 5763
rect 15528 5732 15669 5760
rect 15528 5720 15534 5732
rect 15657 5729 15669 5732
rect 15703 5729 15715 5763
rect 15657 5723 15715 5729
rect 16114 5720 16120 5772
rect 16172 5760 16178 5772
rect 16853 5763 16911 5769
rect 16853 5760 16865 5763
rect 16172 5732 16865 5760
rect 16172 5720 16178 5732
rect 16853 5729 16865 5732
rect 16899 5760 16911 5763
rect 17402 5760 17408 5772
rect 16899 5732 17408 5760
rect 16899 5729 16911 5732
rect 16853 5723 16911 5729
rect 17402 5720 17408 5732
rect 17460 5720 17466 5772
rect 19337 5763 19395 5769
rect 19337 5729 19349 5763
rect 19383 5760 19395 5763
rect 19518 5760 19524 5772
rect 19383 5732 19524 5760
rect 19383 5729 19395 5732
rect 19337 5723 19395 5729
rect 19518 5720 19524 5732
rect 19576 5720 19582 5772
rect 20254 5760 20260 5772
rect 20215 5732 20260 5760
rect 20254 5720 20260 5732
rect 20312 5760 20318 5772
rect 20312 5732 21496 5760
rect 20312 5720 20318 5732
rect 6546 5652 6552 5704
rect 6604 5692 6610 5704
rect 6917 5695 6975 5701
rect 6917 5692 6929 5695
rect 6604 5664 6929 5692
rect 6604 5652 6610 5664
rect 6917 5661 6929 5664
rect 6963 5661 6975 5695
rect 6917 5655 6975 5661
rect 9214 5652 9220 5704
rect 9272 5692 9278 5704
rect 9677 5695 9735 5701
rect 9677 5692 9689 5695
rect 9272 5664 9689 5692
rect 9272 5652 9278 5664
rect 9677 5661 9689 5664
rect 9723 5661 9735 5695
rect 9677 5655 9735 5661
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 12710 5692 12716 5704
rect 11848 5664 12716 5692
rect 11848 5652 11854 5664
rect 12710 5652 12716 5664
rect 12768 5652 12774 5704
rect 15286 5652 15292 5704
rect 15344 5692 15350 5704
rect 15841 5695 15899 5701
rect 15841 5692 15853 5695
rect 15344 5664 15853 5692
rect 15344 5652 15350 5664
rect 15841 5661 15853 5664
rect 15887 5692 15899 5695
rect 16022 5692 16028 5704
rect 15887 5664 16028 5692
rect 15887 5661 15899 5664
rect 15841 5655 15899 5661
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 21468 5701 21496 5732
rect 22738 5720 22744 5772
rect 22796 5760 22802 5772
rect 22833 5763 22891 5769
rect 22833 5760 22845 5763
rect 22796 5732 22845 5760
rect 22796 5720 22802 5732
rect 22833 5729 22845 5732
rect 22879 5729 22891 5763
rect 22833 5723 22891 5729
rect 23382 5720 23388 5772
rect 23440 5760 23446 5772
rect 24489 5763 24547 5769
rect 24489 5760 24501 5763
rect 23440 5732 24501 5760
rect 23440 5720 23446 5732
rect 24489 5729 24501 5732
rect 24535 5760 24547 5763
rect 25038 5760 25044 5772
rect 24535 5732 25044 5760
rect 24535 5729 24547 5732
rect 24489 5723 24547 5729
rect 25038 5720 25044 5732
rect 25096 5720 25102 5772
rect 25406 5720 25412 5772
rect 25464 5760 25470 5772
rect 25774 5760 25780 5772
rect 25464 5732 25780 5760
rect 25464 5720 25470 5732
rect 25774 5720 25780 5732
rect 25832 5720 25838 5772
rect 21453 5695 21511 5701
rect 21453 5661 21465 5695
rect 21499 5692 21511 5695
rect 21726 5692 21732 5704
rect 21499 5664 21732 5692
rect 21499 5661 21511 5664
rect 21453 5655 21511 5661
rect 21726 5652 21732 5664
rect 21784 5652 21790 5704
rect 23014 5692 23020 5704
rect 22975 5664 23020 5692
rect 23014 5652 23020 5664
rect 23072 5652 23078 5704
rect 23934 5692 23940 5704
rect 23308 5664 23940 5692
rect 9122 5624 9128 5636
rect 6012 5596 6960 5624
rect 9035 5596 9128 5624
rect 5592 5584 5598 5596
rect 1762 5556 1768 5568
rect 1723 5528 1768 5556
rect 1762 5516 1768 5528
rect 1820 5516 1826 5568
rect 1854 5516 1860 5568
rect 1912 5556 1918 5568
rect 2225 5559 2283 5565
rect 2225 5556 2237 5559
rect 1912 5528 2237 5556
rect 1912 5516 1918 5528
rect 2225 5525 2237 5528
rect 2271 5525 2283 5559
rect 2225 5519 2283 5525
rect 3237 5559 3295 5565
rect 3237 5525 3249 5559
rect 3283 5556 3295 5559
rect 3881 5559 3939 5565
rect 3881 5556 3893 5559
rect 3283 5528 3893 5556
rect 3283 5525 3295 5528
rect 3237 5519 3295 5525
rect 3881 5525 3893 5528
rect 3927 5556 3939 5559
rect 3970 5556 3976 5568
rect 3927 5528 3976 5556
rect 3927 5525 3939 5528
rect 3881 5519 3939 5525
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 6362 5556 6368 5568
rect 6323 5528 6368 5556
rect 6362 5516 6368 5528
rect 6420 5516 6426 5568
rect 6932 5556 6960 5596
rect 9048 5556 9076 5596
rect 9122 5584 9128 5596
rect 9180 5624 9186 5636
rect 9180 5596 9352 5624
rect 9180 5584 9186 5596
rect 9214 5556 9220 5568
rect 6932 5528 9076 5556
rect 9175 5528 9220 5556
rect 9214 5516 9220 5528
rect 9272 5516 9278 5568
rect 9324 5556 9352 5596
rect 13814 5584 13820 5636
rect 13872 5624 13878 5636
rect 15013 5627 15071 5633
rect 15013 5624 15025 5627
rect 13872 5596 15025 5624
rect 13872 5584 13878 5596
rect 15013 5593 15025 5596
rect 15059 5624 15071 5627
rect 15378 5624 15384 5636
rect 15059 5596 15384 5624
rect 15059 5593 15071 5596
rect 15013 5587 15071 5593
rect 15378 5584 15384 5596
rect 15436 5584 15442 5636
rect 18230 5624 18236 5636
rect 18191 5596 18236 5624
rect 18230 5584 18236 5596
rect 18288 5584 18294 5636
rect 20901 5627 20959 5633
rect 20901 5593 20913 5627
rect 20947 5624 20959 5627
rect 21542 5624 21548 5636
rect 20947 5596 21548 5624
rect 20947 5593 20959 5596
rect 20901 5587 20959 5593
rect 21542 5584 21548 5596
rect 21600 5624 21606 5636
rect 22002 5624 22008 5636
rect 21600 5596 22008 5624
rect 21600 5584 21606 5596
rect 22002 5584 22008 5596
rect 22060 5584 22066 5636
rect 22373 5627 22431 5633
rect 22373 5593 22385 5627
rect 22419 5624 22431 5627
rect 23308 5624 23336 5664
rect 23934 5652 23940 5664
rect 23992 5652 23998 5704
rect 24578 5652 24584 5704
rect 24636 5692 24642 5704
rect 24762 5692 24768 5704
rect 24636 5664 24768 5692
rect 24636 5652 24642 5664
rect 24762 5652 24768 5664
rect 24820 5652 24826 5704
rect 22419 5596 23336 5624
rect 22419 5593 22431 5596
rect 22373 5587 22431 5593
rect 18046 5556 18052 5568
rect 9324 5528 18052 5556
rect 18046 5516 18052 5528
rect 18104 5516 18110 5568
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 19521 5559 19579 5565
rect 19521 5556 19533 5559
rect 19392 5528 19533 5556
rect 19392 5516 19398 5528
rect 19521 5525 19533 5528
rect 19567 5525 19579 5559
rect 19521 5519 19579 5525
rect 20717 5559 20775 5565
rect 20717 5525 20729 5559
rect 20763 5556 20775 5559
rect 21450 5556 21456 5568
rect 20763 5528 21456 5556
rect 20763 5525 20775 5528
rect 20717 5519 20775 5525
rect 21450 5516 21456 5528
rect 21508 5516 21514 5568
rect 21818 5516 21824 5568
rect 21876 5556 21882 5568
rect 22388 5556 22416 5587
rect 23474 5584 23480 5636
rect 23532 5624 23538 5636
rect 24029 5627 24087 5633
rect 24029 5624 24041 5627
rect 23532 5596 24041 5624
rect 23532 5584 23538 5596
rect 24029 5593 24041 5596
rect 24075 5593 24087 5627
rect 24029 5587 24087 5593
rect 24946 5584 24952 5636
rect 25004 5624 25010 5636
rect 25777 5627 25835 5633
rect 25777 5624 25789 5627
rect 25004 5596 25789 5624
rect 25004 5584 25010 5596
rect 25777 5593 25789 5596
rect 25823 5593 25835 5627
rect 25777 5587 25835 5593
rect 25406 5556 25412 5568
rect 21876 5528 22416 5556
rect 25367 5528 25412 5556
rect 21876 5516 21882 5528
rect 25406 5516 25412 5528
rect 25464 5516 25470 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 2777 5355 2835 5361
rect 2777 5321 2789 5355
rect 2823 5352 2835 5355
rect 2958 5352 2964 5364
rect 2823 5324 2964 5352
rect 2823 5321 2835 5324
rect 2777 5315 2835 5321
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 3145 5355 3203 5361
rect 3145 5321 3157 5355
rect 3191 5352 3203 5355
rect 3234 5352 3240 5364
rect 3191 5324 3240 5352
rect 3191 5321 3203 5324
rect 3145 5315 3203 5321
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 6273 5355 6331 5361
rect 6273 5321 6285 5355
rect 6319 5352 6331 5355
rect 6822 5352 6828 5364
rect 6319 5324 6828 5352
rect 6319 5321 6331 5324
rect 6273 5315 6331 5321
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 7101 5355 7159 5361
rect 7101 5352 7113 5355
rect 7064 5324 7113 5352
rect 7064 5312 7070 5324
rect 7101 5321 7113 5324
rect 7147 5321 7159 5355
rect 7101 5315 7159 5321
rect 7561 5355 7619 5361
rect 7561 5321 7573 5355
rect 7607 5352 7619 5355
rect 7834 5352 7840 5364
rect 7607 5324 7840 5352
rect 7607 5321 7619 5324
rect 7561 5315 7619 5321
rect 1673 5287 1731 5293
rect 1673 5253 1685 5287
rect 1719 5284 1731 5287
rect 2130 5284 2136 5296
rect 1719 5256 2136 5284
rect 1719 5253 1731 5256
rect 1673 5247 1731 5253
rect 2130 5244 2136 5256
rect 2188 5284 2194 5296
rect 2682 5284 2688 5296
rect 2188 5256 2688 5284
rect 2188 5244 2194 5256
rect 2682 5244 2688 5256
rect 2740 5244 2746 5296
rect 1762 5176 1768 5228
rect 1820 5216 1826 5228
rect 2225 5219 2283 5225
rect 2225 5216 2237 5219
rect 1820 5188 2237 5216
rect 1820 5176 1826 5188
rect 2225 5185 2237 5188
rect 2271 5216 2283 5219
rect 5718 5216 5724 5228
rect 2271 5188 3372 5216
rect 5679 5188 5724 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 2038 5148 2044 5160
rect 1999 5120 2044 5148
rect 2038 5108 2044 5120
rect 2096 5108 2102 5160
rect 2133 5151 2191 5157
rect 2133 5117 2145 5151
rect 2179 5148 2191 5151
rect 2498 5148 2504 5160
rect 2179 5120 2504 5148
rect 2179 5117 2191 5120
rect 2133 5111 2191 5117
rect 2498 5108 2504 5120
rect 2556 5108 2562 5160
rect 3234 5148 3240 5160
rect 3195 5120 3240 5148
rect 3234 5108 3240 5120
rect 3292 5108 3298 5160
rect 3344 5148 3372 5188
rect 5718 5176 5724 5188
rect 5776 5176 5782 5228
rect 3510 5157 3516 5160
rect 3504 5148 3516 5157
rect 3344 5120 3516 5148
rect 3504 5111 3516 5120
rect 3510 5108 3516 5111
rect 3568 5108 3574 5160
rect 7116 5148 7144 5315
rect 7834 5312 7840 5324
rect 7892 5352 7898 5364
rect 8662 5352 8668 5364
rect 7892 5324 8156 5352
rect 8623 5324 8668 5352
rect 7892 5312 7898 5324
rect 7653 5287 7711 5293
rect 7653 5253 7665 5287
rect 7699 5284 7711 5287
rect 7926 5284 7932 5296
rect 7699 5256 7932 5284
rect 7699 5253 7711 5256
rect 7653 5247 7711 5253
rect 7926 5244 7932 5256
rect 7984 5244 7990 5296
rect 8128 5225 8156 5324
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 10502 5352 10508 5364
rect 10463 5324 10508 5352
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 12437 5355 12495 5361
rect 12437 5321 12449 5355
rect 12483 5352 12495 5355
rect 12618 5352 12624 5364
rect 12483 5324 12624 5352
rect 12483 5321 12495 5324
rect 12437 5315 12495 5321
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 13906 5352 13912 5364
rect 13867 5324 13912 5352
rect 13906 5312 13912 5324
rect 13964 5312 13970 5364
rect 15013 5355 15071 5361
rect 15013 5321 15025 5355
rect 15059 5352 15071 5355
rect 15286 5352 15292 5364
rect 15059 5324 15292 5352
rect 15059 5321 15071 5324
rect 15013 5315 15071 5321
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 16577 5355 16635 5361
rect 16577 5321 16589 5355
rect 16623 5352 16635 5355
rect 17126 5352 17132 5364
rect 16623 5324 17132 5352
rect 16623 5321 16635 5324
rect 16577 5315 16635 5321
rect 17126 5312 17132 5324
rect 17184 5312 17190 5364
rect 17497 5355 17555 5361
rect 17497 5321 17509 5355
rect 17543 5352 17555 5355
rect 17678 5352 17684 5364
rect 17543 5324 17684 5352
rect 17543 5321 17555 5324
rect 17497 5315 17555 5321
rect 17678 5312 17684 5324
rect 17736 5352 17742 5364
rect 19337 5355 19395 5361
rect 19337 5352 19349 5355
rect 17736 5324 19349 5352
rect 17736 5312 17742 5324
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5216 8355 5219
rect 8680 5216 8708 5312
rect 16114 5244 16120 5296
rect 16172 5284 16178 5296
rect 16853 5287 16911 5293
rect 16853 5284 16865 5287
rect 16172 5256 16865 5284
rect 16172 5244 16178 5256
rect 16853 5253 16865 5256
rect 16899 5253 16911 5287
rect 16853 5247 16911 5253
rect 17865 5287 17923 5293
rect 17865 5253 17877 5287
rect 17911 5284 17923 5287
rect 18322 5284 18328 5296
rect 17911 5256 18328 5284
rect 17911 5253 17923 5256
rect 17865 5247 17923 5253
rect 18322 5244 18328 5256
rect 18380 5244 18386 5296
rect 8343 5188 8708 5216
rect 10045 5219 10103 5225
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 10045 5185 10057 5219
rect 10091 5216 10103 5219
rect 10870 5216 10876 5228
rect 10091 5188 10876 5216
rect 10091 5185 10103 5188
rect 10045 5179 10103 5185
rect 10870 5176 10876 5188
rect 10928 5176 10934 5228
rect 11146 5216 11152 5228
rect 11107 5188 11152 5216
rect 11146 5176 11152 5188
rect 11204 5216 11210 5228
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 11204 5188 11529 5216
rect 11204 5176 11210 5188
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5216 12311 5219
rect 12989 5219 13047 5225
rect 12989 5216 13001 5219
rect 12299 5188 13001 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 12989 5185 13001 5188
rect 13035 5216 13047 5219
rect 13446 5216 13452 5228
rect 13035 5188 13452 5216
rect 13035 5185 13047 5188
rect 12989 5179 13047 5185
rect 13446 5176 13452 5188
rect 13504 5176 13510 5228
rect 16022 5216 16028 5228
rect 15983 5188 16028 5216
rect 16022 5176 16028 5188
rect 16080 5176 16086 5228
rect 18524 5225 18552 5324
rect 19337 5321 19349 5324
rect 19383 5352 19395 5355
rect 19518 5352 19524 5364
rect 19383 5324 19524 5352
rect 19383 5321 19395 5324
rect 19337 5315 19395 5321
rect 19518 5312 19524 5324
rect 19576 5312 19582 5364
rect 19978 5312 19984 5364
rect 20036 5352 20042 5364
rect 20530 5352 20536 5364
rect 20036 5324 20536 5352
rect 20036 5312 20042 5324
rect 20530 5312 20536 5324
rect 20588 5352 20594 5364
rect 20625 5355 20683 5361
rect 20625 5352 20637 5355
rect 20588 5324 20637 5352
rect 20588 5312 20594 5324
rect 20625 5321 20637 5324
rect 20671 5321 20683 5355
rect 20990 5352 20996 5364
rect 20951 5324 20996 5352
rect 20625 5315 20683 5321
rect 20990 5312 20996 5324
rect 21048 5352 21054 5364
rect 22557 5355 22615 5361
rect 21048 5324 21772 5352
rect 21048 5312 21054 5324
rect 19613 5287 19671 5293
rect 19613 5253 19625 5287
rect 19659 5284 19671 5287
rect 19659 5256 21680 5284
rect 19659 5253 19671 5256
rect 19613 5247 19671 5253
rect 21652 5228 21680 5256
rect 18509 5219 18567 5225
rect 18509 5185 18521 5219
rect 18555 5185 18567 5219
rect 18509 5179 18567 5185
rect 18601 5219 18659 5225
rect 18601 5185 18613 5219
rect 18647 5185 18659 5219
rect 20162 5216 20168 5228
rect 20123 5188 20168 5216
rect 18601 5179 18659 5185
rect 8018 5148 8024 5160
rect 7116 5120 8024 5148
rect 8018 5108 8024 5120
rect 8076 5108 8082 5160
rect 10888 5148 10916 5176
rect 11882 5148 11888 5160
rect 10888 5120 11888 5148
rect 10318 5040 10324 5092
rect 10376 5080 10382 5092
rect 10888 5089 10916 5120
rect 11882 5108 11888 5120
rect 11940 5108 11946 5160
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5148 12955 5151
rect 13722 5148 13728 5160
rect 12943 5120 13728 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 13722 5108 13728 5120
rect 13780 5108 13786 5160
rect 14274 5108 14280 5160
rect 14332 5148 14338 5160
rect 14369 5151 14427 5157
rect 14369 5148 14381 5151
rect 14332 5120 14381 5148
rect 14332 5108 14338 5120
rect 14369 5117 14381 5120
rect 14415 5117 14427 5151
rect 14369 5111 14427 5117
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 15841 5151 15899 5157
rect 15841 5148 15853 5151
rect 15436 5120 15853 5148
rect 15436 5108 15442 5120
rect 15841 5117 15853 5120
rect 15887 5117 15899 5151
rect 15841 5111 15899 5117
rect 18414 5108 18420 5160
rect 18472 5148 18478 5160
rect 18616 5148 18644 5179
rect 20162 5176 20168 5188
rect 20220 5176 20226 5228
rect 21634 5216 21640 5228
rect 21547 5188 21640 5216
rect 21634 5176 21640 5188
rect 21692 5176 21698 5228
rect 21744 5225 21772 5324
rect 22557 5321 22569 5355
rect 22603 5352 22615 5355
rect 22738 5352 22744 5364
rect 22603 5324 22744 5352
rect 22603 5321 22615 5324
rect 22557 5315 22615 5321
rect 22738 5312 22744 5324
rect 22796 5312 22802 5364
rect 22922 5352 22928 5364
rect 22883 5324 22928 5352
rect 22922 5312 22928 5324
rect 22980 5312 22986 5364
rect 23658 5352 23664 5364
rect 23619 5324 23664 5352
rect 23658 5312 23664 5324
rect 23716 5312 23722 5364
rect 24762 5352 24768 5364
rect 24723 5324 24768 5352
rect 24762 5312 24768 5324
rect 24820 5312 24826 5364
rect 25038 5352 25044 5364
rect 24999 5324 25044 5352
rect 25038 5312 25044 5324
rect 25096 5312 25102 5364
rect 25866 5352 25872 5364
rect 25827 5324 25872 5352
rect 25866 5312 25872 5324
rect 25924 5312 25930 5364
rect 22186 5244 22192 5296
rect 22244 5284 22250 5296
rect 25222 5284 25228 5296
rect 22244 5256 25228 5284
rect 22244 5244 22250 5256
rect 25222 5244 25228 5256
rect 25280 5244 25286 5296
rect 21729 5219 21787 5225
rect 21729 5185 21741 5219
rect 21775 5185 21787 5219
rect 21729 5179 21787 5185
rect 22094 5176 22100 5228
rect 22152 5216 22158 5228
rect 23385 5219 23443 5225
rect 23385 5216 23397 5219
rect 22152 5188 23397 5216
rect 22152 5176 22158 5188
rect 23385 5185 23397 5188
rect 23431 5216 23443 5219
rect 23431 5188 23888 5216
rect 23431 5185 23443 5188
rect 23385 5179 23443 5185
rect 18472 5120 18644 5148
rect 18472 5108 18478 5120
rect 19058 5108 19064 5160
rect 19116 5148 19122 5160
rect 20073 5151 20131 5157
rect 20073 5148 20085 5151
rect 19116 5120 20085 5148
rect 19116 5108 19122 5120
rect 20073 5117 20085 5120
rect 20119 5148 20131 5151
rect 21542 5148 21548 5160
rect 20119 5120 21404 5148
rect 21503 5120 21548 5148
rect 20119 5117 20131 5120
rect 20073 5111 20131 5117
rect 10873 5083 10931 5089
rect 10376 5052 10456 5080
rect 10376 5040 10382 5052
rect 4614 5012 4620 5024
rect 4575 4984 4620 5012
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 5261 5015 5319 5021
rect 5261 4981 5273 5015
rect 5307 5012 5319 5015
rect 5350 5012 5356 5024
rect 5307 4984 5356 5012
rect 5307 4981 5319 4984
rect 5261 4975 5319 4981
rect 5350 4972 5356 4984
rect 5408 5012 5414 5024
rect 5537 5015 5595 5021
rect 5537 5012 5549 5015
rect 5408 4984 5549 5012
rect 5408 4972 5414 4984
rect 5537 4981 5549 4984
rect 5583 4981 5595 5015
rect 6546 5012 6552 5024
rect 6507 4984 6552 5012
rect 5537 4975 5595 4981
rect 6546 4972 6552 4984
rect 6604 5012 6610 5024
rect 7742 5012 7748 5024
rect 6604 4984 7748 5012
rect 6604 4972 6610 4984
rect 7742 4972 7748 4984
rect 7800 5012 7806 5024
rect 9309 5015 9367 5021
rect 9309 5012 9321 5015
rect 7800 4984 9321 5012
rect 7800 4972 7806 4984
rect 9309 4981 9321 4984
rect 9355 4981 9367 5015
rect 9490 5012 9496 5024
rect 9451 4984 9496 5012
rect 9309 4975 9367 4981
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 10428 5021 10456 5052
rect 10873 5049 10885 5083
rect 10919 5049 10931 5083
rect 10873 5043 10931 5049
rect 11514 5040 11520 5092
rect 11572 5080 11578 5092
rect 12805 5083 12863 5089
rect 12805 5080 12817 5083
rect 11572 5052 12817 5080
rect 11572 5040 11578 5052
rect 12805 5049 12817 5052
rect 12851 5049 12863 5083
rect 12805 5043 12863 5049
rect 15102 5040 15108 5092
rect 15160 5080 15166 5092
rect 15933 5083 15991 5089
rect 15933 5080 15945 5083
rect 15160 5052 15945 5080
rect 15160 5040 15166 5052
rect 15933 5049 15945 5052
rect 15979 5080 15991 5083
rect 19981 5083 20039 5089
rect 15979 5052 18092 5080
rect 15979 5049 15991 5052
rect 15933 5043 15991 5049
rect 10413 5015 10471 5021
rect 10413 4981 10425 5015
rect 10459 5012 10471 5015
rect 10965 5015 11023 5021
rect 10965 5012 10977 5015
rect 10459 4984 10977 5012
rect 10459 4981 10471 4984
rect 10413 4975 10471 4981
rect 10965 4981 10977 4984
rect 11011 5012 11023 5015
rect 11330 5012 11336 5024
rect 11011 4984 11336 5012
rect 11011 4981 11023 4984
rect 10965 4975 11023 4981
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 12710 4972 12716 5024
rect 12768 5012 12774 5024
rect 12986 5012 12992 5024
rect 12768 4984 12992 5012
rect 12768 4972 12774 4984
rect 12986 4972 12992 4984
rect 13044 5012 13050 5024
rect 13449 5015 13507 5021
rect 13449 5012 13461 5015
rect 13044 4984 13461 5012
rect 13044 4972 13050 4984
rect 13449 4981 13461 4984
rect 13495 4981 13507 5015
rect 13449 4975 13507 4981
rect 13998 4972 14004 5024
rect 14056 5012 14062 5024
rect 14185 5015 14243 5021
rect 14185 5012 14197 5015
rect 14056 4984 14197 5012
rect 14056 4972 14062 4984
rect 14185 4981 14197 4984
rect 14231 4981 14243 5015
rect 14550 5012 14556 5024
rect 14511 4984 14556 5012
rect 14185 4975 14243 4981
rect 14550 4972 14556 4984
rect 14608 4972 14614 5024
rect 15378 5012 15384 5024
rect 15339 4984 15384 5012
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 15473 5015 15531 5021
rect 15473 4981 15485 5015
rect 15519 5012 15531 5015
rect 16482 5012 16488 5024
rect 15519 4984 16488 5012
rect 15519 4981 15531 4984
rect 15473 4975 15531 4981
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 18064 5021 18092 5052
rect 19981 5049 19993 5083
rect 20027 5080 20039 5083
rect 20162 5080 20168 5092
rect 20027 5052 20168 5080
rect 20027 5049 20039 5052
rect 19981 5043 20039 5049
rect 20162 5040 20168 5052
rect 20220 5040 20226 5092
rect 18049 5015 18107 5021
rect 18049 4981 18061 5015
rect 18095 4981 18107 5015
rect 18049 4975 18107 4981
rect 18322 4972 18328 5024
rect 18380 5012 18386 5024
rect 18417 5015 18475 5021
rect 18417 5012 18429 5015
rect 18380 4984 18429 5012
rect 18380 4972 18386 4984
rect 18417 4981 18429 4984
rect 18463 4981 18475 5015
rect 21174 5012 21180 5024
rect 21135 4984 21180 5012
rect 18417 4975 18475 4981
rect 21174 4972 21180 4984
rect 21232 4972 21238 5024
rect 21376 5012 21404 5120
rect 21542 5108 21548 5120
rect 21600 5108 21606 5160
rect 23032 5120 23796 5148
rect 21450 5040 21456 5092
rect 21508 5080 21514 5092
rect 22646 5080 22652 5092
rect 21508 5052 22652 5080
rect 21508 5040 21514 5052
rect 22646 5040 22652 5052
rect 22704 5040 22710 5092
rect 23032 5012 23060 5120
rect 21376 4984 23060 5012
rect 23768 5012 23796 5120
rect 23860 5080 23888 5188
rect 23934 5176 23940 5228
rect 23992 5216 23998 5228
rect 24302 5216 24308 5228
rect 23992 5188 24308 5216
rect 23992 5176 23998 5188
rect 24302 5176 24308 5188
rect 24360 5176 24366 5228
rect 24026 5148 24032 5160
rect 23987 5120 24032 5148
rect 24026 5108 24032 5120
rect 24084 5108 24090 5160
rect 25225 5151 25283 5157
rect 25225 5117 25237 5151
rect 25271 5148 25283 5151
rect 25866 5148 25872 5160
rect 25271 5120 25872 5148
rect 25271 5117 25283 5120
rect 25225 5111 25283 5117
rect 25866 5108 25872 5120
rect 25924 5108 25930 5160
rect 24121 5083 24179 5089
rect 24121 5080 24133 5083
rect 23860 5052 24133 5080
rect 24121 5049 24133 5052
rect 24167 5049 24179 5083
rect 26145 5083 26203 5089
rect 26145 5080 26157 5083
rect 24121 5043 24179 5049
rect 24228 5052 26157 5080
rect 24228 5012 24256 5052
rect 26145 5049 26157 5052
rect 26191 5049 26203 5083
rect 26145 5043 26203 5049
rect 23768 4984 24256 5012
rect 25222 4972 25228 5024
rect 25280 5012 25286 5024
rect 25409 5015 25467 5021
rect 25409 5012 25421 5015
rect 25280 4984 25421 5012
rect 25280 4972 25286 4984
rect 25409 4981 25421 4984
rect 25455 4981 25467 5015
rect 25409 4975 25467 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 2314 4808 2320 4820
rect 2275 4780 2320 4808
rect 2314 4768 2320 4780
rect 2372 4768 2378 4820
rect 2409 4811 2467 4817
rect 2409 4777 2421 4811
rect 2455 4808 2467 4811
rect 2682 4808 2688 4820
rect 2455 4780 2688 4808
rect 2455 4777 2467 4780
rect 2409 4771 2467 4777
rect 2682 4768 2688 4780
rect 2740 4768 2746 4820
rect 2777 4811 2835 4817
rect 2777 4777 2789 4811
rect 2823 4808 2835 4811
rect 4062 4808 4068 4820
rect 2823 4780 4068 4808
rect 2823 4777 2835 4780
rect 2777 4771 2835 4777
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 4798 4768 4804 4820
rect 4856 4808 4862 4820
rect 8938 4808 8944 4820
rect 4856 4780 8944 4808
rect 4856 4768 4862 4780
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 10413 4811 10471 4817
rect 10413 4808 10425 4811
rect 9732 4780 10425 4808
rect 9732 4768 9738 4780
rect 10413 4777 10425 4780
rect 10459 4777 10471 4811
rect 10870 4808 10876 4820
rect 10831 4780 10876 4808
rect 10413 4771 10471 4777
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 11514 4808 11520 4820
rect 11475 4780 11520 4808
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 13633 4811 13691 4817
rect 13633 4777 13645 4811
rect 13679 4808 13691 4811
rect 13814 4808 13820 4820
rect 13679 4780 13820 4808
rect 13679 4777 13691 4780
rect 13633 4771 13691 4777
rect 13814 4768 13820 4780
rect 13872 4768 13878 4820
rect 14001 4811 14059 4817
rect 14001 4777 14013 4811
rect 14047 4808 14059 4811
rect 14366 4808 14372 4820
rect 14047 4780 14372 4808
rect 14047 4777 14059 4780
rect 14001 4771 14059 4777
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 15102 4808 15108 4820
rect 15063 4780 15108 4808
rect 15102 4768 15108 4780
rect 15160 4768 15166 4820
rect 18141 4811 18199 4817
rect 18141 4777 18153 4811
rect 18187 4808 18199 4811
rect 18874 4808 18880 4820
rect 18187 4780 18880 4808
rect 18187 4777 18199 4780
rect 18141 4771 18199 4777
rect 18874 4768 18880 4780
rect 18932 4768 18938 4820
rect 20714 4808 20720 4820
rect 20675 4780 20720 4808
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 21726 4768 21732 4820
rect 21784 4808 21790 4820
rect 21913 4811 21971 4817
rect 21913 4808 21925 4811
rect 21784 4780 21925 4808
rect 21784 4768 21790 4780
rect 21913 4777 21925 4780
rect 21959 4777 21971 4811
rect 21913 4771 21971 4777
rect 22373 4811 22431 4817
rect 22373 4777 22385 4811
rect 22419 4808 22431 4811
rect 23014 4808 23020 4820
rect 22419 4780 23020 4808
rect 22419 4777 22431 4780
rect 22373 4771 22431 4777
rect 23014 4768 23020 4780
rect 23072 4768 23078 4820
rect 23753 4811 23811 4817
rect 23753 4777 23765 4811
rect 23799 4808 23811 4811
rect 24026 4808 24032 4820
rect 23799 4780 24032 4808
rect 23799 4777 23811 4780
rect 23753 4771 23811 4777
rect 24026 4768 24032 4780
rect 24084 4768 24090 4820
rect 24121 4811 24179 4817
rect 24121 4777 24133 4811
rect 24167 4808 24179 4811
rect 24302 4808 24308 4820
rect 24167 4780 24308 4808
rect 24167 4777 24179 4780
rect 24121 4771 24179 4777
rect 24302 4768 24308 4780
rect 24360 4768 24366 4820
rect 3881 4743 3939 4749
rect 3881 4740 3893 4743
rect 2332 4712 3893 4740
rect 2332 4684 2360 4712
rect 3881 4709 3893 4712
rect 3927 4740 3939 4743
rect 4332 4743 4390 4749
rect 4332 4740 4344 4743
rect 3927 4712 4344 4740
rect 3927 4709 3939 4712
rect 3881 4703 3939 4709
rect 4332 4709 4344 4712
rect 4378 4740 4390 4743
rect 4614 4740 4620 4752
rect 4378 4712 4620 4740
rect 4378 4709 4390 4712
rect 4332 4703 4390 4709
rect 4614 4700 4620 4712
rect 4672 4700 4678 4752
rect 5994 4700 6000 4752
rect 6052 4740 6058 4752
rect 6089 4743 6147 4749
rect 6089 4740 6101 4743
rect 6052 4712 6101 4740
rect 6052 4700 6058 4712
rect 6089 4709 6101 4712
rect 6135 4740 6147 4743
rect 8294 4740 8300 4752
rect 6135 4712 8300 4740
rect 6135 4709 6147 4712
rect 6089 4703 6147 4709
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 9950 4740 9956 4752
rect 9911 4712 9956 4740
rect 9950 4700 9956 4712
rect 10008 4700 10014 4752
rect 13170 4740 13176 4752
rect 13083 4712 13176 4740
rect 13170 4700 13176 4712
rect 13228 4740 13234 4752
rect 17862 4740 17868 4752
rect 13228 4712 17868 4740
rect 13228 4700 13234 4712
rect 17862 4700 17868 4712
rect 17920 4700 17926 4752
rect 18598 4700 18604 4752
rect 18656 4740 18662 4752
rect 19061 4743 19119 4749
rect 19061 4740 19073 4743
rect 18656 4712 19073 4740
rect 18656 4700 18662 4712
rect 19061 4709 19073 4712
rect 19107 4709 19119 4743
rect 20732 4740 20760 4768
rect 22925 4743 22983 4749
rect 20732 4712 21496 4740
rect 19061 4703 19119 4709
rect 2314 4632 2320 4684
rect 2372 4632 2378 4684
rect 2869 4675 2927 4681
rect 2869 4641 2881 4675
rect 2915 4672 2927 4675
rect 3418 4672 3424 4684
rect 2915 4644 3424 4672
rect 2915 4641 2927 4644
rect 2869 4635 2927 4641
rect 3418 4632 3424 4644
rect 3476 4632 3482 4684
rect 6805 4675 6863 4681
rect 6805 4672 6817 4675
rect 6380 4644 6817 4672
rect 2958 4564 2964 4616
rect 3016 4604 3022 4616
rect 3053 4607 3111 4613
rect 3053 4604 3065 4607
rect 3016 4576 3065 4604
rect 3016 4564 3022 4576
rect 3053 4573 3065 4576
rect 3099 4604 3111 4607
rect 3510 4604 3516 4616
rect 3099 4576 3516 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 3510 4564 3516 4576
rect 3568 4564 3574 4616
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 3234 4496 3240 4548
rect 3292 4536 3298 4548
rect 4080 4536 4108 4567
rect 6380 4545 6408 4644
rect 6805 4641 6817 4644
rect 6851 4641 6863 4675
rect 10778 4672 10784 4684
rect 10739 4644 10784 4672
rect 6805 4635 6863 4641
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 12434 4632 12440 4684
rect 12492 4672 12498 4684
rect 13541 4675 13599 4681
rect 12492 4644 12537 4672
rect 12492 4632 12498 4644
rect 13541 4641 13553 4675
rect 13587 4672 13599 4675
rect 13722 4672 13728 4684
rect 13587 4644 13728 4672
rect 13587 4641 13599 4644
rect 13541 4635 13599 4641
rect 6546 4604 6552 4616
rect 6507 4576 6552 4604
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 11057 4607 11115 4613
rect 11057 4573 11069 4607
rect 11103 4604 11115 4607
rect 11146 4604 11152 4616
rect 11103 4576 11152 4604
rect 11103 4573 11115 4576
rect 11057 4567 11115 4573
rect 11146 4564 11152 4576
rect 11204 4564 11210 4616
rect 12526 4604 12532 4616
rect 12487 4576 12532 4604
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 12713 4607 12771 4613
rect 12713 4573 12725 4607
rect 12759 4604 12771 4607
rect 13556 4604 13584 4635
rect 13722 4632 13728 4644
rect 13780 4672 13786 4684
rect 16384 4675 16442 4681
rect 16384 4672 16396 4675
rect 13780 4644 16396 4672
rect 13780 4632 13786 4644
rect 14090 4604 14096 4616
rect 12759 4576 13584 4604
rect 14051 4576 14096 4604
rect 12759 4573 12771 4576
rect 12713 4567 12771 4573
rect 6365 4539 6423 4545
rect 6365 4536 6377 4539
rect 3292 4508 4108 4536
rect 5460 4508 6377 4536
rect 3292 4496 3298 4508
rect 1949 4471 2007 4477
rect 1949 4437 1961 4471
rect 1995 4468 2007 4471
rect 3513 4471 3571 4477
rect 3513 4468 3525 4471
rect 1995 4440 3525 4468
rect 1995 4437 2007 4440
rect 1949 4431 2007 4437
rect 3513 4437 3525 4440
rect 3559 4468 3571 4471
rect 3970 4468 3976 4480
rect 3559 4440 3976 4468
rect 3559 4437 3571 4440
rect 3513 4431 3571 4437
rect 3970 4428 3976 4440
rect 4028 4428 4034 4480
rect 4246 4428 4252 4480
rect 4304 4468 4310 4480
rect 5460 4477 5488 4508
rect 6365 4505 6377 4508
rect 6411 4505 6423 4539
rect 6365 4499 6423 4505
rect 11977 4539 12035 4545
rect 11977 4505 11989 4539
rect 12023 4536 12035 4539
rect 12728 4536 12756 4567
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 14292 4613 14320 4644
rect 16384 4641 16396 4644
rect 16430 4672 16442 4675
rect 17218 4672 17224 4684
rect 16430 4644 17224 4672
rect 16430 4641 16442 4644
rect 16384 4635 16442 4641
rect 17218 4632 17224 4644
rect 17276 4672 17282 4684
rect 18414 4672 18420 4684
rect 17276 4644 18420 4672
rect 17276 4632 17282 4644
rect 18414 4632 18420 4644
rect 18472 4632 18478 4684
rect 18966 4672 18972 4684
rect 18927 4644 18972 4672
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 21266 4672 21272 4684
rect 21227 4644 21272 4672
rect 21266 4632 21272 4644
rect 21324 4632 21330 4684
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 15654 4564 15660 4616
rect 15712 4604 15718 4616
rect 16114 4604 16120 4616
rect 15712 4576 16120 4604
rect 15712 4564 15718 4576
rect 16114 4564 16120 4576
rect 16172 4564 16178 4616
rect 19150 4604 19156 4616
rect 19111 4576 19156 4604
rect 19150 4564 19156 4576
rect 19208 4604 19214 4616
rect 19613 4607 19671 4613
rect 19613 4604 19625 4607
rect 19208 4576 19625 4604
rect 19208 4564 19214 4576
rect 19613 4573 19625 4576
rect 19659 4573 19671 4607
rect 19613 4567 19671 4573
rect 20714 4564 20720 4616
rect 20772 4604 20778 4616
rect 21468 4613 21496 4712
rect 22925 4709 22937 4743
rect 22971 4740 22983 4743
rect 23106 4740 23112 4752
rect 22971 4712 23112 4740
rect 22971 4709 22983 4712
rect 22925 4703 22983 4709
rect 23106 4700 23112 4712
rect 23164 4700 23170 4752
rect 25038 4740 25044 4752
rect 24999 4712 25044 4740
rect 25038 4700 25044 4712
rect 25096 4700 25102 4752
rect 22830 4672 22836 4684
rect 22791 4644 22836 4672
rect 22830 4632 22836 4644
rect 22888 4632 22894 4684
rect 24489 4675 24547 4681
rect 24489 4641 24501 4675
rect 24535 4672 24547 4675
rect 24670 4672 24676 4684
rect 24535 4644 24676 4672
rect 24535 4641 24547 4644
rect 24489 4635 24547 4641
rect 24670 4632 24676 4644
rect 24728 4632 24734 4684
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 20772 4576 21373 4604
rect 20772 4564 20778 4576
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 21361 4567 21419 4573
rect 21453 4607 21511 4613
rect 21453 4573 21465 4607
rect 21499 4604 21511 4607
rect 23014 4604 23020 4616
rect 21499 4576 23020 4604
rect 21499 4573 21511 4576
rect 21453 4567 21511 4573
rect 23014 4564 23020 4576
rect 23072 4564 23078 4616
rect 23658 4564 23664 4616
rect 23716 4604 23722 4616
rect 24210 4604 24216 4616
rect 23716 4576 24216 4604
rect 23716 4564 23722 4576
rect 24210 4564 24216 4576
rect 24268 4564 24274 4616
rect 12023 4508 12756 4536
rect 12023 4505 12035 4508
rect 11977 4499 12035 4505
rect 18782 4496 18788 4548
rect 18840 4536 18846 4548
rect 23290 4536 23296 4548
rect 18840 4508 23296 4536
rect 18840 4496 18846 4508
rect 23290 4496 23296 4508
rect 23348 4496 23354 4548
rect 23382 4496 23388 4548
rect 23440 4536 23446 4548
rect 25777 4539 25835 4545
rect 25777 4536 25789 4539
rect 23440 4508 25789 4536
rect 23440 4496 23446 4508
rect 25777 4505 25789 4508
rect 25823 4505 25835 4539
rect 25777 4499 25835 4505
rect 5445 4471 5503 4477
rect 5445 4468 5457 4471
rect 4304 4440 5457 4468
rect 4304 4428 4310 4440
rect 5445 4437 5457 4440
rect 5491 4437 5503 4471
rect 5445 4431 5503 4437
rect 7929 4471 7987 4477
rect 7929 4437 7941 4471
rect 7975 4468 7987 4471
rect 8573 4471 8631 4477
rect 8573 4468 8585 4471
rect 7975 4440 8585 4468
rect 7975 4437 7987 4440
rect 7929 4431 7987 4437
rect 8573 4437 8585 4440
rect 8619 4468 8631 4471
rect 8846 4468 8852 4480
rect 8619 4440 8852 4468
rect 8619 4437 8631 4440
rect 8573 4431 8631 4437
rect 8846 4428 8852 4440
rect 8904 4428 8910 4480
rect 9401 4471 9459 4477
rect 9401 4437 9413 4471
rect 9447 4468 9459 4471
rect 9490 4468 9496 4480
rect 9447 4440 9496 4468
rect 9447 4437 9459 4440
rect 9401 4431 9459 4437
rect 9490 4428 9496 4440
rect 9548 4428 9554 4480
rect 10318 4468 10324 4480
rect 10279 4440 10324 4468
rect 10318 4428 10324 4440
rect 10376 4428 10382 4480
rect 12066 4468 12072 4480
rect 12027 4440 12072 4468
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 14734 4468 14740 4480
rect 14695 4440 14740 4468
rect 14734 4428 14740 4440
rect 14792 4428 14798 4480
rect 15565 4471 15623 4477
rect 15565 4437 15577 4471
rect 15611 4468 15623 4471
rect 16022 4468 16028 4480
rect 15611 4440 16028 4468
rect 15611 4437 15623 4440
rect 15565 4431 15623 4437
rect 16022 4428 16028 4440
rect 16080 4468 16086 4480
rect 16850 4468 16856 4480
rect 16080 4440 16856 4468
rect 16080 4428 16086 4440
rect 16850 4428 16856 4440
rect 16908 4468 16914 4480
rect 17497 4471 17555 4477
rect 17497 4468 17509 4471
rect 16908 4440 17509 4468
rect 16908 4428 16914 4440
rect 17497 4437 17509 4440
rect 17543 4437 17555 4471
rect 17497 4431 17555 4437
rect 18601 4471 18659 4477
rect 18601 4437 18613 4471
rect 18647 4468 18659 4471
rect 18690 4468 18696 4480
rect 18647 4440 18696 4468
rect 18647 4437 18659 4440
rect 18601 4431 18659 4437
rect 18690 4428 18696 4440
rect 18748 4428 18754 4480
rect 19978 4468 19984 4480
rect 19939 4440 19984 4468
rect 19978 4428 19984 4440
rect 20036 4428 20042 4480
rect 20901 4471 20959 4477
rect 20901 4437 20913 4471
rect 20947 4468 20959 4471
rect 21910 4468 21916 4480
rect 20947 4440 21916 4468
rect 20947 4437 20959 4440
rect 20901 4431 20959 4437
rect 21910 4428 21916 4440
rect 21968 4428 21974 4480
rect 22465 4471 22523 4477
rect 22465 4437 22477 4471
rect 22511 4468 22523 4471
rect 23566 4468 23572 4480
rect 22511 4440 23572 4468
rect 22511 4437 22523 4440
rect 22465 4431 22523 4437
rect 23566 4428 23572 4440
rect 23624 4428 23630 4480
rect 24210 4428 24216 4480
rect 24268 4468 24274 4480
rect 24673 4471 24731 4477
rect 24673 4468 24685 4471
rect 24268 4440 24685 4468
rect 24268 4428 24274 4440
rect 24673 4437 24685 4440
rect 24719 4437 24731 4471
rect 24673 4431 24731 4437
rect 24762 4428 24768 4480
rect 24820 4468 24826 4480
rect 25409 4471 25467 4477
rect 25409 4468 25421 4471
rect 24820 4440 25421 4468
rect 24820 4428 24826 4440
rect 25409 4437 25421 4440
rect 25455 4437 25467 4471
rect 26234 4468 26240 4480
rect 26195 4440 26240 4468
rect 25409 4431 25467 4437
rect 26234 4428 26240 4440
rect 26292 4428 26298 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 2958 4264 2964 4276
rect 2919 4236 2964 4264
rect 2958 4224 2964 4236
rect 3016 4224 3022 4276
rect 3418 4264 3424 4276
rect 3379 4236 3424 4264
rect 3418 4224 3424 4236
rect 3476 4224 3482 4276
rect 5350 4224 5356 4276
rect 5408 4264 5414 4276
rect 18966 4264 18972 4276
rect 5408 4236 9536 4264
rect 5408 4224 5414 4236
rect 1765 4199 1823 4205
rect 1765 4165 1777 4199
rect 1811 4196 1823 4199
rect 2314 4196 2320 4208
rect 1811 4168 2320 4196
rect 1811 4165 1823 4168
rect 1765 4159 1823 4165
rect 2314 4156 2320 4168
rect 2372 4196 2378 4208
rect 2372 4168 2452 4196
rect 2372 4156 2378 4168
rect 2424 4137 2452 4168
rect 5442 4156 5448 4208
rect 5500 4196 5506 4208
rect 6086 4196 6092 4208
rect 5500 4168 6092 4196
rect 5500 4156 5506 4168
rect 6086 4156 6092 4168
rect 6144 4156 6150 4208
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4097 2467 4131
rect 3970 4128 3976 4140
rect 3931 4100 3976 4128
rect 2409 4091 2467 4097
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 4982 4128 4988 4140
rect 4943 4100 4988 4128
rect 4982 4088 4988 4100
rect 5040 4128 5046 4140
rect 5813 4131 5871 4137
rect 5040 4100 5580 4128
rect 5040 4088 5046 4100
rect 2130 4020 2136 4072
rect 2188 4060 2194 4072
rect 2225 4063 2283 4069
rect 2225 4060 2237 4063
rect 2188 4032 2237 4060
rect 2188 4020 2194 4032
rect 2225 4029 2237 4032
rect 2271 4029 2283 4063
rect 2225 4023 2283 4029
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 2682 4060 2688 4072
rect 2363 4032 2688 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 5552 4069 5580 4100
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 6196 4128 6224 4236
rect 9508 4208 9536 4236
rect 14016 4236 18972 4264
rect 9490 4156 9496 4208
rect 9548 4196 9554 4208
rect 13538 4196 13544 4208
rect 9548 4168 9904 4196
rect 9548 4156 9554 4168
rect 9122 4128 9128 4140
rect 5859 4100 6224 4128
rect 9035 4100 9128 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 9122 4088 9128 4100
rect 9180 4128 9186 4140
rect 9876 4137 9904 4168
rect 12452 4168 13544 4196
rect 12452 4140 12480 4168
rect 13538 4156 13544 4168
rect 13596 4156 13602 4208
rect 9769 4131 9827 4137
rect 9769 4128 9781 4131
rect 9180 4100 9781 4128
rect 9180 4088 9186 4100
rect 9769 4097 9781 4100
rect 9815 4097 9827 4131
rect 9769 4091 9827 4097
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4097 9919 4131
rect 11514 4128 11520 4140
rect 11427 4100 11520 4128
rect 9861 4091 9919 4097
rect 11514 4088 11520 4100
rect 11572 4128 11578 4140
rect 12342 4128 12348 4140
rect 11572 4100 12348 4128
rect 11572 4088 11578 4100
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 12434 4088 12440 4140
rect 12492 4088 12498 4140
rect 13170 4128 13176 4140
rect 13131 4100 13176 4128
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4128 13415 4131
rect 13446 4128 13452 4140
rect 13403 4100 13452 4128
rect 13403 4097 13415 4100
rect 13357 4091 13415 4097
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 14016 4128 14044 4236
rect 18966 4224 18972 4236
rect 19024 4264 19030 4276
rect 19061 4267 19119 4273
rect 19061 4264 19073 4267
rect 19024 4236 19073 4264
rect 19024 4224 19030 4236
rect 19061 4233 19073 4236
rect 19107 4233 19119 4267
rect 19061 4227 19119 4233
rect 19613 4267 19671 4273
rect 19613 4233 19625 4267
rect 19659 4264 19671 4267
rect 20162 4264 20168 4276
rect 19659 4236 20168 4264
rect 19659 4233 19671 4236
rect 19613 4227 19671 4233
rect 20162 4224 20168 4236
rect 20220 4224 20226 4276
rect 22557 4267 22615 4273
rect 22557 4233 22569 4267
rect 22603 4264 22615 4267
rect 23106 4264 23112 4276
rect 22603 4236 23112 4264
rect 22603 4233 22615 4236
rect 22557 4227 22615 4233
rect 23106 4224 23112 4236
rect 23164 4224 23170 4276
rect 24670 4264 24676 4276
rect 24631 4236 24676 4264
rect 24670 4224 24676 4236
rect 24728 4224 24734 4276
rect 24857 4267 24915 4273
rect 24857 4233 24869 4267
rect 24903 4264 24915 4267
rect 25222 4264 25228 4276
rect 24903 4236 25228 4264
rect 24903 4233 24915 4236
rect 24857 4227 24915 4233
rect 25222 4224 25228 4236
rect 25280 4224 25286 4276
rect 14090 4156 14096 4208
rect 14148 4196 14154 4208
rect 14185 4199 14243 4205
rect 14185 4196 14197 4199
rect 14148 4168 14197 4196
rect 14148 4156 14154 4168
rect 14185 4165 14197 4168
rect 14231 4196 14243 4199
rect 15010 4196 15016 4208
rect 14231 4168 15016 4196
rect 14231 4165 14243 4168
rect 14185 4159 14243 4165
rect 15010 4156 15016 4168
rect 15068 4156 15074 4208
rect 15378 4156 15384 4208
rect 15436 4196 15442 4208
rect 15436 4168 16988 4196
rect 15436 4156 15442 4168
rect 14918 4128 14924 4140
rect 13648 4100 14044 4128
rect 14879 4100 14924 4128
rect 5537 4063 5595 4069
rect 5537 4029 5549 4063
rect 5583 4060 5595 4063
rect 6086 4060 6092 4072
rect 5583 4032 6092 4060
rect 5583 4029 5595 4032
rect 5537 4023 5595 4029
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 6178 4020 6184 4072
rect 6236 4060 6242 4072
rect 6362 4060 6368 4072
rect 6236 4032 6368 4060
rect 6236 4020 6242 4032
rect 6362 4020 6368 4032
rect 6420 4020 6426 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6564 4032 6837 4060
rect 1872 3964 2452 3992
rect 1872 3933 1900 3964
rect 1857 3927 1915 3933
rect 1857 3893 1869 3927
rect 1903 3893 1915 3927
rect 2424 3924 2452 3964
rect 2498 3952 2504 4004
rect 2556 3992 2562 4004
rect 3329 3995 3387 4001
rect 3329 3992 3341 3995
rect 2556 3964 3341 3992
rect 2556 3952 2562 3964
rect 3329 3961 3341 3964
rect 3375 3992 3387 3995
rect 3878 3992 3884 4004
rect 3375 3964 3884 3992
rect 3375 3961 3387 3964
rect 3329 3955 3387 3961
rect 3878 3952 3884 3964
rect 3936 3952 3942 4004
rect 4154 3952 4160 4004
rect 4212 3992 4218 4004
rect 5258 3992 5264 4004
rect 4212 3964 5264 3992
rect 4212 3952 4218 3964
rect 5258 3952 5264 3964
rect 5316 3992 5322 4004
rect 5629 3995 5687 4001
rect 5629 3992 5641 3995
rect 5316 3964 5641 3992
rect 5316 3952 5322 3964
rect 5629 3961 5641 3964
rect 5675 3961 5687 3995
rect 5629 3955 5687 3961
rect 6564 3936 6592 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 9306 4020 9312 4072
rect 9364 4060 9370 4072
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 9364 4032 9689 4060
rect 9364 4020 9370 4032
rect 9677 4029 9689 4032
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 11054 4020 11060 4072
rect 11112 4060 11118 4072
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 11112 4032 12173 4060
rect 11112 4020 11118 4032
rect 12161 4029 12173 4032
rect 12207 4060 12219 4063
rect 13081 4063 13139 4069
rect 13081 4060 13093 4063
rect 12207 4032 13093 4060
rect 12207 4029 12219 4032
rect 12161 4023 12219 4029
rect 13081 4029 13093 4032
rect 13127 4060 13139 4063
rect 13648 4060 13676 4100
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 15286 4128 15292 4140
rect 15247 4100 15292 4128
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 16117 4131 16175 4137
rect 16117 4097 16129 4131
rect 16163 4128 16175 4131
rect 16390 4128 16396 4140
rect 16163 4100 16396 4128
rect 16163 4097 16175 4100
rect 16117 4091 16175 4097
rect 16390 4088 16396 4100
rect 16448 4128 16454 4140
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16448 4100 16681 4128
rect 16448 4088 16454 4100
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16850 4128 16856 4140
rect 16811 4100 16856 4128
rect 16669 4091 16727 4097
rect 16850 4088 16856 4100
rect 16908 4088 16914 4140
rect 16960 4128 16988 4168
rect 18414 4156 18420 4208
rect 18472 4196 18478 4208
rect 18472 4168 18644 4196
rect 18472 4156 18478 4168
rect 18616 4137 18644 4168
rect 18690 4156 18696 4208
rect 18748 4196 18754 4208
rect 18748 4168 19288 4196
rect 18748 4156 18754 4168
rect 17773 4131 17831 4137
rect 17773 4128 17785 4131
rect 16960 4100 17785 4128
rect 17773 4097 17785 4100
rect 17819 4128 17831 4131
rect 18509 4131 18567 4137
rect 18509 4128 18521 4131
rect 17819 4100 18521 4128
rect 17819 4097 17831 4100
rect 17773 4091 17831 4097
rect 18509 4097 18521 4100
rect 18555 4097 18567 4131
rect 18509 4091 18567 4097
rect 18601 4131 18659 4137
rect 18601 4097 18613 4131
rect 18647 4097 18659 4131
rect 19260 4128 19288 4168
rect 19978 4156 19984 4208
rect 20036 4196 20042 4208
rect 26234 4196 26240 4208
rect 20036 4168 20208 4196
rect 20036 4156 20042 4168
rect 20180 4137 20208 4168
rect 20640 4168 26240 4196
rect 20165 4131 20223 4137
rect 19260 4100 20116 4128
rect 18601 4091 18659 4097
rect 13127 4032 13676 4060
rect 13817 4063 13875 4069
rect 13127 4029 13139 4032
rect 13081 4023 13139 4029
rect 13817 4029 13829 4063
rect 13863 4060 13875 4063
rect 14366 4060 14372 4072
rect 13863 4032 14372 4060
rect 13863 4029 13875 4032
rect 13817 4023 13875 4029
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 14642 4060 14648 4072
rect 14603 4032 14648 4060
rect 14642 4020 14648 4032
rect 14700 4020 14706 4072
rect 15304 4060 15332 4088
rect 16577 4063 16635 4069
rect 16577 4060 16589 4063
rect 15304 4032 16589 4060
rect 16577 4029 16589 4032
rect 16623 4029 16635 4063
rect 16577 4023 16635 4029
rect 17218 4020 17224 4072
rect 17276 4060 17282 4072
rect 17405 4063 17463 4069
rect 17405 4060 17417 4063
rect 17276 4032 17417 4060
rect 17276 4020 17282 4032
rect 17405 4029 17417 4032
rect 17451 4029 17463 4063
rect 17405 4023 17463 4029
rect 18230 4020 18236 4072
rect 18288 4060 18294 4072
rect 18417 4063 18475 4069
rect 18417 4060 18429 4063
rect 18288 4032 18429 4060
rect 18288 4020 18294 4032
rect 18417 4029 18429 4032
rect 18463 4060 18475 4063
rect 18874 4060 18880 4072
rect 18463 4032 18880 4060
rect 18463 4029 18475 4032
rect 18417 4023 18475 4029
rect 18874 4020 18880 4032
rect 18932 4020 18938 4072
rect 20088 4069 20116 4100
rect 20165 4097 20177 4131
rect 20211 4097 20223 4131
rect 20165 4091 20223 4097
rect 20073 4063 20131 4069
rect 20073 4029 20085 4063
rect 20119 4060 20131 4063
rect 20254 4060 20260 4072
rect 20119 4032 20260 4060
rect 20119 4029 20131 4032
rect 20073 4023 20131 4029
rect 20254 4020 20260 4032
rect 20312 4020 20318 4072
rect 20346 4020 20352 4072
rect 20404 4060 20410 4072
rect 20640 4060 20668 4168
rect 26234 4156 26240 4168
rect 26292 4156 26298 4208
rect 21726 4128 21732 4140
rect 21687 4100 21732 4128
rect 21726 4088 21732 4100
rect 21784 4088 21790 4140
rect 23474 4088 23480 4140
rect 23532 4128 23538 4140
rect 24213 4131 24271 4137
rect 24213 4128 24225 4131
rect 23532 4100 24225 4128
rect 23532 4088 23538 4100
rect 24213 4097 24225 4100
rect 24259 4097 24271 4131
rect 24213 4091 24271 4097
rect 24946 4088 24952 4140
rect 25004 4128 25010 4140
rect 25004 4100 25268 4128
rect 25004 4088 25010 4100
rect 20404 4032 20668 4060
rect 20404 4020 20410 4032
rect 20990 4020 20996 4072
rect 21048 4060 21054 4072
rect 21545 4063 21603 4069
rect 21545 4060 21557 4063
rect 21048 4032 21557 4060
rect 21048 4020 21054 4032
rect 21545 4029 21557 4032
rect 21591 4029 21603 4063
rect 21545 4023 21603 4029
rect 22554 4020 22560 4072
rect 22612 4060 22618 4072
rect 23750 4060 23756 4072
rect 22612 4032 23756 4060
rect 22612 4020 22618 4032
rect 23750 4020 23756 4032
rect 23808 4020 23814 4072
rect 24857 4063 24915 4069
rect 24857 4060 24869 4063
rect 23860 4032 24869 4060
rect 7092 3995 7150 4001
rect 7092 3961 7104 3995
rect 7138 3992 7150 3995
rect 7466 3992 7472 4004
rect 7138 3964 7472 3992
rect 7138 3961 7150 3964
rect 7092 3955 7150 3961
rect 7466 3952 7472 3964
rect 7524 3992 7530 4004
rect 14734 3992 14740 4004
rect 7524 3964 8892 3992
rect 7524 3952 7530 3964
rect 8864 3936 8892 3964
rect 12728 3964 14740 3992
rect 2682 3924 2688 3936
rect 2424 3896 2688 3924
rect 1857 3887 1915 3893
rect 2682 3884 2688 3896
rect 2740 3884 2746 3936
rect 3786 3924 3792 3936
rect 3747 3896 3792 3924
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 4525 3927 4583 3933
rect 4525 3893 4537 3927
rect 4571 3924 4583 3927
rect 4614 3924 4620 3936
rect 4571 3896 4620 3924
rect 4571 3893 4583 3896
rect 4525 3887 4583 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 5074 3884 5080 3936
rect 5132 3924 5138 3936
rect 5169 3927 5227 3933
rect 5169 3924 5181 3927
rect 5132 3896 5181 3924
rect 5132 3884 5138 3896
rect 5169 3893 5181 3896
rect 5215 3893 5227 3927
rect 6178 3924 6184 3936
rect 6139 3896 6184 3924
rect 5169 3887 5227 3893
rect 6178 3884 6184 3896
rect 6236 3924 6242 3936
rect 6546 3924 6552 3936
rect 6236 3896 6552 3924
rect 6236 3884 6242 3896
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 6972 3896 8217 3924
rect 6972 3884 6978 3896
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 8846 3924 8852 3936
rect 8807 3896 8852 3924
rect 8205 3887 8263 3893
rect 8846 3884 8852 3896
rect 8904 3884 8910 3936
rect 9309 3927 9367 3933
rect 9309 3893 9321 3927
rect 9355 3924 9367 3927
rect 9398 3924 9404 3936
rect 9355 3896 9404 3924
rect 9355 3893 9367 3896
rect 9309 3887 9367 3893
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 10505 3927 10563 3933
rect 10505 3893 10517 3927
rect 10551 3924 10563 3927
rect 10778 3924 10784 3936
rect 10551 3896 10784 3924
rect 10551 3893 10563 3896
rect 10505 3887 10563 3893
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 10873 3927 10931 3933
rect 10873 3893 10885 3927
rect 10919 3924 10931 3927
rect 10962 3924 10968 3936
rect 10919 3896 10968 3924
rect 10919 3893 10931 3896
rect 10873 3887 10931 3893
rect 10962 3884 10968 3896
rect 11020 3884 11026 3936
rect 11885 3927 11943 3933
rect 11885 3893 11897 3927
rect 11931 3924 11943 3927
rect 11974 3924 11980 3936
rect 11931 3896 11980 3924
rect 11931 3893 11943 3896
rect 11885 3887 11943 3893
rect 11974 3884 11980 3896
rect 12032 3924 12038 3936
rect 12526 3924 12532 3936
rect 12032 3896 12532 3924
rect 12032 3884 12038 3896
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 12728 3933 12756 3964
rect 14734 3952 14740 3964
rect 14792 3952 14798 4004
rect 20162 3952 20168 4004
rect 20220 3992 20226 4004
rect 21085 3995 21143 4001
rect 21085 3992 21097 3995
rect 20220 3964 21097 3992
rect 20220 3952 20226 3964
rect 21085 3961 21097 3964
rect 21131 3992 21143 3995
rect 21637 3995 21695 4001
rect 21637 3992 21649 3995
rect 21131 3964 21649 3992
rect 21131 3961 21143 3964
rect 21085 3955 21143 3961
rect 21637 3961 21649 3964
rect 21683 3992 21695 3995
rect 22094 3992 22100 4004
rect 21683 3964 22100 3992
rect 21683 3961 21695 3964
rect 21637 3955 21695 3961
rect 22094 3952 22100 3964
rect 22152 3952 22158 4004
rect 22186 3952 22192 4004
rect 22244 3992 22250 4004
rect 23860 3992 23888 4032
rect 24857 4029 24869 4032
rect 24903 4029 24915 4063
rect 25038 4060 25044 4072
rect 24999 4032 25044 4060
rect 24857 4023 24915 4029
rect 25038 4020 25044 4032
rect 25096 4020 25102 4072
rect 25240 4069 25268 4100
rect 25225 4063 25283 4069
rect 25225 4029 25237 4063
rect 25271 4060 25283 4063
rect 25777 4063 25835 4069
rect 25777 4060 25789 4063
rect 25271 4032 25789 4060
rect 25271 4029 25283 4032
rect 25225 4023 25283 4029
rect 25777 4029 25789 4032
rect 25823 4029 25835 4063
rect 25777 4023 25835 4029
rect 22244 3964 23888 3992
rect 22244 3952 22250 3964
rect 23934 3952 23940 4004
rect 23992 3992 23998 4004
rect 24121 3995 24179 4001
rect 24121 3992 24133 3995
rect 23992 3964 24133 3992
rect 23992 3952 23998 3964
rect 24121 3961 24133 3964
rect 24167 3992 24179 3995
rect 26237 3995 26295 4001
rect 26237 3992 26249 3995
rect 24167 3964 26249 3992
rect 24167 3961 24179 3964
rect 24121 3955 24179 3961
rect 26237 3961 26249 3964
rect 26283 3961 26295 3995
rect 26237 3955 26295 3961
rect 12713 3927 12771 3933
rect 12713 3893 12725 3927
rect 12759 3893 12771 3927
rect 14274 3924 14280 3936
rect 14235 3896 14280 3924
rect 12713 3887 12771 3893
rect 14274 3884 14280 3896
rect 14332 3884 14338 3936
rect 15286 3884 15292 3936
rect 15344 3924 15350 3936
rect 15654 3924 15660 3936
rect 15344 3896 15660 3924
rect 15344 3884 15350 3896
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 16206 3924 16212 3936
rect 16167 3896 16212 3924
rect 16206 3884 16212 3896
rect 16264 3884 16270 3936
rect 18046 3924 18052 3936
rect 18007 3896 18052 3924
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 19426 3924 19432 3936
rect 19387 3896 19432 3924
rect 19426 3884 19432 3896
rect 19484 3924 19490 3936
rect 19981 3927 20039 3933
rect 19981 3924 19993 3927
rect 19484 3896 19993 3924
rect 19484 3884 19490 3896
rect 19981 3893 19993 3896
rect 20027 3893 20039 3927
rect 19981 3887 20039 3893
rect 20717 3927 20775 3933
rect 20717 3893 20729 3927
rect 20763 3924 20775 3927
rect 20990 3924 20996 3936
rect 20763 3896 20996 3924
rect 20763 3893 20775 3896
rect 20717 3887 20775 3893
rect 20990 3884 20996 3896
rect 21048 3884 21054 3936
rect 21174 3924 21180 3936
rect 21135 3896 21180 3924
rect 21174 3884 21180 3896
rect 21232 3884 21238 3936
rect 22830 3924 22836 3936
rect 22791 3896 22836 3924
rect 22830 3884 22836 3896
rect 22888 3884 22894 3936
rect 23382 3924 23388 3936
rect 23343 3896 23388 3924
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 23661 3927 23719 3933
rect 23661 3893 23673 3927
rect 23707 3924 23719 3927
rect 23750 3924 23756 3936
rect 23707 3896 23756 3924
rect 23707 3893 23719 3896
rect 23661 3887 23719 3893
rect 23750 3884 23756 3896
rect 23808 3884 23814 3936
rect 24026 3924 24032 3936
rect 23987 3896 24032 3924
rect 24026 3884 24032 3896
rect 24084 3884 24090 3936
rect 25406 3924 25412 3936
rect 25367 3896 25412 3924
rect 25406 3884 25412 3896
rect 25464 3884 25470 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 2409 3723 2467 3729
rect 2409 3689 2421 3723
rect 2455 3720 2467 3723
rect 2682 3720 2688 3732
rect 2455 3692 2688 3720
rect 2455 3689 2467 3692
rect 2409 3683 2467 3689
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 3513 3723 3571 3729
rect 3513 3689 3525 3723
rect 3559 3720 3571 3723
rect 3786 3720 3792 3732
rect 3559 3692 3792 3720
rect 3559 3689 3571 3692
rect 3513 3683 3571 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 4062 3720 4068 3732
rect 4023 3692 4068 3720
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 4522 3720 4528 3732
rect 4483 3692 4528 3720
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 5258 3720 5264 3732
rect 5219 3692 5264 3720
rect 5258 3680 5264 3692
rect 5316 3680 5322 3732
rect 9306 3720 9312 3732
rect 9267 3692 9312 3720
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 10134 3720 10140 3732
rect 9732 3692 9777 3720
rect 10095 3692 10140 3720
rect 9732 3680 9738 3692
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 10781 3723 10839 3729
rect 10781 3689 10793 3723
rect 10827 3720 10839 3723
rect 10870 3720 10876 3732
rect 10827 3692 10876 3720
rect 10827 3689 10839 3692
rect 10781 3683 10839 3689
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 13078 3720 13084 3732
rect 11204 3692 13084 3720
rect 11204 3680 11210 3692
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 13722 3720 13728 3732
rect 13683 3692 13728 3720
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 14182 3720 14188 3732
rect 14143 3692 14188 3720
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 14642 3680 14648 3732
rect 14700 3720 14706 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 14700 3692 15025 3720
rect 14700 3680 14706 3692
rect 15013 3689 15025 3692
rect 15059 3689 15071 3723
rect 15013 3683 15071 3689
rect 15470 3680 15476 3732
rect 15528 3720 15534 3732
rect 16298 3720 16304 3732
rect 15528 3692 16304 3720
rect 15528 3680 15534 3692
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 16482 3680 16488 3732
rect 16540 3720 16546 3732
rect 17865 3723 17923 3729
rect 17865 3720 17877 3723
rect 16540 3692 17877 3720
rect 16540 3680 16546 3692
rect 17865 3689 17877 3692
rect 17911 3689 17923 3723
rect 18598 3720 18604 3732
rect 18559 3692 18604 3720
rect 17865 3683 17923 3689
rect 18598 3680 18604 3692
rect 18656 3680 18662 3732
rect 18969 3723 19027 3729
rect 18969 3689 18981 3723
rect 19015 3720 19027 3723
rect 19058 3720 19064 3732
rect 19015 3692 19064 3720
rect 19015 3689 19027 3692
rect 18969 3683 19027 3689
rect 19058 3680 19064 3692
rect 19116 3680 19122 3732
rect 19429 3723 19487 3729
rect 19429 3689 19441 3723
rect 19475 3720 19487 3723
rect 20346 3720 20352 3732
rect 19475 3692 20352 3720
rect 19475 3689 19487 3692
rect 19429 3683 19487 3689
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 20901 3723 20959 3729
rect 20901 3689 20913 3723
rect 20947 3689 20959 3723
rect 21358 3720 21364 3732
rect 21319 3692 21364 3720
rect 20901 3683 20959 3689
rect 2314 3652 2320 3664
rect 2227 3624 2320 3652
rect 2314 3612 2320 3624
rect 2372 3652 2378 3664
rect 2372 3624 3004 3652
rect 2372 3612 2378 3624
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3584 2007 3587
rect 2038 3584 2044 3596
rect 1995 3556 2044 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 1412 3516 1440 3547
rect 2038 3544 2044 3556
rect 2096 3584 2102 3596
rect 2777 3587 2835 3593
rect 2777 3584 2789 3587
rect 2096 3556 2789 3584
rect 2096 3544 2102 3556
rect 2777 3553 2789 3556
rect 2823 3553 2835 3587
rect 2777 3547 2835 3553
rect 2222 3516 2228 3528
rect 1412 3488 2228 3516
rect 2222 3476 2228 3488
rect 2280 3476 2286 3528
rect 2976 3525 3004 3624
rect 4614 3612 4620 3664
rect 4672 3652 4678 3664
rect 5629 3655 5687 3661
rect 5629 3652 5641 3655
rect 4672 3624 5641 3652
rect 4672 3612 4678 3624
rect 5629 3621 5641 3624
rect 5675 3652 5687 3655
rect 6178 3652 6184 3664
rect 5675 3624 6184 3652
rect 5675 3621 5687 3624
rect 5629 3615 5687 3621
rect 4430 3584 4436 3596
rect 4391 3556 4436 3584
rect 4430 3544 4436 3556
rect 4488 3544 4494 3596
rect 5828 3593 5856 3624
rect 6178 3612 6184 3624
rect 6236 3612 6242 3664
rect 8846 3612 8852 3664
rect 8904 3652 8910 3664
rect 11517 3655 11575 3661
rect 11517 3652 11529 3655
rect 8904 3624 11529 3652
rect 8904 3612 8910 3624
rect 5813 3587 5871 3593
rect 4724 3556 5304 3584
rect 2869 3519 2927 3525
rect 2869 3485 2881 3519
rect 2915 3485 2927 3519
rect 2869 3479 2927 3485
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3485 3019 3519
rect 2961 3479 3019 3485
rect 3881 3519 3939 3525
rect 3881 3485 3893 3519
rect 3927 3516 3939 3519
rect 3970 3516 3976 3528
rect 3927 3488 3976 3516
rect 3927 3485 3939 3488
rect 3881 3479 3939 3485
rect 2884 3448 2912 3479
rect 3970 3476 3976 3488
rect 4028 3516 4034 3528
rect 4724 3525 4752 3556
rect 4709 3519 4767 3525
rect 4709 3516 4721 3519
rect 4028 3488 4721 3516
rect 4028 3476 4034 3488
rect 4709 3485 4721 3488
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 5166 3476 5172 3528
rect 5224 3476 5230 3528
rect 5184 3448 5212 3476
rect 2884 3420 5212 3448
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3380 1639 3383
rect 4798 3380 4804 3392
rect 1627 3352 4804 3380
rect 1627 3349 1639 3352
rect 1581 3343 1639 3349
rect 4798 3340 4804 3352
rect 4856 3340 4862 3392
rect 5276 3380 5304 3556
rect 5813 3553 5825 3587
rect 5859 3553 5871 3587
rect 5813 3547 5871 3553
rect 5902 3544 5908 3596
rect 5960 3584 5966 3596
rect 6069 3587 6127 3593
rect 6069 3584 6081 3587
rect 5960 3556 6081 3584
rect 5960 3544 5966 3556
rect 6069 3553 6081 3556
rect 6115 3553 6127 3587
rect 8570 3584 8576 3596
rect 8531 3556 8576 3584
rect 6069 3547 6127 3553
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 9858 3544 9864 3596
rect 9916 3584 9922 3596
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 9916 3556 10057 3584
rect 9916 3544 9922 3556
rect 10045 3553 10057 3556
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 10336 3525 10364 3624
rect 11517 3621 11529 3624
rect 11563 3652 11575 3655
rect 11606 3652 11612 3664
rect 11563 3624 11612 3652
rect 11563 3621 11575 3624
rect 11517 3615 11575 3621
rect 11606 3612 11612 3624
rect 11664 3612 11670 3664
rect 14093 3655 14151 3661
rect 14093 3621 14105 3655
rect 14139 3652 14151 3655
rect 16500 3652 16528 3680
rect 14139 3624 16528 3652
rect 14139 3621 14151 3624
rect 14093 3615 14151 3621
rect 16758 3612 16764 3664
rect 16816 3652 16822 3664
rect 17221 3655 17279 3661
rect 17221 3652 17233 3655
rect 16816 3624 17233 3652
rect 16816 3612 16822 3624
rect 17221 3621 17233 3624
rect 17267 3652 17279 3655
rect 17586 3652 17592 3664
rect 17267 3624 17592 3652
rect 17267 3621 17279 3624
rect 17221 3615 17279 3621
rect 17586 3612 17592 3624
rect 17644 3612 17650 3664
rect 17770 3652 17776 3664
rect 17731 3624 17776 3652
rect 17770 3612 17776 3624
rect 17828 3612 17834 3664
rect 19337 3655 19395 3661
rect 19337 3621 19349 3655
rect 19383 3652 19395 3655
rect 19518 3652 19524 3664
rect 19383 3624 19524 3652
rect 19383 3621 19395 3624
rect 19337 3615 19395 3621
rect 11149 3587 11207 3593
rect 11149 3553 11161 3587
rect 11195 3584 11207 3587
rect 11238 3584 11244 3596
rect 11195 3556 11244 3584
rect 11195 3553 11207 3556
rect 11149 3547 11207 3553
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 11968 3587 12026 3593
rect 11968 3553 11980 3587
rect 12014 3584 12026 3587
rect 12250 3584 12256 3596
rect 12014 3556 12256 3584
rect 12014 3553 12026 3556
rect 11968 3547 12026 3553
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 16209 3587 16267 3593
rect 16209 3553 16221 3587
rect 16255 3584 16267 3587
rect 17034 3584 17040 3596
rect 16255 3556 17040 3584
rect 16255 3553 16267 3556
rect 16209 3547 16267 3553
rect 17034 3544 17040 3556
rect 17092 3544 17098 3596
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 11606 3476 11612 3528
rect 11664 3516 11670 3528
rect 11701 3519 11759 3525
rect 11701 3516 11713 3519
rect 11664 3488 11713 3516
rect 11664 3476 11670 3488
rect 11701 3485 11713 3488
rect 11747 3485 11759 3519
rect 11701 3479 11759 3485
rect 14737 3519 14795 3525
rect 14737 3485 14749 3519
rect 14783 3516 14795 3519
rect 14918 3516 14924 3528
rect 14783 3488 14924 3516
rect 14783 3485 14795 3488
rect 14737 3479 14795 3485
rect 14918 3476 14924 3488
rect 14976 3516 14982 3528
rect 15378 3516 15384 3528
rect 14976 3488 15384 3516
rect 14976 3476 14982 3488
rect 15378 3476 15384 3488
rect 15436 3516 15442 3528
rect 16485 3519 16543 3525
rect 16485 3516 16497 3519
rect 15436 3488 16497 3516
rect 15436 3476 15442 3488
rect 16485 3485 16497 3488
rect 16531 3516 16543 3519
rect 16850 3516 16856 3528
rect 16531 3488 16856 3516
rect 16531 3485 16543 3488
rect 16485 3479 16543 3485
rect 16850 3476 16856 3488
rect 16908 3476 16914 3528
rect 16945 3519 17003 3525
rect 16945 3485 16957 3519
rect 16991 3516 17003 3519
rect 17218 3516 17224 3528
rect 16991 3488 17224 3516
rect 16991 3485 17003 3488
rect 16945 3479 17003 3485
rect 17218 3476 17224 3488
rect 17276 3476 17282 3528
rect 17954 3516 17960 3528
rect 17915 3488 17960 3516
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 7193 3451 7251 3457
rect 7193 3417 7205 3451
rect 7239 3448 7251 3451
rect 7834 3448 7840 3460
rect 7239 3420 7840 3448
rect 7239 3417 7251 3420
rect 7193 3411 7251 3417
rect 7208 3380 7236 3411
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 14458 3408 14464 3460
rect 14516 3448 14522 3460
rect 19352 3448 19380 3615
rect 19518 3612 19524 3624
rect 19576 3612 19582 3664
rect 20916 3652 20944 3683
rect 21358 3680 21364 3692
rect 21416 3680 21422 3732
rect 23566 3680 23572 3732
rect 23624 3720 23630 3732
rect 24397 3723 24455 3729
rect 24397 3720 24409 3723
rect 23624 3692 24409 3720
rect 23624 3680 23630 3692
rect 24397 3689 24409 3692
rect 24443 3720 24455 3723
rect 24762 3720 24768 3732
rect 24443 3692 24768 3720
rect 24443 3689 24455 3692
rect 24397 3683 24455 3689
rect 24762 3680 24768 3692
rect 24820 3680 24826 3732
rect 21450 3652 21456 3664
rect 20916 3624 21456 3652
rect 21450 3612 21456 3624
rect 21508 3612 21514 3664
rect 23474 3652 23480 3664
rect 23435 3624 23480 3652
rect 23474 3612 23480 3624
rect 23532 3612 23538 3664
rect 25409 3655 25467 3661
rect 25409 3652 25421 3655
rect 23952 3624 25421 3652
rect 21266 3584 21272 3596
rect 21227 3556 21272 3584
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 22094 3544 22100 3596
rect 22152 3584 22158 3596
rect 22833 3587 22891 3593
rect 22833 3584 22845 3587
rect 22152 3556 22845 3584
rect 22152 3544 22158 3556
rect 22833 3553 22845 3556
rect 22879 3584 22891 3587
rect 23952 3584 23980 3624
rect 25409 3621 25421 3624
rect 25455 3621 25467 3655
rect 25409 3615 25467 3621
rect 22879 3556 23980 3584
rect 24489 3587 24547 3593
rect 22879 3553 22891 3556
rect 22833 3547 22891 3553
rect 24489 3553 24501 3587
rect 24535 3584 24547 3587
rect 26237 3587 26295 3593
rect 26237 3584 26249 3587
rect 24535 3556 26249 3584
rect 24535 3553 24547 3556
rect 24489 3547 24547 3553
rect 26237 3553 26249 3556
rect 26283 3553 26295 3587
rect 26237 3547 26295 3553
rect 19613 3519 19671 3525
rect 19613 3485 19625 3519
rect 19659 3516 19671 3519
rect 19978 3516 19984 3528
rect 19659 3488 19984 3516
rect 19659 3485 19671 3488
rect 19613 3479 19671 3485
rect 19978 3476 19984 3488
rect 20036 3476 20042 3528
rect 21453 3519 21511 3525
rect 21453 3516 21465 3519
rect 20640 3488 21465 3516
rect 14516 3420 19380 3448
rect 14516 3408 14522 3420
rect 5276 3352 7236 3380
rect 7282 3340 7288 3392
rect 7340 3380 7346 3392
rect 7745 3383 7803 3389
rect 7745 3380 7757 3383
rect 7340 3352 7757 3380
rect 7340 3340 7346 3352
rect 7745 3349 7757 3352
rect 7791 3349 7803 3383
rect 7745 3343 7803 3349
rect 8481 3383 8539 3389
rect 8481 3349 8493 3383
rect 8527 3380 8539 3383
rect 8662 3380 8668 3392
rect 8527 3352 8668 3380
rect 8527 3349 8539 3352
rect 8481 3343 8539 3349
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 8754 3340 8760 3392
rect 8812 3380 8818 3392
rect 15562 3380 15568 3392
rect 8812 3352 8857 3380
rect 15523 3352 15568 3380
rect 8812 3340 8818 3352
rect 15562 3340 15568 3352
rect 15620 3340 15626 3392
rect 15838 3380 15844 3392
rect 15799 3352 15844 3380
rect 15838 3340 15844 3352
rect 15896 3340 15902 3392
rect 17402 3380 17408 3392
rect 17363 3352 17408 3380
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 19978 3380 19984 3392
rect 19939 3352 19984 3380
rect 19978 3340 19984 3352
rect 20036 3380 20042 3392
rect 20640 3389 20668 3488
rect 21453 3485 21465 3488
rect 21499 3516 21511 3519
rect 21726 3516 21732 3528
rect 21499 3488 21732 3516
rect 21499 3485 21511 3488
rect 21453 3479 21511 3485
rect 21726 3476 21732 3488
rect 21784 3516 21790 3528
rect 21913 3519 21971 3525
rect 21913 3516 21925 3519
rect 21784 3488 21925 3516
rect 21784 3476 21790 3488
rect 21913 3485 21925 3488
rect 21959 3485 21971 3519
rect 21913 3479 21971 3485
rect 22002 3476 22008 3528
rect 22060 3516 22066 3528
rect 22922 3516 22928 3528
rect 22060 3488 22928 3516
rect 22060 3476 22066 3488
rect 22922 3476 22928 3488
rect 22980 3476 22986 3528
rect 23109 3519 23167 3525
rect 23109 3485 23121 3519
rect 23155 3485 23167 3519
rect 23109 3479 23167 3485
rect 22373 3451 22431 3457
rect 22373 3417 22385 3451
rect 22419 3448 22431 3451
rect 23014 3448 23020 3460
rect 22419 3420 23020 3448
rect 22419 3417 22431 3420
rect 22373 3411 22431 3417
rect 23014 3408 23020 3420
rect 23072 3448 23078 3460
rect 23124 3448 23152 3479
rect 23658 3476 23664 3528
rect 23716 3516 23722 3528
rect 24504 3516 24532 3547
rect 24670 3516 24676 3528
rect 23716 3488 24532 3516
rect 24631 3488 24676 3516
rect 23716 3476 23722 3488
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 24026 3448 24032 3460
rect 23072 3420 23152 3448
rect 23939 3420 24032 3448
rect 23072 3408 23078 3420
rect 24026 3408 24032 3420
rect 24084 3448 24090 3460
rect 25041 3451 25099 3457
rect 25041 3448 25053 3451
rect 24084 3420 25053 3448
rect 24084 3408 24090 3420
rect 25041 3417 25053 3420
rect 25087 3417 25099 3451
rect 25041 3411 25099 3417
rect 20625 3383 20683 3389
rect 20625 3380 20637 3383
rect 20036 3352 20637 3380
rect 20036 3340 20042 3352
rect 20625 3349 20637 3352
rect 20671 3349 20683 3383
rect 20625 3343 20683 3349
rect 22465 3383 22523 3389
rect 22465 3349 22477 3383
rect 22511 3380 22523 3383
rect 23474 3380 23480 3392
rect 22511 3352 23480 3380
rect 22511 3349 22523 3352
rect 22465 3343 22523 3349
rect 23474 3340 23480 3352
rect 23532 3340 23538 3392
rect 23842 3380 23848 3392
rect 23803 3352 23848 3380
rect 23842 3340 23848 3352
rect 23900 3340 23906 3392
rect 24762 3340 24768 3392
rect 24820 3380 24826 3392
rect 25777 3383 25835 3389
rect 25777 3380 25789 3383
rect 24820 3352 25789 3380
rect 24820 3340 24826 3352
rect 25777 3349 25789 3352
rect 25823 3349 25835 3383
rect 25777 3343 25835 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 2038 3176 2044 3188
rect 1999 3148 2044 3176
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 3605 3179 3663 3185
rect 3605 3176 3617 3179
rect 3068 3148 3617 3176
rect 1762 3068 1768 3120
rect 1820 3108 1826 3120
rect 2682 3108 2688 3120
rect 1820 3080 2688 3108
rect 1820 3068 1826 3080
rect 2682 3068 2688 3080
rect 2740 3068 2746 3120
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3040 2007 3043
rect 2593 3043 2651 3049
rect 2593 3040 2605 3043
rect 1995 3012 2605 3040
rect 1995 3009 2007 3012
rect 1949 3003 2007 3009
rect 2593 3009 2605 3012
rect 2639 3040 2651 3043
rect 2958 3040 2964 3052
rect 2639 3012 2964 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 2498 2972 2504 2984
rect 2459 2944 2504 2972
rect 2498 2932 2504 2944
rect 2556 2932 2562 2984
rect 3068 2972 3096 3148
rect 3605 3145 3617 3148
rect 3651 3176 3663 3179
rect 3694 3176 3700 3188
rect 3651 3148 3700 3176
rect 3651 3145 3663 3148
rect 3605 3139 3663 3145
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 4982 3176 4988 3188
rect 4488 3148 4988 3176
rect 4488 3136 4494 3148
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 5166 3176 5172 3188
rect 5127 3148 5172 3176
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 6178 3136 6184 3188
rect 6236 3176 6242 3188
rect 7190 3176 7196 3188
rect 6236 3148 7196 3176
rect 6236 3136 6242 3148
rect 7190 3136 7196 3148
rect 7248 3136 7254 3188
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 10321 3179 10379 3185
rect 10321 3176 10333 3179
rect 9916 3148 10333 3176
rect 9916 3136 9922 3148
rect 10321 3145 10333 3148
rect 10367 3145 10379 3179
rect 10321 3139 10379 3145
rect 10870 3136 10876 3188
rect 10928 3176 10934 3188
rect 11146 3176 11152 3188
rect 10928 3148 11152 3176
rect 10928 3136 10934 3148
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 12250 3176 12256 3188
rect 12211 3148 12256 3176
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 14369 3179 14427 3185
rect 14369 3145 14381 3179
rect 14415 3176 14427 3179
rect 15470 3176 15476 3188
rect 14415 3148 15476 3176
rect 14415 3145 14427 3148
rect 14369 3139 14427 3145
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 15562 3136 15568 3188
rect 15620 3176 15626 3188
rect 16209 3179 16267 3185
rect 16209 3176 16221 3179
rect 15620 3148 16221 3176
rect 15620 3136 15626 3148
rect 3510 3068 3516 3120
rect 3568 3108 3574 3120
rect 4522 3108 4528 3120
rect 3568 3080 4528 3108
rect 3568 3068 3574 3080
rect 4522 3068 4528 3080
rect 4580 3108 4586 3120
rect 4617 3111 4675 3117
rect 4617 3108 4629 3111
rect 4580 3080 4629 3108
rect 4580 3068 4586 3080
rect 4617 3077 4629 3080
rect 4663 3077 4675 3111
rect 6822 3108 6828 3120
rect 6783 3080 6828 3108
rect 4617 3071 4675 3077
rect 6822 3068 6828 3080
rect 6880 3068 6886 3120
rect 10134 3068 10140 3120
rect 10192 3108 10198 3120
rect 10689 3111 10747 3117
rect 10689 3108 10701 3111
rect 10192 3080 10701 3108
rect 10192 3068 10198 3080
rect 10689 3077 10701 3080
rect 10735 3077 10747 3111
rect 12158 3108 12164 3120
rect 10689 3071 10747 3077
rect 11164 3080 12164 3108
rect 11164 3052 11192 3080
rect 12158 3068 12164 3080
rect 12216 3068 12222 3120
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3040 3203 3043
rect 3970 3040 3976 3052
rect 3191 3012 3976 3040
rect 3191 3009 3203 3012
rect 3145 3003 3203 3009
rect 3970 3000 3976 3012
rect 4028 3040 4034 3052
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 4028 3012 4169 3040
rect 4028 3000 4034 3012
rect 4157 3009 4169 3012
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 5534 3000 5540 3052
rect 5592 3040 5598 3052
rect 5813 3043 5871 3049
rect 5813 3040 5825 3043
rect 5592 3012 5825 3040
rect 5592 3000 5598 3012
rect 5813 3009 5825 3012
rect 5859 3040 5871 3043
rect 7282 3040 7288 3052
rect 5859 3012 7288 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 7466 3040 7472 3052
rect 7427 3012 7472 3040
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 11146 3000 11152 3052
rect 11204 3000 11210 3052
rect 11422 3000 11428 3052
rect 11480 3040 11486 3052
rect 12250 3040 12256 3052
rect 11480 3012 12256 3040
rect 11480 3000 11486 3012
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13722 3040 13728 3052
rect 13219 3012 13728 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 13722 3000 13728 3012
rect 13780 3040 13786 3052
rect 13817 3043 13875 3049
rect 13817 3040 13829 3043
rect 13780 3012 13829 3040
rect 13780 3000 13786 3012
rect 13817 3009 13829 3012
rect 13863 3009 13875 3043
rect 13817 3003 13875 3009
rect 2608 2944 3096 2972
rect 3237 2975 3295 2981
rect 2409 2907 2467 2913
rect 2409 2873 2421 2907
rect 2455 2904 2467 2907
rect 2608 2904 2636 2944
rect 3237 2941 3249 2975
rect 3283 2972 3295 2975
rect 3513 2975 3571 2981
rect 3513 2972 3525 2975
rect 3283 2944 3525 2972
rect 3283 2941 3295 2944
rect 3237 2935 3295 2941
rect 3513 2941 3525 2944
rect 3559 2972 3571 2975
rect 4065 2975 4123 2981
rect 4065 2972 4077 2975
rect 3559 2944 4077 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 4065 2941 4077 2944
rect 4111 2972 4123 2975
rect 5994 2972 6000 2984
rect 4111 2944 6000 2972
rect 4111 2941 4123 2944
rect 4065 2935 4123 2941
rect 5994 2932 6000 2944
rect 6052 2932 6058 2984
rect 6273 2975 6331 2981
rect 6273 2941 6285 2975
rect 6319 2972 6331 2975
rect 7190 2972 7196 2984
rect 6319 2944 7196 2972
rect 6319 2941 6331 2944
rect 6273 2935 6331 2941
rect 7190 2932 7196 2944
rect 7248 2972 7254 2984
rect 8110 2972 8116 2984
rect 7248 2944 8116 2972
rect 7248 2932 7254 2944
rect 8110 2932 8116 2944
rect 8168 2932 8174 2984
rect 8202 2932 8208 2984
rect 8260 2972 8266 2984
rect 8662 2981 8668 2984
rect 8389 2975 8447 2981
rect 8389 2972 8401 2975
rect 8260 2944 8401 2972
rect 8260 2932 8266 2944
rect 8389 2941 8401 2944
rect 8435 2941 8447 2975
rect 8656 2972 8668 2981
rect 8623 2944 8668 2972
rect 8389 2935 8447 2941
rect 8656 2935 8668 2944
rect 8662 2932 8668 2935
rect 8720 2932 8726 2984
rect 9766 2932 9772 2984
rect 9824 2932 9830 2984
rect 11238 2972 11244 2984
rect 11199 2944 11244 2972
rect 11238 2932 11244 2944
rect 11296 2932 11302 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 14660 2944 14841 2972
rect 2455 2876 2636 2904
rect 2455 2873 2467 2876
rect 2409 2867 2467 2873
rect 2682 2864 2688 2916
rect 2740 2904 2746 2916
rect 5537 2907 5595 2913
rect 2740 2876 3740 2904
rect 2740 2864 2746 2876
rect 3712 2848 3740 2876
rect 5537 2873 5549 2907
rect 5583 2904 5595 2907
rect 6362 2904 6368 2916
rect 5583 2876 6368 2904
rect 5583 2873 5595 2876
rect 5537 2867 5595 2873
rect 6362 2864 6368 2876
rect 6420 2864 6426 2916
rect 7098 2904 7104 2916
rect 6472 2876 7104 2904
rect 1210 2796 1216 2848
rect 1268 2836 1274 2848
rect 3237 2839 3295 2845
rect 3237 2836 3249 2839
rect 1268 2808 3249 2836
rect 1268 2796 1274 2808
rect 3237 2805 3249 2808
rect 3283 2805 3295 2839
rect 3237 2799 3295 2805
rect 3694 2796 3700 2848
rect 3752 2836 3758 2848
rect 3973 2839 4031 2845
rect 3973 2836 3985 2839
rect 3752 2808 3985 2836
rect 3752 2796 3758 2808
rect 3973 2805 3985 2808
rect 4019 2805 4031 2839
rect 3973 2799 4031 2805
rect 5629 2839 5687 2845
rect 5629 2805 5641 2839
rect 5675 2836 5687 2839
rect 6472 2836 6500 2876
rect 7098 2864 7104 2876
rect 7156 2864 7162 2916
rect 7285 2907 7343 2913
rect 7285 2873 7297 2907
rect 7331 2904 7343 2907
rect 9784 2904 9812 2932
rect 7331 2876 9812 2904
rect 12805 2907 12863 2913
rect 7331 2873 7343 2876
rect 7285 2867 7343 2873
rect 12805 2873 12817 2907
rect 12851 2904 12863 2907
rect 13725 2907 13783 2913
rect 12851 2876 13676 2904
rect 12851 2873 12863 2876
rect 12805 2867 12863 2873
rect 5675 2808 6500 2836
rect 6641 2839 6699 2845
rect 5675 2805 5687 2808
rect 5629 2799 5687 2805
rect 6641 2805 6653 2839
rect 6687 2836 6699 2839
rect 7300 2836 7328 2867
rect 13648 2848 13676 2876
rect 13725 2873 13737 2907
rect 13771 2904 13783 2907
rect 13998 2904 14004 2916
rect 13771 2876 14004 2904
rect 13771 2873 13783 2876
rect 13725 2867 13783 2873
rect 13998 2864 14004 2876
rect 14056 2864 14062 2916
rect 7926 2836 7932 2848
rect 6687 2808 7328 2836
rect 7887 2808 7932 2836
rect 6687 2805 6699 2808
rect 6641 2799 6699 2805
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 8202 2836 8208 2848
rect 8163 2808 8208 2836
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 9766 2836 9772 2848
rect 9727 2808 9772 2836
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 11422 2836 11428 2848
rect 11383 2808 11428 2836
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 11790 2836 11796 2848
rect 11664 2808 11796 2836
rect 11664 2796 11670 2808
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 13262 2836 13268 2848
rect 13223 2808 13268 2836
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 13630 2836 13636 2848
rect 13591 2808 13636 2836
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 14458 2796 14464 2848
rect 14516 2836 14522 2848
rect 14660 2845 14688 2944
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 14918 2932 14924 2984
rect 14976 2972 14982 2984
rect 15096 2975 15154 2981
rect 15096 2972 15108 2975
rect 14976 2944 15108 2972
rect 14976 2932 14982 2944
rect 15096 2941 15108 2944
rect 15142 2972 15154 2975
rect 15378 2972 15384 2984
rect 15142 2944 15384 2972
rect 15142 2941 15154 2944
rect 15096 2935 15154 2941
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 15562 2932 15568 2984
rect 15620 2972 15626 2984
rect 15856 2972 15884 3148
rect 16209 3145 16221 3148
rect 16255 3176 16267 3179
rect 17773 3179 17831 3185
rect 17773 3176 17785 3179
rect 16255 3148 17785 3176
rect 16255 3145 16267 3148
rect 16209 3139 16267 3145
rect 17773 3145 17785 3148
rect 17819 3176 17831 3179
rect 17954 3176 17960 3188
rect 17819 3148 17960 3176
rect 17819 3145 17831 3148
rect 17773 3139 17831 3145
rect 17954 3136 17960 3148
rect 18012 3136 18018 3188
rect 18782 3136 18788 3188
rect 18840 3176 18846 3188
rect 19242 3176 19248 3188
rect 18840 3148 19248 3176
rect 18840 3136 18846 3148
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 19613 3179 19671 3185
rect 19613 3145 19625 3179
rect 19659 3176 19671 3179
rect 20714 3176 20720 3188
rect 19659 3148 20720 3176
rect 19659 3145 19671 3148
rect 19613 3139 19671 3145
rect 20714 3136 20720 3148
rect 20772 3136 20778 3188
rect 21177 3179 21235 3185
rect 21177 3145 21189 3179
rect 21223 3176 21235 3179
rect 22002 3176 22008 3188
rect 21223 3148 22008 3176
rect 21223 3145 21235 3148
rect 21177 3139 21235 3145
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 22278 3176 22284 3188
rect 22239 3148 22284 3176
rect 22278 3136 22284 3148
rect 22336 3136 22342 3188
rect 23658 3176 23664 3188
rect 23619 3148 23664 3176
rect 23658 3136 23664 3148
rect 23716 3136 23722 3188
rect 24670 3176 24676 3188
rect 24631 3148 24676 3176
rect 24670 3136 24676 3148
rect 24728 3136 24734 3188
rect 16850 3068 16856 3120
rect 16908 3108 16914 3120
rect 17129 3111 17187 3117
rect 17129 3108 17141 3111
rect 16908 3080 17141 3108
rect 16908 3068 16914 3080
rect 17129 3077 17141 3080
rect 17175 3077 17187 3111
rect 17129 3071 17187 3077
rect 17972 3040 18000 3136
rect 19978 3068 19984 3120
rect 20036 3108 20042 3120
rect 23477 3111 23535 3117
rect 20036 3080 20208 3108
rect 20036 3068 20042 3080
rect 18601 3043 18659 3049
rect 18601 3040 18613 3043
rect 17972 3012 18613 3040
rect 18601 3009 18613 3012
rect 18647 3040 18659 3043
rect 19061 3043 19119 3049
rect 19061 3040 19073 3043
rect 18647 3012 19073 3040
rect 18647 3009 18659 3012
rect 18601 3003 18659 3009
rect 19061 3009 19073 3012
rect 19107 3009 19119 3043
rect 20070 3040 20076 3052
rect 20031 3012 20076 3040
rect 19061 3003 19119 3009
rect 20070 3000 20076 3012
rect 20128 3000 20134 3052
rect 20180 3049 20208 3080
rect 23477 3077 23489 3111
rect 23523 3108 23535 3111
rect 23566 3108 23572 3120
rect 23523 3080 23572 3108
rect 23523 3077 23535 3080
rect 23477 3071 23535 3077
rect 23566 3068 23572 3080
rect 23624 3108 23630 3120
rect 24210 3108 24216 3120
rect 23624 3080 24216 3108
rect 23624 3068 23630 3080
rect 24210 3068 24216 3080
rect 24268 3068 24274 3120
rect 20165 3043 20223 3049
rect 20165 3009 20177 3043
rect 20211 3009 20223 3043
rect 21726 3040 21732 3052
rect 21687 3012 21732 3040
rect 20165 3003 20223 3009
rect 21726 3000 21732 3012
rect 21784 3040 21790 3052
rect 22925 3043 22983 3049
rect 22925 3040 22937 3043
rect 21784 3012 22937 3040
rect 21784 3000 21790 3012
rect 22925 3009 22937 3012
rect 22971 3009 22983 3043
rect 22925 3003 22983 3009
rect 24026 3000 24032 3052
rect 24084 3040 24090 3052
rect 24121 3043 24179 3049
rect 24121 3040 24133 3043
rect 24084 3012 24133 3040
rect 24084 3000 24090 3012
rect 24121 3009 24133 3012
rect 24167 3009 24179 3043
rect 24302 3040 24308 3052
rect 24263 3012 24308 3040
rect 24121 3003 24179 3009
rect 24302 3000 24308 3012
rect 24360 3000 24366 3052
rect 26234 3040 26240 3052
rect 26195 3012 26240 3040
rect 26234 3000 26240 3012
rect 26292 3000 26298 3052
rect 15620 2944 15884 2972
rect 16853 2975 16911 2981
rect 15620 2932 15626 2944
rect 16853 2941 16865 2975
rect 16899 2972 16911 2975
rect 17034 2972 17040 2984
rect 16899 2944 17040 2972
rect 16899 2941 16911 2944
rect 16853 2935 16911 2941
rect 17034 2932 17040 2944
rect 17092 2932 17098 2984
rect 17586 2932 17592 2984
rect 17644 2972 17650 2984
rect 18138 2972 18144 2984
rect 17644 2944 18144 2972
rect 17644 2932 17650 2944
rect 18138 2932 18144 2944
rect 18196 2932 18202 2984
rect 18414 2972 18420 2984
rect 18375 2944 18420 2972
rect 18414 2932 18420 2944
rect 18472 2932 18478 2984
rect 18506 2932 18512 2984
rect 18564 2972 18570 2984
rect 19521 2975 19579 2981
rect 18564 2944 18609 2972
rect 18564 2932 18570 2944
rect 19521 2941 19533 2975
rect 19567 2972 19579 2975
rect 19981 2975 20039 2981
rect 19981 2972 19993 2975
rect 19567 2944 19993 2972
rect 19567 2941 19579 2944
rect 19521 2935 19579 2941
rect 19981 2941 19993 2944
rect 20027 2972 20039 2975
rect 20806 2972 20812 2984
rect 20027 2944 20812 2972
rect 20027 2941 20039 2944
rect 19981 2935 20039 2941
rect 20806 2932 20812 2944
rect 20864 2932 20870 2984
rect 21266 2972 21272 2984
rect 20916 2944 21272 2972
rect 18156 2904 18184 2932
rect 18598 2904 18604 2916
rect 18156 2876 18604 2904
rect 18598 2864 18604 2876
rect 18656 2864 18662 2916
rect 20714 2904 20720 2916
rect 20675 2876 20720 2904
rect 20714 2864 20720 2876
rect 20772 2904 20778 2916
rect 20916 2904 20944 2944
rect 21266 2932 21272 2944
rect 21324 2932 21330 2984
rect 21637 2975 21695 2981
rect 21637 2941 21649 2975
rect 21683 2972 21695 2975
rect 22278 2972 22284 2984
rect 21683 2944 22284 2972
rect 21683 2941 21695 2944
rect 21637 2935 21695 2941
rect 22278 2932 22284 2944
rect 22336 2932 22342 2984
rect 22462 2932 22468 2984
rect 22520 2972 22526 2984
rect 23566 2972 23572 2984
rect 22520 2944 23572 2972
rect 22520 2932 22526 2944
rect 23566 2932 23572 2944
rect 23624 2932 23630 2984
rect 23750 2932 23756 2984
rect 23808 2972 23814 2984
rect 24670 2972 24676 2984
rect 23808 2944 24676 2972
rect 23808 2932 23814 2944
rect 24670 2932 24676 2944
rect 24728 2932 24734 2984
rect 25225 2975 25283 2981
rect 25225 2941 25237 2975
rect 25271 2972 25283 2975
rect 25774 2972 25780 2984
rect 25271 2944 25780 2972
rect 25271 2941 25283 2944
rect 25225 2935 25283 2941
rect 25774 2932 25780 2944
rect 25832 2932 25838 2984
rect 20772 2876 20944 2904
rect 20772 2864 20778 2876
rect 20990 2864 20996 2916
rect 21048 2904 21054 2916
rect 21085 2907 21143 2913
rect 21085 2904 21097 2907
rect 21048 2876 21097 2904
rect 21048 2864 21054 2876
rect 21085 2873 21097 2876
rect 21131 2904 21143 2907
rect 21545 2907 21603 2913
rect 21545 2904 21557 2907
rect 21131 2876 21557 2904
rect 21131 2873 21143 2876
rect 21085 2867 21143 2873
rect 21545 2873 21557 2876
rect 21591 2873 21603 2907
rect 25682 2904 25688 2916
rect 21545 2867 21603 2873
rect 23768 2876 25688 2904
rect 23768 2848 23796 2876
rect 25682 2864 25688 2876
rect 25740 2864 25746 2916
rect 14645 2839 14703 2845
rect 14645 2836 14657 2839
rect 14516 2808 14657 2836
rect 14516 2796 14522 2808
rect 14645 2805 14657 2808
rect 14691 2805 14703 2839
rect 18046 2836 18052 2848
rect 18007 2808 18052 2836
rect 14645 2799 14703 2805
rect 18046 2796 18052 2808
rect 18104 2796 18110 2848
rect 21358 2796 21364 2848
rect 21416 2836 21422 2848
rect 22649 2839 22707 2845
rect 22649 2836 22661 2839
rect 21416 2808 22661 2836
rect 21416 2796 21422 2808
rect 22649 2805 22661 2808
rect 22695 2836 22707 2839
rect 23106 2836 23112 2848
rect 22695 2808 23112 2836
rect 22695 2805 22707 2808
rect 22649 2799 22707 2805
rect 23106 2796 23112 2808
rect 23164 2796 23170 2848
rect 23750 2796 23756 2848
rect 23808 2796 23814 2848
rect 24029 2839 24087 2845
rect 24029 2805 24041 2839
rect 24075 2836 24087 2839
rect 24210 2836 24216 2848
rect 24075 2808 24216 2836
rect 24075 2805 24087 2808
rect 24029 2799 24087 2805
rect 24210 2796 24216 2808
rect 24268 2796 24274 2848
rect 25038 2836 25044 2848
rect 24999 2808 25044 2836
rect 25038 2796 25044 2808
rect 25096 2796 25102 2848
rect 25130 2796 25136 2848
rect 25188 2836 25194 2848
rect 25409 2839 25467 2845
rect 25409 2836 25421 2839
rect 25188 2808 25421 2836
rect 25188 2796 25194 2808
rect 25409 2805 25421 2808
rect 25455 2805 25467 2839
rect 25409 2799 25467 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 2222 2592 2228 2644
rect 2280 2632 2286 2644
rect 2409 2635 2467 2641
rect 2409 2632 2421 2635
rect 2280 2604 2421 2632
rect 2280 2592 2286 2604
rect 2409 2601 2421 2604
rect 2455 2601 2467 2635
rect 2866 2632 2872 2644
rect 2827 2604 2872 2632
rect 2409 2595 2467 2601
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 5721 2635 5779 2641
rect 5721 2632 5733 2635
rect 5592 2604 5733 2632
rect 5592 2592 5598 2604
rect 5721 2601 5733 2604
rect 5767 2601 5779 2635
rect 5721 2595 5779 2601
rect 6546 2592 6552 2644
rect 6604 2632 6610 2644
rect 6641 2635 6699 2641
rect 6641 2632 6653 2635
rect 6604 2604 6653 2632
rect 6604 2592 6610 2604
rect 6641 2601 6653 2604
rect 6687 2601 6699 2635
rect 8294 2632 8300 2644
rect 8255 2604 8300 2632
rect 6641 2595 6699 2601
rect 2774 2524 2780 2576
rect 2832 2564 2838 2576
rect 3694 2564 3700 2576
rect 2832 2536 2877 2564
rect 3655 2536 3700 2564
rect 2832 2524 2838 2536
rect 3694 2524 3700 2536
rect 3752 2524 3758 2576
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 1946 2496 1952 2508
rect 1443 2468 1952 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2496 4399 2499
rect 4430 2496 4436 2508
rect 4387 2468 4436 2496
rect 4387 2465 4399 2468
rect 4341 2459 4399 2465
rect 4430 2456 4436 2468
rect 4488 2456 4494 2508
rect 4608 2499 4666 2505
rect 4608 2465 4620 2499
rect 4654 2496 4666 2499
rect 5074 2496 5080 2508
rect 4654 2468 5080 2496
rect 4654 2465 4666 2468
rect 4608 2459 4666 2465
rect 5074 2456 5080 2468
rect 5132 2496 5138 2508
rect 6273 2499 6331 2505
rect 6273 2496 6285 2499
rect 5132 2468 6285 2496
rect 5132 2456 5138 2468
rect 6273 2465 6285 2468
rect 6319 2465 6331 2499
rect 6656 2496 6684 2595
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 14277 2635 14335 2641
rect 14277 2601 14289 2635
rect 14323 2632 14335 2635
rect 14550 2632 14556 2644
rect 14323 2604 14556 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 14918 2632 14924 2644
rect 14879 2604 14924 2632
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 18049 2635 18107 2641
rect 18049 2601 18061 2635
rect 18095 2632 18107 2635
rect 18785 2635 18843 2641
rect 18785 2632 18797 2635
rect 18095 2604 18797 2632
rect 18095 2601 18107 2604
rect 18049 2595 18107 2601
rect 18785 2601 18797 2604
rect 18831 2632 18843 2635
rect 18966 2632 18972 2644
rect 18831 2604 18972 2632
rect 18831 2601 18843 2604
rect 18785 2595 18843 2601
rect 18966 2592 18972 2604
rect 19024 2592 19030 2644
rect 21177 2635 21235 2641
rect 21177 2601 21189 2635
rect 21223 2632 21235 2635
rect 22002 2632 22008 2644
rect 21223 2604 22008 2632
rect 21223 2601 21235 2604
rect 21177 2595 21235 2601
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 22278 2632 22284 2644
rect 22239 2604 22284 2632
rect 22278 2592 22284 2604
rect 22336 2592 22342 2644
rect 23934 2592 23940 2644
rect 23992 2632 23998 2644
rect 24029 2635 24087 2641
rect 24029 2632 24041 2635
rect 23992 2604 24041 2632
rect 23992 2592 23998 2604
rect 24029 2601 24041 2604
rect 24075 2601 24087 2635
rect 24029 2595 24087 2601
rect 7184 2567 7242 2573
rect 7184 2533 7196 2567
rect 7230 2564 7242 2567
rect 7926 2564 7932 2576
rect 7230 2536 7932 2564
rect 7230 2533 7242 2536
rect 7184 2527 7242 2533
rect 7926 2524 7932 2536
rect 7984 2524 7990 2576
rect 10036 2567 10094 2573
rect 10036 2533 10048 2567
rect 10082 2564 10094 2567
rect 10870 2564 10876 2576
rect 10082 2536 10876 2564
rect 10082 2533 10094 2536
rect 10036 2527 10094 2533
rect 10870 2524 10876 2536
rect 10928 2524 10934 2576
rect 12069 2567 12127 2573
rect 12069 2533 12081 2567
rect 12115 2564 12127 2567
rect 13164 2567 13222 2573
rect 13164 2564 13176 2567
rect 12115 2536 13176 2564
rect 12115 2533 12127 2536
rect 12069 2527 12127 2533
rect 13164 2533 13176 2536
rect 13210 2564 13222 2567
rect 13722 2564 13728 2576
rect 13210 2536 13728 2564
rect 13210 2533 13222 2536
rect 13164 2527 13222 2533
rect 13722 2524 13728 2536
rect 13780 2524 13786 2576
rect 15562 2524 15568 2576
rect 15620 2564 15626 2576
rect 15718 2567 15776 2573
rect 15718 2564 15730 2567
rect 15620 2536 15730 2564
rect 15620 2524 15626 2536
rect 15718 2533 15730 2536
rect 15764 2533 15776 2567
rect 15718 2527 15776 2533
rect 18138 2524 18144 2576
rect 18196 2564 18202 2576
rect 18196 2536 18920 2564
rect 18196 2524 18202 2536
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6656 2468 6929 2496
rect 6273 2459 6331 2465
rect 6917 2465 6929 2468
rect 6963 2496 6975 2499
rect 8202 2496 8208 2508
rect 6963 2468 8208 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 8202 2456 8208 2468
rect 8260 2496 8266 2508
rect 8849 2499 8907 2505
rect 8849 2496 8861 2499
rect 8260 2468 8861 2496
rect 8260 2456 8266 2468
rect 8849 2465 8861 2468
rect 8895 2496 8907 2499
rect 9493 2499 9551 2505
rect 9493 2496 9505 2499
rect 8895 2468 9505 2496
rect 8895 2465 8907 2468
rect 8849 2459 8907 2465
rect 9493 2465 9505 2468
rect 9539 2496 9551 2499
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9539 2468 9781 2496
rect 9539 2465 9551 2468
rect 9493 2459 9551 2465
rect 9769 2465 9781 2468
rect 9815 2496 9827 2499
rect 11790 2496 11796 2508
rect 9815 2468 11796 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 11790 2456 11796 2468
rect 11848 2496 11854 2508
rect 12345 2499 12403 2505
rect 12345 2496 12357 2499
rect 11848 2468 12357 2496
rect 11848 2456 11854 2468
rect 12345 2465 12357 2468
rect 12391 2496 12403 2499
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 12391 2468 12909 2496
rect 12391 2465 12403 2468
rect 12345 2459 12403 2465
rect 12897 2465 12909 2468
rect 12943 2496 12955 2499
rect 12986 2496 12992 2508
rect 12943 2468 12992 2496
rect 12943 2465 12955 2468
rect 12897 2459 12955 2465
rect 12986 2456 12992 2468
rect 13044 2496 13050 2508
rect 14458 2496 14464 2508
rect 13044 2468 14464 2496
rect 13044 2456 13050 2468
rect 14458 2456 14464 2468
rect 14516 2496 14522 2508
rect 15197 2499 15255 2505
rect 15197 2496 15209 2499
rect 14516 2468 15209 2496
rect 14516 2456 14522 2468
rect 15197 2465 15209 2468
rect 15243 2496 15255 2499
rect 15286 2496 15292 2508
rect 15243 2468 15292 2496
rect 15243 2465 15255 2468
rect 15197 2459 15255 2465
rect 15286 2456 15292 2468
rect 15344 2496 15350 2508
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15344 2468 15485 2496
rect 15344 2456 15350 2468
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 15473 2459 15531 2465
rect 18693 2499 18751 2505
rect 18693 2465 18705 2499
rect 18739 2465 18751 2499
rect 18693 2459 18751 2465
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2428 2375 2431
rect 2961 2431 3019 2437
rect 2961 2428 2973 2431
rect 2363 2400 2973 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 2961 2397 2973 2400
rect 3007 2428 3019 2431
rect 4246 2428 4252 2440
rect 3007 2400 4252 2428
rect 3007 2397 3019 2400
rect 2961 2391 3019 2397
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 18708 2372 18736 2459
rect 18892 2437 18920 2536
rect 20898 2524 20904 2576
rect 20956 2564 20962 2576
rect 21637 2567 21695 2573
rect 21637 2564 21649 2567
rect 20956 2536 21649 2564
rect 20956 2524 20962 2536
rect 21637 2533 21649 2536
rect 21683 2564 21695 2567
rect 22554 2564 22560 2576
rect 21683 2536 22560 2564
rect 21683 2533 21695 2536
rect 21637 2527 21695 2533
rect 22554 2524 22560 2536
rect 22612 2524 22618 2576
rect 23474 2524 23480 2576
rect 23532 2564 23538 2576
rect 24397 2567 24455 2573
rect 24397 2564 24409 2567
rect 23532 2536 24409 2564
rect 23532 2524 23538 2536
rect 24397 2533 24409 2536
rect 24443 2564 24455 2567
rect 24762 2564 24768 2576
rect 24443 2536 24768 2564
rect 24443 2533 24455 2536
rect 24397 2527 24455 2533
rect 24762 2524 24768 2536
rect 24820 2524 24826 2576
rect 19705 2499 19763 2505
rect 19705 2465 19717 2499
rect 19751 2496 19763 2499
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19751 2468 19901 2496
rect 19751 2465 19763 2468
rect 19705 2459 19763 2465
rect 19889 2465 19901 2468
rect 19935 2496 19947 2499
rect 20070 2496 20076 2508
rect 19935 2468 20076 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 20070 2456 20076 2468
rect 20128 2456 20134 2508
rect 21545 2499 21603 2505
rect 21545 2465 21557 2499
rect 21591 2465 21603 2499
rect 22738 2496 22744 2508
rect 22699 2468 22744 2496
rect 21545 2459 21603 2465
rect 18877 2431 18935 2437
rect 18877 2397 18889 2431
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 17681 2363 17739 2369
rect 17681 2360 17693 2363
rect 16684 2332 17693 2360
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 1946 2292 1952 2304
rect 1907 2264 1952 2292
rect 1946 2252 1952 2264
rect 2004 2252 2010 2304
rect 11149 2295 11207 2301
rect 11149 2261 11161 2295
rect 11195 2292 11207 2295
rect 11238 2292 11244 2304
rect 11195 2264 11244 2292
rect 11195 2261 11207 2264
rect 11149 2255 11207 2261
rect 11238 2252 11244 2264
rect 11296 2252 11302 2304
rect 14550 2252 14556 2304
rect 14608 2292 14614 2304
rect 16684 2292 16712 2332
rect 17681 2329 17693 2332
rect 17727 2360 17739 2363
rect 18690 2360 18696 2372
rect 17727 2332 18696 2360
rect 17727 2329 17739 2332
rect 17681 2323 17739 2329
rect 18690 2320 18696 2332
rect 18748 2320 18754 2372
rect 20530 2360 20536 2372
rect 20491 2332 20536 2360
rect 20530 2320 20536 2332
rect 20588 2360 20594 2372
rect 21560 2360 21588 2459
rect 22738 2456 22744 2468
rect 22796 2456 22802 2508
rect 23014 2456 23020 2508
rect 23072 2496 23078 2508
rect 23385 2499 23443 2505
rect 23385 2496 23397 2499
rect 23072 2468 23397 2496
rect 23072 2456 23078 2468
rect 23385 2465 23397 2468
rect 23431 2496 23443 2499
rect 23661 2499 23719 2505
rect 23661 2496 23673 2499
rect 23431 2468 23673 2496
rect 23431 2465 23443 2468
rect 23385 2459 23443 2465
rect 23661 2465 23673 2468
rect 23707 2496 23719 2499
rect 24302 2496 24308 2508
rect 23707 2468 24308 2496
rect 23707 2465 23719 2468
rect 23661 2459 23719 2465
rect 24302 2456 24308 2468
rect 24360 2456 24366 2508
rect 24486 2496 24492 2508
rect 24447 2468 24492 2496
rect 24486 2456 24492 2468
rect 24544 2456 24550 2508
rect 24670 2456 24676 2508
rect 24728 2496 24734 2508
rect 25593 2499 25651 2505
rect 25593 2496 25605 2499
rect 24728 2468 25605 2496
rect 24728 2456 24734 2468
rect 25593 2465 25605 2468
rect 25639 2496 25651 2499
rect 26053 2499 26111 2505
rect 26053 2496 26065 2499
rect 25639 2468 26065 2496
rect 25639 2465 25651 2468
rect 25593 2459 25651 2465
rect 26053 2465 26065 2468
rect 26099 2465 26111 2499
rect 26418 2496 26424 2508
rect 26379 2468 26424 2496
rect 26053 2459 26111 2465
rect 26418 2456 26424 2468
rect 26476 2456 26482 2508
rect 21726 2428 21732 2440
rect 21687 2400 21732 2428
rect 21726 2388 21732 2400
rect 21784 2428 21790 2440
rect 22557 2431 22615 2437
rect 22557 2428 22569 2431
rect 21784 2400 22569 2428
rect 21784 2388 21790 2400
rect 22557 2397 22569 2400
rect 22603 2397 22615 2431
rect 22557 2391 22615 2397
rect 22922 2388 22928 2440
rect 22980 2428 22986 2440
rect 24578 2428 24584 2440
rect 22980 2400 23060 2428
rect 24539 2400 24584 2428
rect 22980 2388 22986 2400
rect 20588 2332 21588 2360
rect 23032 2360 23060 2400
rect 24578 2388 24584 2400
rect 24636 2428 24642 2440
rect 25041 2431 25099 2437
rect 25041 2428 25053 2431
rect 24636 2400 25053 2428
rect 24636 2388 24642 2400
rect 25041 2397 25053 2400
rect 25087 2397 25099 2431
rect 25041 2391 25099 2397
rect 25409 2363 25467 2369
rect 25409 2360 25421 2363
rect 23032 2332 25421 2360
rect 20588 2320 20594 2332
rect 25409 2329 25421 2332
rect 25455 2329 25467 2363
rect 25409 2323 25467 2329
rect 16850 2292 16856 2304
rect 14608 2264 16712 2292
rect 16811 2264 16856 2292
rect 14608 2252 14614 2264
rect 16850 2252 16856 2264
rect 16908 2252 16914 2304
rect 18322 2292 18328 2304
rect 18283 2264 18328 2292
rect 18322 2252 18328 2264
rect 18380 2252 18386 2304
rect 19886 2252 19892 2304
rect 19944 2292 19950 2304
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 19944 2264 20085 2292
rect 19944 2252 19950 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 20898 2292 20904 2304
rect 20859 2264 20904 2292
rect 20073 2255 20131 2261
rect 20898 2252 20904 2264
rect 20956 2252 20962 2304
rect 22922 2292 22928 2304
rect 22883 2264 22928 2292
rect 22922 2252 22928 2264
rect 22980 2252 22986 2304
rect 24762 2252 24768 2304
rect 24820 2292 24826 2304
rect 25498 2292 25504 2304
rect 24820 2264 25504 2292
rect 24820 2252 24826 2264
rect 25498 2252 25504 2264
rect 25556 2252 25562 2304
rect 25774 2292 25780 2304
rect 25735 2264 25780 2292
rect 25774 2252 25780 2264
rect 25832 2252 25838 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 11330 2048 11336 2100
rect 11388 2088 11394 2100
rect 17402 2088 17408 2100
rect 11388 2060 17408 2088
rect 11388 2048 11394 2060
rect 17402 2048 17408 2060
rect 17460 2048 17466 2100
rect 14642 1844 14648 1896
rect 14700 1884 14706 1896
rect 17494 1884 17500 1896
rect 14700 1856 17500 1884
rect 14700 1844 14706 1856
rect 17494 1844 17500 1856
rect 17552 1844 17558 1896
rect 5626 1640 5632 1692
rect 5684 1680 5690 1692
rect 6638 1680 6644 1692
rect 5684 1652 6644 1680
rect 5684 1640 5690 1652
rect 6638 1640 6644 1652
rect 6696 1640 6702 1692
rect 15102 1572 15108 1624
rect 15160 1612 15166 1624
rect 17954 1612 17960 1624
rect 15160 1584 17960 1612
rect 15160 1572 15166 1584
rect 17954 1572 17960 1584
rect 18012 1572 18018 1624
rect 24946 552 24952 604
rect 25004 592 25010 604
rect 25406 592 25412 604
rect 25004 564 25412 592
rect 25004 552 25010 564
rect 25406 552 25412 564
rect 25464 552 25470 604
rect 14826 212 14832 264
rect 14884 252 14890 264
rect 18138 252 18144 264
rect 14884 224 18144 252
rect 14884 212 14890 224
rect 18138 212 18144 224
rect 18196 212 18202 264
<< via1 >>
rect 20720 26800 20772 26852
rect 23756 26800 23808 26852
rect 18512 26664 18564 26716
rect 24768 26664 24820 26716
rect 20352 26528 20404 26580
rect 13544 26460 13596 26512
rect 23296 26460 23348 26512
rect 7380 26120 7432 26172
rect 20444 26256 20496 26308
rect 23756 26256 23808 26308
rect 10784 26188 10836 26240
rect 21364 26188 21416 26240
rect 25044 26120 25096 26172
rect 2688 26095 2740 26104
rect 2688 26061 2697 26095
rect 2697 26061 2731 26095
rect 2731 26061 2740 26095
rect 2688 26052 2740 26061
rect 5172 26052 5224 26104
rect 11520 26052 11572 26104
rect 10876 25984 10928 26036
rect 22928 26052 22980 26104
rect 18420 25984 18472 26036
rect 26608 25984 26660 26036
rect 5080 25916 5132 25968
rect 16948 25916 17000 25968
rect 18236 25916 18288 25968
rect 18328 25916 18380 25968
rect 19248 25916 19300 25968
rect 20904 25916 20956 25968
rect 20996 25916 21048 25968
rect 22744 25916 22796 25968
rect 6828 25848 6880 25900
rect 11704 25848 11756 25900
rect 23756 25848 23808 25900
rect 11336 25780 11388 25832
rect 15568 25780 15620 25832
rect 9956 25644 10008 25696
rect 18880 25712 18932 25764
rect 19984 25780 20036 25832
rect 20720 25780 20772 25832
rect 24584 25712 24636 25764
rect 16672 25644 16724 25696
rect 23480 25644 23532 25696
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5540 25440 5592 25492
rect 9496 25440 9548 25492
rect 9956 25483 10008 25492
rect 9956 25449 9965 25483
rect 9965 25449 9999 25483
rect 9999 25449 10008 25483
rect 9956 25440 10008 25449
rect 1492 25372 1544 25424
rect 5264 25372 5316 25424
rect 11704 25440 11756 25492
rect 12808 25440 12860 25492
rect 12900 25440 12952 25492
rect 14188 25440 14240 25492
rect 2136 25304 2188 25356
rect 2504 25347 2556 25356
rect 2504 25313 2513 25347
rect 2513 25313 2547 25347
rect 2547 25313 2556 25347
rect 2504 25304 2556 25313
rect 4068 25347 4120 25356
rect 4068 25313 4077 25347
rect 4077 25313 4111 25347
rect 4111 25313 4120 25347
rect 4068 25304 4120 25313
rect 6552 25304 6604 25356
rect 9772 25347 9824 25356
rect 9772 25313 9781 25347
rect 9781 25313 9815 25347
rect 9815 25313 9824 25347
rect 9772 25304 9824 25313
rect 11336 25347 11388 25356
rect 2228 25236 2280 25288
rect 4344 25168 4396 25220
rect 5172 25168 5224 25220
rect 572 25100 624 25152
rect 2044 25143 2096 25152
rect 2044 25109 2053 25143
rect 2053 25109 2087 25143
rect 2087 25109 2096 25143
rect 2044 25100 2096 25109
rect 2320 25143 2372 25152
rect 2320 25109 2329 25143
rect 2329 25109 2363 25143
rect 2363 25109 2372 25143
rect 2320 25100 2372 25109
rect 2872 25100 2924 25152
rect 3148 25143 3200 25152
rect 3148 25109 3157 25143
rect 3157 25109 3191 25143
rect 3191 25109 3200 25143
rect 3148 25100 3200 25109
rect 3424 25143 3476 25152
rect 3424 25109 3433 25143
rect 3433 25109 3467 25143
rect 3467 25109 3476 25143
rect 3424 25100 3476 25109
rect 3700 25100 3752 25152
rect 4712 25143 4764 25152
rect 4712 25109 4721 25143
rect 4721 25109 4755 25143
rect 4755 25109 4764 25143
rect 4712 25100 4764 25109
rect 4988 25143 5040 25152
rect 4988 25109 4997 25143
rect 4997 25109 5031 25143
rect 5031 25109 5040 25143
rect 4988 25100 5040 25109
rect 6460 25100 6512 25152
rect 7932 25168 7984 25220
rect 11336 25313 11345 25347
rect 11345 25313 11379 25347
rect 11379 25313 11388 25347
rect 11336 25304 11388 25313
rect 11060 25236 11112 25288
rect 14096 25372 14148 25424
rect 15476 25440 15528 25492
rect 19524 25440 19576 25492
rect 19984 25440 20036 25492
rect 20628 25440 20680 25492
rect 23020 25440 23072 25492
rect 21272 25372 21324 25424
rect 12072 25304 12124 25356
rect 12900 25236 12952 25288
rect 13084 25279 13136 25288
rect 13084 25245 13093 25279
rect 13093 25245 13127 25279
rect 13127 25245 13136 25279
rect 13084 25236 13136 25245
rect 14004 25236 14056 25288
rect 14372 25304 14424 25356
rect 15936 25304 15988 25356
rect 16856 25304 16908 25356
rect 16948 25304 17000 25356
rect 17500 25304 17552 25356
rect 18604 25304 18656 25356
rect 18696 25347 18748 25356
rect 18696 25313 18705 25347
rect 18705 25313 18739 25347
rect 18739 25313 18748 25347
rect 18696 25304 18748 25313
rect 19064 25304 19116 25356
rect 20720 25304 20772 25356
rect 21180 25347 21232 25356
rect 21180 25313 21189 25347
rect 21189 25313 21223 25347
rect 21223 25313 21232 25347
rect 21180 25304 21232 25313
rect 22376 25304 22428 25356
rect 24216 25304 24268 25356
rect 17316 25279 17368 25288
rect 17316 25245 17325 25279
rect 17325 25245 17359 25279
rect 17359 25245 17368 25279
rect 17316 25236 17368 25245
rect 7656 25100 7708 25152
rect 7840 25100 7892 25152
rect 18972 25279 19024 25288
rect 18972 25245 18981 25279
rect 18981 25245 19015 25279
rect 19015 25245 19024 25279
rect 18972 25236 19024 25245
rect 19248 25236 19300 25288
rect 23204 25236 23256 25288
rect 8760 25100 8812 25152
rect 9772 25100 9824 25152
rect 11980 25143 12032 25152
rect 11980 25109 11989 25143
rect 11989 25109 12023 25143
rect 12023 25109 12032 25143
rect 11980 25100 12032 25109
rect 12440 25143 12492 25152
rect 12440 25109 12449 25143
rect 12449 25109 12483 25143
rect 12483 25109 12492 25143
rect 12440 25100 12492 25109
rect 12992 25100 13044 25152
rect 13176 25100 13228 25152
rect 14832 25143 14884 25152
rect 14832 25109 14841 25143
rect 14841 25109 14875 25143
rect 14875 25109 14884 25143
rect 14832 25100 14884 25109
rect 15292 25100 15344 25152
rect 16672 25143 16724 25152
rect 16672 25109 16681 25143
rect 16681 25109 16715 25143
rect 16715 25109 16724 25143
rect 16672 25100 16724 25109
rect 17316 25100 17368 25152
rect 18144 25143 18196 25152
rect 18144 25109 18153 25143
rect 18153 25109 18187 25143
rect 18187 25109 18196 25143
rect 18144 25100 18196 25109
rect 18236 25100 18288 25152
rect 18788 25100 18840 25152
rect 21732 25143 21784 25152
rect 21732 25109 21741 25143
rect 21741 25109 21775 25143
rect 21775 25109 21784 25143
rect 21732 25100 21784 25109
rect 26056 25100 26108 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 6736 24896 6788 24948
rect 3424 24828 3476 24880
rect 4712 24828 4764 24880
rect 7932 24828 7984 24880
rect 11060 24871 11112 24880
rect 1584 24692 1636 24744
rect 2412 24692 2464 24744
rect 4988 24692 5040 24744
rect 7472 24692 7524 24744
rect 10232 24803 10284 24812
rect 10232 24769 10241 24803
rect 10241 24769 10275 24803
rect 10275 24769 10284 24803
rect 10232 24760 10284 24769
rect 11060 24837 11069 24871
rect 11069 24837 11103 24871
rect 11103 24837 11112 24871
rect 11060 24828 11112 24837
rect 11520 24828 11572 24880
rect 12256 24760 12308 24812
rect 9496 24692 9548 24744
rect 12348 24692 12400 24744
rect 13084 24896 13136 24948
rect 14096 24896 14148 24948
rect 12992 24828 13044 24880
rect 15660 24828 15712 24880
rect 15752 24828 15804 24880
rect 18880 24828 18932 24880
rect 13452 24760 13504 24812
rect 14004 24760 14056 24812
rect 14832 24803 14884 24812
rect 14832 24769 14841 24803
rect 14841 24769 14875 24803
rect 14875 24769 14884 24803
rect 14832 24760 14884 24769
rect 14372 24692 14424 24744
rect 14464 24692 14516 24744
rect 17316 24760 17368 24812
rect 17408 24760 17460 24812
rect 18236 24760 18288 24812
rect 18604 24803 18656 24812
rect 18604 24769 18613 24803
rect 18613 24769 18647 24803
rect 18647 24769 18656 24803
rect 18604 24760 18656 24769
rect 18972 24760 19024 24812
rect 20628 24828 20680 24880
rect 24768 24828 24820 24880
rect 20352 24760 20404 24812
rect 20720 24803 20772 24812
rect 20720 24769 20729 24803
rect 20729 24769 20763 24803
rect 20763 24769 20772 24803
rect 20720 24760 20772 24769
rect 18144 24692 18196 24744
rect 19984 24735 20036 24744
rect 19984 24701 19993 24735
rect 19993 24701 20027 24735
rect 20027 24701 20036 24735
rect 19984 24692 20036 24701
rect 21732 24692 21784 24744
rect 1400 24556 1452 24608
rect 2136 24556 2188 24608
rect 2412 24556 2464 24608
rect 3056 24556 3108 24608
rect 3792 24556 3844 24608
rect 4068 24599 4120 24608
rect 4068 24565 4077 24599
rect 4077 24565 4111 24599
rect 4111 24565 4120 24599
rect 4068 24556 4120 24565
rect 6000 24556 6052 24608
rect 6552 24599 6604 24608
rect 6552 24565 6561 24599
rect 6561 24565 6595 24599
rect 6595 24565 6604 24599
rect 6552 24556 6604 24565
rect 7932 24599 7984 24608
rect 7932 24565 7941 24599
rect 7941 24565 7975 24599
rect 7975 24565 7984 24599
rect 7932 24556 7984 24565
rect 8116 24599 8168 24608
rect 8116 24565 8125 24599
rect 8125 24565 8159 24599
rect 8159 24565 8168 24599
rect 8116 24556 8168 24565
rect 8208 24556 8260 24608
rect 8760 24556 8812 24608
rect 9496 24599 9548 24608
rect 9496 24565 9505 24599
rect 9505 24565 9539 24599
rect 9539 24565 9548 24599
rect 9496 24556 9548 24565
rect 9680 24599 9732 24608
rect 9680 24565 9689 24599
rect 9689 24565 9723 24599
rect 9723 24565 9732 24599
rect 9680 24556 9732 24565
rect 11428 24599 11480 24608
rect 11428 24565 11437 24599
rect 11437 24565 11471 24599
rect 11471 24565 11480 24599
rect 11428 24556 11480 24565
rect 12256 24599 12308 24608
rect 12256 24565 12265 24599
rect 12265 24565 12299 24599
rect 12299 24565 12308 24599
rect 12256 24556 12308 24565
rect 12716 24556 12768 24608
rect 13452 24556 13504 24608
rect 14556 24556 14608 24608
rect 14924 24624 14976 24676
rect 16304 24667 16356 24676
rect 16304 24633 16313 24667
rect 16313 24633 16347 24667
rect 16347 24633 16356 24667
rect 16304 24624 16356 24633
rect 17592 24624 17644 24676
rect 18512 24667 18564 24676
rect 18512 24633 18521 24667
rect 18521 24633 18555 24667
rect 18555 24633 18564 24667
rect 18512 24624 18564 24633
rect 18696 24624 18748 24676
rect 15384 24556 15436 24608
rect 15936 24556 15988 24608
rect 16396 24599 16448 24608
rect 16396 24565 16405 24599
rect 16405 24565 16439 24599
rect 16439 24565 16448 24599
rect 16396 24556 16448 24565
rect 16488 24556 16540 24608
rect 17500 24599 17552 24608
rect 17500 24565 17509 24599
rect 17509 24565 17543 24599
rect 17543 24565 17552 24599
rect 17500 24556 17552 24565
rect 17960 24556 18012 24608
rect 20536 24624 20588 24676
rect 21180 24556 21232 24608
rect 21640 24556 21692 24608
rect 21824 24599 21876 24608
rect 21824 24565 21833 24599
rect 21833 24565 21867 24599
rect 21867 24565 21876 24599
rect 21824 24556 21876 24565
rect 22376 24599 22428 24608
rect 22376 24565 22385 24599
rect 22385 24565 22419 24599
rect 22419 24565 22428 24599
rect 22376 24556 22428 24565
rect 23572 24556 23624 24608
rect 24032 24599 24084 24608
rect 24032 24565 24041 24599
rect 24041 24565 24075 24599
rect 24075 24565 24084 24599
rect 24032 24556 24084 24565
rect 24400 24599 24452 24608
rect 24400 24565 24409 24599
rect 24409 24565 24443 24599
rect 24443 24565 24452 24599
rect 24400 24556 24452 24565
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 4988 24352 5040 24404
rect 5264 24352 5316 24404
rect 14832 24352 14884 24404
rect 15752 24352 15804 24404
rect 16488 24395 16540 24404
rect 16488 24361 16497 24395
rect 16497 24361 16531 24395
rect 16531 24361 16540 24395
rect 16488 24352 16540 24361
rect 18788 24352 18840 24404
rect 20628 24395 20680 24404
rect 20628 24361 20637 24395
rect 20637 24361 20671 24395
rect 20671 24361 20680 24395
rect 20628 24352 20680 24361
rect 24124 24352 24176 24404
rect 24676 24395 24728 24404
rect 24676 24361 24685 24395
rect 24685 24361 24719 24395
rect 24719 24361 24728 24395
rect 24676 24352 24728 24361
rect 1124 24284 1176 24336
rect 6184 24327 6236 24336
rect 1860 24216 1912 24268
rect 2228 24216 2280 24268
rect 6184 24293 6193 24327
rect 6193 24293 6227 24327
rect 6227 24293 6236 24327
rect 6184 24284 6236 24293
rect 7104 24284 7156 24336
rect 9404 24284 9456 24336
rect 14188 24284 14240 24336
rect 15384 24284 15436 24336
rect 5540 24216 5592 24268
rect 7196 24216 7248 24268
rect 10140 24216 10192 24268
rect 12992 24216 13044 24268
rect 1952 24148 2004 24200
rect 2136 24191 2188 24200
rect 2136 24157 2145 24191
rect 2145 24157 2179 24191
rect 2179 24157 2188 24191
rect 2136 24148 2188 24157
rect 2964 24148 3016 24200
rect 5080 24148 5132 24200
rect 6644 24191 6696 24200
rect 3884 24080 3936 24132
rect 2228 24012 2280 24064
rect 2504 24012 2556 24064
rect 4068 24012 4120 24064
rect 4344 24055 4396 24064
rect 4344 24021 4353 24055
rect 4353 24021 4387 24055
rect 4387 24021 4396 24055
rect 4344 24012 4396 24021
rect 6644 24157 6653 24191
rect 6653 24157 6687 24191
rect 6687 24157 6696 24191
rect 6644 24148 6696 24157
rect 10416 24191 10468 24200
rect 10416 24157 10425 24191
rect 10425 24157 10459 24191
rect 10459 24157 10468 24191
rect 10416 24148 10468 24157
rect 11428 24148 11480 24200
rect 12164 24148 12216 24200
rect 13360 24191 13412 24200
rect 13360 24157 13369 24191
rect 13369 24157 13403 24191
rect 13403 24157 13412 24191
rect 13360 24148 13412 24157
rect 13452 24191 13504 24200
rect 13452 24157 13461 24191
rect 13461 24157 13495 24191
rect 13495 24157 13504 24191
rect 13452 24148 13504 24157
rect 14096 24148 14148 24200
rect 15108 24148 15160 24200
rect 15292 24148 15344 24200
rect 20996 24284 21048 24336
rect 16672 24216 16724 24268
rect 17684 24216 17736 24268
rect 20444 24216 20496 24268
rect 21272 24259 21324 24268
rect 21272 24225 21281 24259
rect 21281 24225 21315 24259
rect 21315 24225 21324 24259
rect 21272 24216 21324 24225
rect 22652 24216 22704 24268
rect 24124 24216 24176 24268
rect 6368 24080 6420 24132
rect 6552 24080 6604 24132
rect 8208 24080 8260 24132
rect 14004 24080 14056 24132
rect 14832 24080 14884 24132
rect 16948 24148 17000 24200
rect 17408 24148 17460 24200
rect 17868 24148 17920 24200
rect 18604 24191 18656 24200
rect 18604 24157 18613 24191
rect 18613 24157 18647 24191
rect 18647 24157 18656 24191
rect 18604 24148 18656 24157
rect 20720 24148 20772 24200
rect 21364 24191 21416 24200
rect 21364 24157 21373 24191
rect 21373 24157 21407 24191
rect 21407 24157 21416 24191
rect 21364 24148 21416 24157
rect 16672 24080 16724 24132
rect 18420 24080 18472 24132
rect 6092 24012 6144 24064
rect 7564 24012 7616 24064
rect 8668 24055 8720 24064
rect 8668 24021 8677 24055
rect 8677 24021 8711 24055
rect 8711 24021 8720 24055
rect 8668 24012 8720 24021
rect 10140 24012 10192 24064
rect 10324 24055 10376 24064
rect 10324 24021 10333 24055
rect 10333 24021 10367 24055
rect 10367 24021 10376 24055
rect 10324 24012 10376 24021
rect 11796 24055 11848 24064
rect 11796 24021 11805 24055
rect 11805 24021 11839 24055
rect 11839 24021 11848 24055
rect 11796 24012 11848 24021
rect 12072 24012 12124 24064
rect 12900 24055 12952 24064
rect 12900 24021 12909 24055
rect 12909 24021 12943 24055
rect 12943 24021 12952 24055
rect 12900 24012 12952 24021
rect 13728 24012 13780 24064
rect 14464 24055 14516 24064
rect 14464 24021 14473 24055
rect 14473 24021 14507 24055
rect 14507 24021 14516 24055
rect 14464 24012 14516 24021
rect 18052 24012 18104 24064
rect 19248 24012 19300 24064
rect 20352 24012 20404 24064
rect 21548 24012 21600 24064
rect 21824 24012 21876 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 3148 23808 3200 23860
rect 5540 23808 5592 23860
rect 7472 23851 7524 23860
rect 7472 23817 7481 23851
rect 7481 23817 7515 23851
rect 7515 23817 7524 23851
rect 7472 23808 7524 23817
rect 12164 23851 12216 23860
rect 12164 23817 12173 23851
rect 12173 23817 12207 23851
rect 12207 23817 12216 23851
rect 12164 23808 12216 23817
rect 14740 23851 14792 23860
rect 2044 23672 2096 23724
rect 2320 23536 2372 23588
rect 10968 23740 11020 23792
rect 4068 23715 4120 23724
rect 4068 23681 4077 23715
rect 4077 23681 4111 23715
rect 4111 23681 4120 23715
rect 4068 23672 4120 23681
rect 3884 23604 3936 23656
rect 4528 23672 4580 23724
rect 4712 23672 4764 23724
rect 5448 23672 5500 23724
rect 6092 23672 6144 23724
rect 10324 23672 10376 23724
rect 11704 23740 11756 23792
rect 14740 23817 14749 23851
rect 14749 23817 14783 23851
rect 14783 23817 14792 23851
rect 14740 23808 14792 23817
rect 15844 23808 15896 23860
rect 16764 23808 16816 23860
rect 17316 23808 17368 23860
rect 15200 23740 15252 23792
rect 2964 23536 3016 23588
rect 6368 23604 6420 23656
rect 7472 23604 7524 23656
rect 5632 23536 5684 23588
rect 6644 23579 6696 23588
rect 6644 23545 6653 23579
rect 6653 23545 6687 23579
rect 6687 23545 6696 23579
rect 8668 23604 8720 23656
rect 11796 23672 11848 23724
rect 13636 23672 13688 23724
rect 12348 23604 12400 23656
rect 15200 23647 15252 23656
rect 6644 23536 6696 23545
rect 10416 23536 10468 23588
rect 15200 23613 15209 23647
rect 15209 23613 15243 23647
rect 15243 23613 15252 23647
rect 15200 23604 15252 23613
rect 21272 23808 21324 23860
rect 21916 23808 21968 23860
rect 24768 23851 24820 23860
rect 24768 23817 24777 23851
rect 24777 23817 24811 23851
rect 24811 23817 24820 23851
rect 24768 23808 24820 23817
rect 19340 23740 19392 23792
rect 20628 23672 20680 23724
rect 20720 23672 20772 23724
rect 21824 23672 21876 23724
rect 24124 23672 24176 23724
rect 18144 23604 18196 23656
rect 19524 23604 19576 23656
rect 21916 23647 21968 23656
rect 21916 23613 21925 23647
rect 21925 23613 21959 23647
rect 21959 23613 21968 23647
rect 21916 23604 21968 23613
rect 12532 23536 12584 23588
rect 13452 23536 13504 23588
rect 13912 23536 13964 23588
rect 15384 23536 15436 23588
rect 20444 23536 20496 23588
rect 1952 23468 2004 23520
rect 7012 23511 7064 23520
rect 7012 23477 7021 23511
rect 7021 23477 7055 23511
rect 7055 23477 7064 23511
rect 7012 23468 7064 23477
rect 9496 23511 9548 23520
rect 9496 23477 9505 23511
rect 9505 23477 9539 23511
rect 9539 23477 9548 23511
rect 9496 23468 9548 23477
rect 10140 23511 10192 23520
rect 10140 23477 10149 23511
rect 10149 23477 10183 23511
rect 10183 23477 10192 23511
rect 10140 23468 10192 23477
rect 10784 23511 10836 23520
rect 10784 23477 10793 23511
rect 10793 23477 10827 23511
rect 10827 23477 10836 23511
rect 10784 23468 10836 23477
rect 11152 23511 11204 23520
rect 11152 23477 11161 23511
rect 11161 23477 11195 23511
rect 11195 23477 11204 23511
rect 11152 23468 11204 23477
rect 13820 23511 13872 23520
rect 13820 23477 13829 23511
rect 13829 23477 13863 23511
rect 13863 23477 13872 23511
rect 13820 23468 13872 23477
rect 14004 23468 14056 23520
rect 16488 23468 16540 23520
rect 17868 23468 17920 23520
rect 19432 23511 19484 23520
rect 19432 23477 19441 23511
rect 19441 23477 19475 23511
rect 19475 23477 19484 23511
rect 19432 23468 19484 23477
rect 20168 23468 20220 23520
rect 20996 23511 21048 23520
rect 20996 23477 21005 23511
rect 21005 23477 21039 23511
rect 21039 23477 21048 23511
rect 20996 23468 21048 23477
rect 21364 23536 21416 23588
rect 22008 23536 22060 23588
rect 22468 23468 22520 23520
rect 22652 23511 22704 23520
rect 22652 23477 22661 23511
rect 22661 23477 22695 23511
rect 22695 23477 22704 23511
rect 22652 23468 22704 23477
rect 24032 23468 24084 23520
rect 25320 23604 25372 23656
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 1584 23307 1636 23316
rect 1584 23273 1593 23307
rect 1593 23273 1627 23307
rect 1627 23273 1636 23307
rect 1584 23264 1636 23273
rect 3056 23264 3108 23316
rect 5264 23264 5316 23316
rect 7196 23307 7248 23316
rect 7196 23273 7205 23307
rect 7205 23273 7239 23307
rect 7239 23273 7248 23307
rect 7196 23264 7248 23273
rect 3516 23196 3568 23248
rect 2780 23171 2832 23180
rect 2780 23137 2789 23171
rect 2789 23137 2823 23171
rect 2823 23137 2832 23171
rect 2780 23128 2832 23137
rect 3240 23128 3292 23180
rect 5080 23196 5132 23248
rect 9680 23264 9732 23316
rect 5448 23128 5500 23180
rect 5632 23128 5684 23180
rect 6000 23128 6052 23180
rect 3516 23035 3568 23044
rect 3516 23001 3525 23035
rect 3525 23001 3559 23035
rect 3559 23001 3568 23035
rect 3516 22992 3568 23001
rect 8024 23035 8076 23044
rect 8024 23001 8033 23035
rect 8033 23001 8067 23035
rect 8067 23001 8076 23035
rect 8024 22992 8076 23001
rect 8484 23103 8536 23112
rect 8484 23069 8493 23103
rect 8493 23069 8527 23103
rect 8527 23069 8536 23103
rect 8484 23060 8536 23069
rect 9496 23196 9548 23248
rect 9680 23128 9732 23180
rect 9036 22992 9088 23044
rect 10324 23103 10376 23112
rect 10324 23069 10333 23103
rect 10333 23069 10367 23103
rect 10367 23069 10376 23103
rect 10968 23264 11020 23316
rect 12532 23264 12584 23316
rect 13084 23264 13136 23316
rect 13728 23264 13780 23316
rect 13912 23307 13964 23316
rect 13912 23273 13921 23307
rect 13921 23273 13955 23307
rect 13955 23273 13964 23307
rect 13912 23264 13964 23273
rect 14832 23264 14884 23316
rect 15568 23264 15620 23316
rect 12808 23196 12860 23248
rect 16764 23239 16816 23248
rect 16764 23205 16798 23239
rect 16798 23205 16816 23239
rect 16764 23196 16816 23205
rect 20168 23264 20220 23316
rect 20444 23264 20496 23316
rect 21824 23264 21876 23316
rect 22008 23264 22060 23316
rect 22652 23264 22704 23316
rect 22744 23264 22796 23316
rect 24768 23307 24820 23316
rect 24768 23273 24777 23307
rect 24777 23273 24811 23307
rect 24811 23273 24820 23307
rect 24768 23264 24820 23273
rect 19892 23196 19944 23248
rect 20260 23196 20312 23248
rect 22284 23239 22336 23248
rect 22284 23205 22293 23239
rect 22293 23205 22327 23239
rect 22327 23205 22336 23239
rect 22284 23196 22336 23205
rect 11060 23128 11112 23180
rect 11888 23128 11940 23180
rect 12900 23128 12952 23180
rect 14740 23128 14792 23180
rect 16212 23128 16264 23180
rect 19340 23171 19392 23180
rect 19340 23137 19349 23171
rect 19349 23137 19383 23171
rect 19383 23137 19392 23171
rect 21272 23171 21324 23180
rect 19340 23128 19392 23137
rect 21272 23137 21281 23171
rect 21281 23137 21315 23171
rect 21315 23137 21324 23171
rect 21272 23128 21324 23137
rect 21456 23128 21508 23180
rect 22836 23171 22888 23180
rect 11796 23103 11848 23112
rect 10324 23060 10376 23069
rect 11796 23069 11805 23103
rect 11805 23069 11839 23103
rect 11839 23069 11848 23103
rect 11796 23060 11848 23069
rect 13360 23103 13412 23112
rect 13360 23069 13369 23103
rect 13369 23069 13403 23103
rect 13403 23069 13412 23103
rect 13360 23060 13412 23069
rect 13820 23060 13872 23112
rect 15200 23060 15252 23112
rect 16488 23103 16540 23112
rect 16488 23069 16497 23103
rect 16497 23069 16531 23103
rect 16531 23069 16540 23103
rect 16488 23060 16540 23069
rect 20168 23060 20220 23112
rect 20720 23060 20772 23112
rect 22836 23137 22845 23171
rect 22845 23137 22879 23171
rect 22879 23137 22888 23171
rect 22836 23128 22888 23137
rect 24676 23128 24728 23180
rect 23204 23060 23256 23112
rect 12992 22992 13044 23044
rect 13084 22992 13136 23044
rect 13452 22992 13504 23044
rect 17868 23035 17920 23044
rect 17868 23001 17877 23035
rect 17877 23001 17911 23035
rect 17911 23001 17920 23035
rect 17868 22992 17920 23001
rect 1860 22967 1912 22976
rect 1860 22933 1869 22967
rect 1869 22933 1903 22967
rect 1903 22933 1912 22967
rect 1860 22924 1912 22933
rect 4160 22924 4212 22976
rect 6000 22924 6052 22976
rect 6276 22967 6328 22976
rect 6276 22933 6285 22967
rect 6285 22933 6319 22967
rect 6319 22933 6328 22967
rect 6276 22924 6328 22933
rect 6920 22967 6972 22976
rect 6920 22933 6929 22967
rect 6929 22933 6963 22967
rect 6963 22933 6972 22967
rect 6920 22924 6972 22933
rect 9496 22967 9548 22976
rect 9496 22933 9505 22967
rect 9505 22933 9539 22967
rect 9539 22933 9548 22967
rect 9496 22924 9548 22933
rect 12808 22967 12860 22976
rect 12808 22933 12817 22967
rect 12817 22933 12851 22967
rect 12851 22933 12860 22967
rect 12808 22924 12860 22933
rect 18604 22924 18656 22976
rect 18788 22924 18840 22976
rect 18972 22967 19024 22976
rect 18972 22933 18981 22967
rect 18981 22933 19015 22967
rect 19015 22933 19024 22967
rect 18972 22924 19024 22933
rect 20260 22967 20312 22976
rect 20260 22933 20269 22967
rect 20269 22933 20303 22967
rect 20303 22933 20312 22967
rect 20260 22924 20312 22933
rect 20444 22924 20496 22976
rect 22008 22924 22060 22976
rect 22100 22924 22152 22976
rect 23480 22967 23532 22976
rect 23480 22933 23489 22967
rect 23489 22933 23523 22967
rect 23523 22933 23532 22967
rect 23480 22924 23532 22933
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 3884 22720 3936 22772
rect 4988 22720 5040 22772
rect 5356 22720 5408 22772
rect 6828 22763 6880 22772
rect 6828 22729 6837 22763
rect 6837 22729 6871 22763
rect 6871 22729 6880 22763
rect 6828 22720 6880 22729
rect 9404 22720 9456 22772
rect 10324 22720 10376 22772
rect 11060 22763 11112 22772
rect 11060 22729 11069 22763
rect 11069 22729 11103 22763
rect 11103 22729 11112 22763
rect 11060 22720 11112 22729
rect 11428 22763 11480 22772
rect 11428 22729 11437 22763
rect 11437 22729 11471 22763
rect 11471 22729 11480 22763
rect 11428 22720 11480 22729
rect 12440 22763 12492 22772
rect 12440 22729 12449 22763
rect 12449 22729 12483 22763
rect 12483 22729 12492 22763
rect 12440 22720 12492 22729
rect 15384 22720 15436 22772
rect 16212 22763 16264 22772
rect 16212 22729 16221 22763
rect 16221 22729 16255 22763
rect 16255 22729 16264 22763
rect 16212 22720 16264 22729
rect 19524 22763 19576 22772
rect 19524 22729 19533 22763
rect 19533 22729 19567 22763
rect 19567 22729 19576 22763
rect 19524 22720 19576 22729
rect 20076 22720 20128 22772
rect 20996 22763 21048 22772
rect 20996 22729 21005 22763
rect 21005 22729 21039 22763
rect 21039 22729 21048 22763
rect 20996 22720 21048 22729
rect 22836 22763 22888 22772
rect 22836 22729 22845 22763
rect 22845 22729 22879 22763
rect 22879 22729 22888 22763
rect 22836 22720 22888 22729
rect 23848 22763 23900 22772
rect 23848 22729 23857 22763
rect 23857 22729 23891 22763
rect 23891 22729 23900 22763
rect 23848 22720 23900 22729
rect 3056 22652 3108 22704
rect 10140 22652 10192 22704
rect 11796 22652 11848 22704
rect 2780 22584 2832 22636
rect 3148 22627 3200 22636
rect 1492 22380 1544 22432
rect 1584 22380 1636 22432
rect 3148 22593 3157 22627
rect 3157 22593 3191 22627
rect 3191 22593 3200 22627
rect 3148 22584 3200 22593
rect 3332 22627 3384 22636
rect 3332 22593 3341 22627
rect 3341 22593 3375 22627
rect 3375 22593 3384 22627
rect 3332 22584 3384 22593
rect 7564 22584 7616 22636
rect 3424 22516 3476 22568
rect 4528 22559 4580 22568
rect 4528 22525 4562 22559
rect 4562 22525 4580 22559
rect 3148 22448 3200 22500
rect 4528 22516 4580 22525
rect 6276 22516 6328 22568
rect 6920 22516 6972 22568
rect 7196 22559 7248 22568
rect 7196 22525 7205 22559
rect 7205 22525 7239 22559
rect 7239 22525 7248 22559
rect 7196 22516 7248 22525
rect 11060 22584 11112 22636
rect 12900 22627 12952 22636
rect 12900 22593 12909 22627
rect 12909 22593 12943 22627
rect 12943 22593 12952 22627
rect 12900 22584 12952 22593
rect 13360 22652 13412 22704
rect 17040 22695 17092 22704
rect 17040 22661 17049 22695
rect 17049 22661 17083 22695
rect 17083 22661 17092 22695
rect 17040 22652 17092 22661
rect 17592 22652 17644 22704
rect 17868 22695 17920 22704
rect 17868 22661 17877 22695
rect 17877 22661 17911 22695
rect 17911 22661 17920 22695
rect 17868 22652 17920 22661
rect 19616 22695 19668 22704
rect 19616 22661 19625 22695
rect 19625 22661 19659 22695
rect 19659 22661 19668 22695
rect 19616 22652 19668 22661
rect 19892 22652 19944 22704
rect 20720 22695 20772 22704
rect 10048 22516 10100 22568
rect 11244 22559 11296 22568
rect 11244 22525 11253 22559
rect 11253 22525 11287 22559
rect 11287 22525 11296 22559
rect 11244 22516 11296 22525
rect 11980 22516 12032 22568
rect 12716 22516 12768 22568
rect 13360 22516 13412 22568
rect 13544 22516 13596 22568
rect 4712 22448 4764 22500
rect 7012 22448 7064 22500
rect 7380 22448 7432 22500
rect 7932 22448 7984 22500
rect 8944 22491 8996 22500
rect 8944 22457 8978 22491
rect 8978 22457 8996 22491
rect 8944 22448 8996 22457
rect 9956 22448 10008 22500
rect 10784 22448 10836 22500
rect 18052 22584 18104 22636
rect 18512 22627 18564 22636
rect 18512 22593 18521 22627
rect 18521 22593 18555 22627
rect 18555 22593 18564 22627
rect 18512 22584 18564 22593
rect 18696 22627 18748 22636
rect 18696 22593 18705 22627
rect 18705 22593 18739 22627
rect 18739 22593 18748 22627
rect 18696 22584 18748 22593
rect 19432 22584 19484 22636
rect 20444 22584 20496 22636
rect 3332 22380 3384 22432
rect 3792 22380 3844 22432
rect 5264 22380 5316 22432
rect 5632 22423 5684 22432
rect 5632 22389 5641 22423
rect 5641 22389 5675 22423
rect 5675 22389 5684 22423
rect 5632 22380 5684 22389
rect 6276 22380 6328 22432
rect 6552 22380 6604 22432
rect 10048 22423 10100 22432
rect 10048 22389 10057 22423
rect 10057 22389 10091 22423
rect 10091 22389 10100 22423
rect 10048 22380 10100 22389
rect 11888 22423 11940 22432
rect 11888 22389 11897 22423
rect 11897 22389 11931 22423
rect 11931 22389 11940 22423
rect 11888 22380 11940 22389
rect 13452 22423 13504 22432
rect 13452 22389 13461 22423
rect 13461 22389 13495 22423
rect 13495 22389 13504 22423
rect 13452 22380 13504 22389
rect 13544 22380 13596 22432
rect 13728 22380 13780 22432
rect 14188 22423 14240 22432
rect 14188 22389 14197 22423
rect 14197 22389 14231 22423
rect 14231 22389 14240 22423
rect 16304 22516 16356 22568
rect 17868 22516 17920 22568
rect 18972 22516 19024 22568
rect 19248 22516 19300 22568
rect 19800 22516 19852 22568
rect 20076 22559 20128 22568
rect 20076 22525 20085 22559
rect 20085 22525 20119 22559
rect 20119 22525 20128 22559
rect 20076 22516 20128 22525
rect 20720 22661 20729 22695
rect 20729 22661 20763 22695
rect 20763 22661 20772 22695
rect 20720 22652 20772 22661
rect 22744 22652 22796 22704
rect 21456 22584 21508 22636
rect 20720 22516 20772 22568
rect 20996 22516 21048 22568
rect 14648 22448 14700 22500
rect 16488 22448 16540 22500
rect 18144 22448 18196 22500
rect 21824 22516 21876 22568
rect 23664 22559 23716 22568
rect 23664 22525 23673 22559
rect 23673 22525 23707 22559
rect 23707 22525 23716 22559
rect 23664 22516 23716 22525
rect 24676 22491 24728 22500
rect 24676 22457 24685 22491
rect 24685 22457 24719 22491
rect 24719 22457 24728 22491
rect 24676 22448 24728 22457
rect 14188 22380 14240 22389
rect 15292 22380 15344 22432
rect 18052 22423 18104 22432
rect 18052 22389 18061 22423
rect 18061 22389 18095 22423
rect 18095 22389 18104 22423
rect 18052 22380 18104 22389
rect 18236 22380 18288 22432
rect 20996 22380 21048 22432
rect 21364 22380 21416 22432
rect 23204 22423 23256 22432
rect 23204 22389 23213 22423
rect 23213 22389 23247 22423
rect 23247 22389 23256 22423
rect 23204 22380 23256 22389
rect 24768 22423 24820 22432
rect 24768 22389 24777 22423
rect 24777 22389 24811 22423
rect 24811 22389 24820 22423
rect 24768 22380 24820 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 1860 22176 1912 22228
rect 1032 22040 1084 22092
rect 1492 22040 1544 22092
rect 1124 21972 1176 22024
rect 4068 22176 4120 22228
rect 4344 22176 4396 22228
rect 5448 22219 5500 22228
rect 5448 22185 5457 22219
rect 5457 22185 5491 22219
rect 5491 22185 5500 22219
rect 5448 22176 5500 22185
rect 6184 22176 6236 22228
rect 8208 22176 8260 22228
rect 9864 22219 9916 22228
rect 9864 22185 9873 22219
rect 9873 22185 9907 22219
rect 9907 22185 9916 22219
rect 9864 22176 9916 22185
rect 10692 22176 10744 22228
rect 13544 22219 13596 22228
rect 13544 22185 13553 22219
rect 13553 22185 13587 22219
rect 13587 22185 13596 22219
rect 13544 22176 13596 22185
rect 2964 22108 3016 22160
rect 3240 22040 3292 22092
rect 2780 21972 2832 22024
rect 1952 21904 2004 21956
rect 4712 22108 4764 22160
rect 5632 22108 5684 22160
rect 8392 22151 8444 22160
rect 4528 22040 4580 22092
rect 6368 22083 6420 22092
rect 6368 22049 6377 22083
rect 6377 22049 6411 22083
rect 6411 22049 6420 22083
rect 6368 22040 6420 22049
rect 3608 21972 3660 22024
rect 4160 21972 4212 22024
rect 4896 22015 4948 22024
rect 4896 21981 4905 22015
rect 4905 21981 4939 22015
rect 4939 21981 4948 22015
rect 4896 21972 4948 21981
rect 4988 22015 5040 22024
rect 4988 21981 4997 22015
rect 4997 21981 5031 22015
rect 5031 21981 5040 22015
rect 8392 22117 8401 22151
rect 8401 22117 8435 22151
rect 8435 22117 8444 22151
rect 8392 22108 8444 22117
rect 10048 22108 10100 22160
rect 9404 22083 9456 22092
rect 9404 22049 9413 22083
rect 9413 22049 9447 22083
rect 9447 22049 9456 22083
rect 9404 22040 9456 22049
rect 9680 22083 9732 22092
rect 9680 22049 9689 22083
rect 9689 22049 9723 22083
rect 9723 22049 9732 22083
rect 9680 22040 9732 22049
rect 12716 22108 12768 22160
rect 13912 22151 13964 22160
rect 13912 22117 13921 22151
rect 13921 22117 13955 22151
rect 13955 22117 13964 22151
rect 13912 22108 13964 22117
rect 11336 22083 11388 22092
rect 11336 22049 11370 22083
rect 11370 22049 11388 22083
rect 11336 22040 11388 22049
rect 16120 22176 16172 22228
rect 16304 22176 16356 22228
rect 16764 22176 16816 22228
rect 16948 22176 17000 22228
rect 17776 22176 17828 22228
rect 20076 22176 20128 22228
rect 20260 22219 20312 22228
rect 20260 22185 20269 22219
rect 20269 22185 20303 22219
rect 20303 22185 20312 22219
rect 20260 22176 20312 22185
rect 21272 22176 21324 22228
rect 16488 22108 16540 22160
rect 18696 22108 18748 22160
rect 20352 22108 20404 22160
rect 15292 22083 15344 22092
rect 15292 22049 15301 22083
rect 15301 22049 15335 22083
rect 15335 22049 15344 22083
rect 15292 22040 15344 22049
rect 15844 22040 15896 22092
rect 15936 22040 15988 22092
rect 4988 21972 5040 21981
rect 6644 21972 6696 22024
rect 6736 21972 6788 22024
rect 7104 22015 7156 22024
rect 7104 21981 7113 22015
rect 7113 21981 7147 22015
rect 7147 21981 7156 22015
rect 7104 21972 7156 21981
rect 8484 22015 8536 22024
rect 8484 21981 8493 22015
rect 8493 21981 8527 22015
rect 8527 21981 8536 22015
rect 8484 21972 8536 21981
rect 6460 21947 6512 21956
rect 6460 21913 6469 21947
rect 6469 21913 6503 21947
rect 6503 21913 6512 21947
rect 6460 21904 6512 21913
rect 8300 21904 8352 21956
rect 9588 21972 9640 22024
rect 11060 22015 11112 22024
rect 11060 21981 11069 22015
rect 11069 21981 11103 22015
rect 11103 21981 11112 22015
rect 11060 21972 11112 21981
rect 14004 22015 14056 22024
rect 14004 21981 14013 22015
rect 14013 21981 14047 22015
rect 14047 21981 14056 22015
rect 14004 21972 14056 21981
rect 12532 21904 12584 21956
rect 12808 21904 12860 21956
rect 16948 22040 17000 22092
rect 17500 22040 17552 22092
rect 17868 22040 17920 22092
rect 18512 22040 18564 22092
rect 18880 22040 18932 22092
rect 19708 22083 19760 22092
rect 17132 21972 17184 22024
rect 18604 22015 18656 22024
rect 18604 21981 18613 22015
rect 18613 21981 18647 22015
rect 18647 21981 18656 22015
rect 18604 21972 18656 21981
rect 18696 22015 18748 22024
rect 18696 21981 18705 22015
rect 18705 21981 18739 22015
rect 18739 21981 18748 22015
rect 18696 21972 18748 21981
rect 19156 21972 19208 22024
rect 19708 22049 19717 22083
rect 19717 22049 19751 22083
rect 19751 22049 19760 22083
rect 19708 22040 19760 22049
rect 20168 22040 20220 22092
rect 20720 22040 20772 22092
rect 20260 21972 20312 22024
rect 20352 21972 20404 22024
rect 22008 22176 22060 22228
rect 22468 22219 22520 22228
rect 22468 22185 22477 22219
rect 22477 22185 22511 22219
rect 22511 22185 22520 22219
rect 22468 22176 22520 22185
rect 23020 22219 23072 22228
rect 23020 22185 23029 22219
rect 23029 22185 23063 22219
rect 23063 22185 23072 22219
rect 23020 22176 23072 22185
rect 22836 22040 22888 22092
rect 24032 22040 24084 22092
rect 24860 22040 24912 22092
rect 25228 22040 25280 22092
rect 21732 22015 21784 22024
rect 21732 21981 21741 22015
rect 21741 21981 21775 22015
rect 21775 21981 21784 22015
rect 21732 21972 21784 21981
rect 22744 21972 22796 22024
rect 23296 22015 23348 22024
rect 23296 21981 23305 22015
rect 23305 21981 23339 22015
rect 23339 21981 23348 22015
rect 23296 21972 23348 21981
rect 16488 21904 16540 21956
rect 17500 21904 17552 21956
rect 17684 21904 17736 21956
rect 19800 21904 19852 21956
rect 20076 21904 20128 21956
rect 24124 21972 24176 22024
rect 24216 21972 24268 22024
rect 23940 21904 23992 21956
rect 3240 21836 3292 21888
rect 3516 21879 3568 21888
rect 3516 21845 3525 21879
rect 3525 21845 3559 21879
rect 3559 21845 3568 21879
rect 3516 21836 3568 21845
rect 3792 21879 3844 21888
rect 3792 21845 3801 21879
rect 3801 21845 3835 21879
rect 3835 21845 3844 21879
rect 3792 21836 3844 21845
rect 6092 21836 6144 21888
rect 6368 21836 6420 21888
rect 7288 21836 7340 21888
rect 7564 21836 7616 21888
rect 10140 21836 10192 21888
rect 13268 21836 13320 21888
rect 14188 21836 14240 21888
rect 14648 21879 14700 21888
rect 14648 21845 14657 21879
rect 14657 21845 14691 21879
rect 14691 21845 14700 21879
rect 14648 21836 14700 21845
rect 19248 21879 19300 21888
rect 19248 21845 19257 21879
rect 19257 21845 19291 21879
rect 19291 21845 19300 21879
rect 19248 21836 19300 21845
rect 19892 21879 19944 21888
rect 19892 21845 19901 21879
rect 19901 21845 19935 21879
rect 19935 21845 19944 21879
rect 19892 21836 19944 21845
rect 20536 21836 20588 21888
rect 20720 21879 20772 21888
rect 20720 21845 20729 21879
rect 20729 21845 20763 21879
rect 20763 21845 20772 21879
rect 20720 21836 20772 21845
rect 22008 21836 22060 21888
rect 23756 21879 23808 21888
rect 23756 21845 23765 21879
rect 23765 21845 23799 21879
rect 23799 21845 23808 21879
rect 23756 21836 23808 21845
rect 24032 21879 24084 21888
rect 24032 21845 24041 21879
rect 24041 21845 24075 21879
rect 24075 21845 24084 21879
rect 24032 21836 24084 21845
rect 24124 21836 24176 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1308 21632 1360 21684
rect 1860 21675 1912 21684
rect 1860 21641 1869 21675
rect 1869 21641 1903 21675
rect 1903 21641 1912 21675
rect 1860 21632 1912 21641
rect 4896 21632 4948 21684
rect 5080 21632 5132 21684
rect 3424 21607 3476 21616
rect 2780 21496 2832 21548
rect 664 21428 716 21480
rect 3424 21573 3433 21607
rect 3433 21573 3467 21607
rect 3467 21573 3476 21607
rect 3424 21564 3476 21573
rect 3884 21564 3936 21616
rect 6828 21564 6880 21616
rect 8944 21632 8996 21684
rect 11060 21632 11112 21684
rect 11336 21632 11388 21684
rect 11888 21632 11940 21684
rect 12624 21632 12676 21684
rect 12808 21675 12860 21684
rect 12808 21641 12817 21675
rect 12817 21641 12851 21675
rect 12851 21641 12860 21675
rect 12808 21632 12860 21641
rect 9220 21564 9272 21616
rect 9680 21564 9732 21616
rect 14004 21632 14056 21684
rect 15292 21675 15344 21684
rect 15292 21641 15301 21675
rect 15301 21641 15335 21675
rect 15335 21641 15344 21675
rect 15292 21632 15344 21641
rect 16764 21632 16816 21684
rect 17040 21632 17092 21684
rect 18052 21632 18104 21684
rect 18604 21632 18656 21684
rect 19708 21632 19760 21684
rect 21088 21675 21140 21684
rect 21088 21641 21097 21675
rect 21097 21641 21131 21675
rect 21131 21641 21140 21675
rect 21088 21632 21140 21641
rect 23020 21675 23072 21684
rect 23020 21641 23029 21675
rect 23029 21641 23063 21675
rect 23063 21641 23072 21675
rect 23020 21632 23072 21641
rect 24860 21632 24912 21684
rect 25412 21675 25464 21684
rect 25412 21641 25421 21675
rect 25421 21641 25455 21675
rect 25455 21641 25464 21675
rect 25412 21632 25464 21641
rect 21456 21564 21508 21616
rect 23296 21564 23348 21616
rect 23756 21564 23808 21616
rect 3516 21496 3568 21548
rect 5540 21539 5592 21548
rect 5540 21505 5549 21539
rect 5549 21505 5583 21539
rect 5583 21505 5592 21539
rect 5540 21496 5592 21505
rect 9864 21496 9916 21548
rect 13268 21539 13320 21548
rect 13268 21505 13277 21539
rect 13277 21505 13311 21539
rect 13311 21505 13320 21539
rect 13268 21496 13320 21505
rect 17592 21496 17644 21548
rect 18144 21496 18196 21548
rect 18604 21539 18656 21548
rect 18604 21505 18613 21539
rect 18613 21505 18647 21539
rect 18647 21505 18656 21539
rect 18604 21496 18656 21505
rect 19800 21496 19852 21548
rect 20444 21496 20496 21548
rect 20904 21496 20956 21548
rect 22376 21496 22428 21548
rect 24032 21496 24084 21548
rect 24400 21496 24452 21548
rect 7104 21428 7156 21480
rect 7564 21428 7616 21480
rect 9680 21428 9732 21480
rect 11152 21428 11204 21480
rect 6184 21360 6236 21412
rect 8300 21360 8352 21412
rect 10692 21360 10744 21412
rect 11796 21360 11848 21412
rect 16396 21428 16448 21480
rect 18696 21428 18748 21480
rect 21180 21428 21232 21480
rect 23020 21428 23072 21480
rect 14004 21360 14056 21412
rect 14464 21360 14516 21412
rect 2044 21292 2096 21344
rect 2596 21292 2648 21344
rect 3516 21292 3568 21344
rect 5448 21335 5500 21344
rect 5448 21301 5457 21335
rect 5457 21301 5491 21335
rect 5491 21301 5500 21335
rect 5448 21292 5500 21301
rect 6736 21292 6788 21344
rect 8392 21292 8444 21344
rect 10140 21292 10192 21344
rect 10876 21292 10928 21344
rect 16672 21360 16724 21412
rect 18512 21360 18564 21412
rect 21088 21360 21140 21412
rect 21916 21360 21968 21412
rect 23940 21360 23992 21412
rect 14740 21292 14792 21344
rect 15844 21292 15896 21344
rect 16396 21335 16448 21344
rect 16396 21301 16405 21335
rect 16405 21301 16439 21335
rect 16439 21301 16448 21335
rect 16396 21292 16448 21301
rect 17040 21292 17092 21344
rect 17868 21292 17920 21344
rect 18604 21292 18656 21344
rect 18696 21292 18748 21344
rect 19340 21292 19392 21344
rect 20628 21292 20680 21344
rect 21732 21292 21784 21344
rect 22468 21292 22520 21344
rect 22744 21335 22796 21344
rect 22744 21301 22753 21335
rect 22753 21301 22787 21335
rect 22787 21301 22796 21335
rect 22744 21292 22796 21301
rect 23756 21292 23808 21344
rect 24584 21292 24636 21344
rect 25780 21335 25832 21344
rect 25780 21301 25789 21335
rect 25789 21301 25823 21335
rect 25823 21301 25832 21335
rect 25780 21292 25832 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1124 21088 1176 21140
rect 2320 21088 2372 21140
rect 3148 21088 3200 21140
rect 4068 21131 4120 21140
rect 4068 21097 4077 21131
rect 4077 21097 4111 21131
rect 4111 21097 4120 21131
rect 4068 21088 4120 21097
rect 5448 21131 5500 21140
rect 5448 21097 5457 21131
rect 5457 21097 5491 21131
rect 5491 21097 5500 21131
rect 5448 21088 5500 21097
rect 7104 21131 7156 21140
rect 7104 21097 7113 21131
rect 7113 21097 7147 21131
rect 7147 21097 7156 21131
rect 7104 21088 7156 21097
rect 8300 21131 8352 21140
rect 8300 21097 8309 21131
rect 8309 21097 8343 21131
rect 8343 21097 8352 21131
rect 9036 21131 9088 21140
rect 8300 21088 8352 21097
rect 3332 21020 3384 21072
rect 6092 21020 6144 21072
rect 8208 21020 8260 21072
rect 9036 21097 9045 21131
rect 9045 21097 9079 21131
rect 9079 21097 9088 21131
rect 9036 21088 9088 21097
rect 11796 21131 11848 21140
rect 11796 21097 11805 21131
rect 11805 21097 11839 21131
rect 11839 21097 11848 21131
rect 11796 21088 11848 21097
rect 12256 21131 12308 21140
rect 12256 21097 12265 21131
rect 12265 21097 12299 21131
rect 12299 21097 12308 21131
rect 12256 21088 12308 21097
rect 13636 21131 13688 21140
rect 13636 21097 13645 21131
rect 13645 21097 13679 21131
rect 13679 21097 13688 21131
rect 13636 21088 13688 21097
rect 14280 21131 14332 21140
rect 14280 21097 14289 21131
rect 14289 21097 14323 21131
rect 14323 21097 14332 21131
rect 14280 21088 14332 21097
rect 14556 21088 14608 21140
rect 15752 21131 15804 21140
rect 15752 21097 15761 21131
rect 15761 21097 15795 21131
rect 15795 21097 15804 21131
rect 15752 21088 15804 21097
rect 17408 21088 17460 21140
rect 20352 21131 20404 21140
rect 20352 21097 20361 21131
rect 20361 21097 20395 21131
rect 20395 21097 20404 21131
rect 20352 21088 20404 21097
rect 20904 21088 20956 21140
rect 21180 21131 21232 21140
rect 21180 21097 21189 21131
rect 21189 21097 21223 21131
rect 21223 21097 21232 21131
rect 21180 21088 21232 21097
rect 24768 21088 24820 21140
rect 1492 20952 1544 21004
rect 2780 20952 2832 21004
rect 4160 20952 4212 21004
rect 6000 20995 6052 21004
rect 5448 20884 5500 20936
rect 2872 20816 2924 20868
rect 3148 20816 3200 20868
rect 6000 20961 6009 20995
rect 6009 20961 6043 20995
rect 6043 20961 6052 20995
rect 6000 20952 6052 20961
rect 7932 20952 7984 21004
rect 9680 20952 9732 21004
rect 9864 20952 9916 21004
rect 6092 20927 6144 20936
rect 6092 20893 6101 20927
rect 6101 20893 6135 20927
rect 6135 20893 6144 20927
rect 6092 20884 6144 20893
rect 6460 20884 6512 20936
rect 11428 21020 11480 21072
rect 13452 21020 13504 21072
rect 15108 21063 15160 21072
rect 15108 21029 15117 21063
rect 15117 21029 15151 21063
rect 15151 21029 15160 21063
rect 15108 21020 15160 21029
rect 16948 21020 17000 21072
rect 18144 21063 18196 21072
rect 18144 21029 18153 21063
rect 18153 21029 18187 21063
rect 18187 21029 18196 21063
rect 18144 21020 18196 21029
rect 18696 21020 18748 21072
rect 20812 21020 20864 21072
rect 21548 21063 21600 21072
rect 21548 21029 21557 21063
rect 21557 21029 21591 21063
rect 21591 21029 21600 21063
rect 21548 21020 21600 21029
rect 22928 21020 22980 21072
rect 24676 21063 24728 21072
rect 24676 21029 24685 21063
rect 24685 21029 24719 21063
rect 24719 21029 24728 21063
rect 24676 21020 24728 21029
rect 12624 20995 12676 21004
rect 12624 20961 12633 20995
rect 12633 20961 12667 20995
rect 12667 20961 12676 20995
rect 12624 20952 12676 20961
rect 12716 20995 12768 21004
rect 12716 20961 12725 20995
rect 12725 20961 12759 20995
rect 12759 20961 12768 20995
rect 12716 20952 12768 20961
rect 14280 20952 14332 21004
rect 15292 20952 15344 21004
rect 12900 20927 12952 20936
rect 7288 20816 7340 20868
rect 8484 20816 8536 20868
rect 9588 20816 9640 20868
rect 12900 20893 12909 20927
rect 12909 20893 12943 20927
rect 12943 20893 12952 20927
rect 12900 20884 12952 20893
rect 15844 20927 15896 20936
rect 15844 20893 15853 20927
rect 15853 20893 15887 20927
rect 15887 20893 15896 20927
rect 15844 20884 15896 20893
rect 17868 20884 17920 20936
rect 18512 20952 18564 21004
rect 19984 20952 20036 21004
rect 21456 20952 21508 21004
rect 23940 20952 23992 21004
rect 19156 20884 19208 20936
rect 12072 20816 12124 20868
rect 12256 20816 12308 20868
rect 14464 20816 14516 20868
rect 17776 20816 17828 20868
rect 18512 20816 18564 20868
rect 19248 20816 19300 20868
rect 20260 20884 20312 20936
rect 20628 20884 20680 20936
rect 20904 20884 20956 20936
rect 24400 20816 24452 20868
rect 3516 20791 3568 20800
rect 3516 20757 3525 20791
rect 3525 20757 3559 20791
rect 3559 20757 3568 20791
rect 3516 20748 3568 20757
rect 4988 20748 5040 20800
rect 6736 20791 6788 20800
rect 6736 20757 6745 20791
rect 6745 20757 6779 20791
rect 6779 20757 6788 20791
rect 6736 20748 6788 20757
rect 6920 20748 6972 20800
rect 9404 20791 9456 20800
rect 9404 20757 9413 20791
rect 9413 20757 9447 20791
rect 9447 20757 9456 20791
rect 9404 20748 9456 20757
rect 14004 20791 14056 20800
rect 14004 20757 14013 20791
rect 14013 20757 14047 20791
rect 14047 20757 14056 20791
rect 14004 20748 14056 20757
rect 21364 20748 21416 20800
rect 21916 20748 21968 20800
rect 22468 20748 22520 20800
rect 23664 20791 23716 20800
rect 23664 20757 23673 20791
rect 23673 20757 23707 20791
rect 23707 20757 23716 20791
rect 23664 20748 23716 20757
rect 24032 20791 24084 20800
rect 24032 20757 24041 20791
rect 24041 20757 24075 20791
rect 24075 20757 24084 20791
rect 24032 20748 24084 20757
rect 24124 20748 24176 20800
rect 24768 20748 24820 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1216 20544 1268 20596
rect 2136 20544 2188 20596
rect 3148 20544 3200 20596
rect 6000 20544 6052 20596
rect 6460 20544 6512 20596
rect 2872 20476 2924 20528
rect 3700 20476 3752 20528
rect 2412 20451 2464 20460
rect 2412 20417 2421 20451
rect 2421 20417 2455 20451
rect 2455 20417 2464 20451
rect 2412 20408 2464 20417
rect 2504 20408 2556 20460
rect 2780 20408 2832 20460
rect 5264 20408 5316 20460
rect 6000 20408 6052 20460
rect 6828 20544 6880 20596
rect 9588 20544 9640 20596
rect 12624 20544 12676 20596
rect 12900 20544 12952 20596
rect 14096 20544 14148 20596
rect 15752 20587 15804 20596
rect 15752 20553 15761 20587
rect 15761 20553 15795 20587
rect 15795 20553 15804 20587
rect 15752 20544 15804 20553
rect 17868 20544 17920 20596
rect 18512 20587 18564 20596
rect 18512 20553 18521 20587
rect 18521 20553 18555 20587
rect 18555 20553 18564 20587
rect 18512 20544 18564 20553
rect 21456 20544 21508 20596
rect 22192 20544 22244 20596
rect 22652 20544 22704 20596
rect 22928 20544 22980 20596
rect 16396 20519 16448 20528
rect 16396 20485 16405 20519
rect 16405 20485 16439 20519
rect 16439 20485 16448 20519
rect 16396 20476 16448 20485
rect 7104 20408 7156 20460
rect 9864 20408 9916 20460
rect 14464 20451 14516 20460
rect 14464 20417 14473 20451
rect 14473 20417 14507 20451
rect 14507 20417 14516 20451
rect 14464 20408 14516 20417
rect 14648 20451 14700 20460
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 16948 20451 17000 20460
rect 16948 20417 16957 20451
rect 16957 20417 16991 20451
rect 16991 20417 17000 20451
rect 16948 20408 17000 20417
rect 18604 20408 18656 20460
rect 21548 20408 21600 20460
rect 22376 20408 22428 20460
rect 3332 20340 3384 20392
rect 4712 20340 4764 20392
rect 5816 20383 5868 20392
rect 5816 20349 5825 20383
rect 5825 20349 5859 20383
rect 5859 20349 5868 20383
rect 5816 20340 5868 20349
rect 6092 20340 6144 20392
rect 3516 20272 3568 20324
rect 4988 20272 5040 20324
rect 7564 20272 7616 20324
rect 7840 20340 7892 20392
rect 9680 20383 9732 20392
rect 9680 20349 9689 20383
rect 9689 20349 9723 20383
rect 9723 20349 9732 20383
rect 9680 20340 9732 20349
rect 11612 20340 11664 20392
rect 10784 20272 10836 20324
rect 13820 20340 13872 20392
rect 19340 20383 19392 20392
rect 19340 20349 19374 20383
rect 19374 20349 19392 20383
rect 19340 20340 19392 20349
rect 23020 20340 23072 20392
rect 25964 20383 26016 20392
rect 25964 20349 25973 20383
rect 25973 20349 26007 20383
rect 26007 20349 26016 20383
rect 25964 20340 26016 20349
rect 11980 20272 12032 20324
rect 13728 20272 13780 20324
rect 14740 20272 14792 20324
rect 16488 20272 16540 20324
rect 20720 20272 20772 20324
rect 2320 20247 2372 20256
rect 2320 20213 2329 20247
rect 2329 20213 2363 20247
rect 2363 20213 2372 20247
rect 2320 20204 2372 20213
rect 4344 20204 4396 20256
rect 5264 20247 5316 20256
rect 5264 20213 5273 20247
rect 5273 20213 5307 20247
rect 5307 20213 5316 20247
rect 5264 20204 5316 20213
rect 7196 20247 7248 20256
rect 7196 20213 7205 20247
rect 7205 20213 7239 20247
rect 7239 20213 7248 20247
rect 7196 20204 7248 20213
rect 8760 20204 8812 20256
rect 10048 20247 10100 20256
rect 10048 20213 10057 20247
rect 10057 20213 10091 20247
rect 10091 20213 10100 20247
rect 10048 20204 10100 20213
rect 12900 20247 12952 20256
rect 12900 20213 12909 20247
rect 12909 20213 12943 20247
rect 12943 20213 12952 20247
rect 12900 20204 12952 20213
rect 14280 20204 14332 20256
rect 16212 20247 16264 20256
rect 16212 20213 16221 20247
rect 16221 20213 16255 20247
rect 16255 20213 16264 20247
rect 16212 20204 16264 20213
rect 17316 20204 17368 20256
rect 18328 20204 18380 20256
rect 19340 20204 19392 20256
rect 20444 20247 20496 20256
rect 20444 20213 20453 20247
rect 20453 20213 20487 20247
rect 20487 20213 20496 20247
rect 20444 20204 20496 20213
rect 21548 20247 21600 20256
rect 21548 20213 21557 20247
rect 21557 20213 21591 20247
rect 21591 20213 21600 20247
rect 21548 20204 21600 20213
rect 23664 20204 23716 20256
rect 24032 20204 24084 20256
rect 25780 20204 25832 20256
rect 25964 20204 26016 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 940 20000 992 20052
rect 2320 20000 2372 20052
rect 4988 20000 5040 20052
rect 7196 20000 7248 20052
rect 7840 20043 7892 20052
rect 7840 20009 7849 20043
rect 7849 20009 7883 20043
rect 7883 20009 7892 20043
rect 7840 20000 7892 20009
rect 8300 20043 8352 20052
rect 8300 20009 8309 20043
rect 8309 20009 8343 20043
rect 8343 20009 8352 20043
rect 8300 20000 8352 20009
rect 9680 20043 9732 20052
rect 9680 20009 9689 20043
rect 9689 20009 9723 20043
rect 9723 20009 9732 20043
rect 9680 20000 9732 20009
rect 10140 20000 10192 20052
rect 10784 20000 10836 20052
rect 11060 20000 11112 20052
rect 11520 20000 11572 20052
rect 12900 20000 12952 20052
rect 15108 20043 15160 20052
rect 15108 20009 15117 20043
rect 15117 20009 15151 20043
rect 15151 20009 15160 20043
rect 15108 20000 15160 20009
rect 15660 20000 15712 20052
rect 16488 20043 16540 20052
rect 16488 20009 16497 20043
rect 16497 20009 16531 20043
rect 16531 20009 16540 20043
rect 16488 20000 16540 20009
rect 16856 20000 16908 20052
rect 17408 20043 17460 20052
rect 17408 20009 17417 20043
rect 17417 20009 17451 20043
rect 17451 20009 17460 20043
rect 17408 20000 17460 20009
rect 18144 20043 18196 20052
rect 18144 20009 18153 20043
rect 18153 20009 18187 20043
rect 18187 20009 18196 20043
rect 18144 20000 18196 20009
rect 18972 20000 19024 20052
rect 2872 19975 2924 19984
rect 2872 19941 2881 19975
rect 2881 19941 2915 19975
rect 2915 19941 2924 19975
rect 2872 19932 2924 19941
rect 3516 19975 3568 19984
rect 3516 19941 3525 19975
rect 3525 19941 3559 19975
rect 3559 19941 3568 19975
rect 3516 19932 3568 19941
rect 3792 19864 3844 19916
rect 3056 19839 3108 19848
rect 3056 19805 3065 19839
rect 3065 19805 3099 19839
rect 3099 19805 3108 19839
rect 3056 19796 3108 19805
rect 4160 19932 4212 19984
rect 17132 19932 17184 19984
rect 17776 19932 17828 19984
rect 19432 20000 19484 20052
rect 22100 20000 22152 20052
rect 24676 20000 24728 20052
rect 24860 20043 24912 20052
rect 24860 20009 24869 20043
rect 24869 20009 24903 20043
rect 24903 20009 24912 20043
rect 24860 20000 24912 20009
rect 25136 20043 25188 20052
rect 25136 20009 25145 20043
rect 25145 20009 25179 20043
rect 25179 20009 25188 20043
rect 25136 20000 25188 20009
rect 19248 19932 19300 19984
rect 21272 19932 21324 19984
rect 23112 19932 23164 19984
rect 24584 19932 24636 19984
rect 4068 19907 4120 19916
rect 4068 19873 4077 19907
rect 4077 19873 4111 19907
rect 4111 19873 4120 19907
rect 4068 19864 4120 19873
rect 4712 19907 4764 19916
rect 4712 19873 4721 19907
rect 4721 19873 4755 19907
rect 4755 19873 4764 19907
rect 4712 19864 4764 19873
rect 4988 19864 5040 19916
rect 5540 19864 5592 19916
rect 6736 19864 6788 19916
rect 8024 19864 8076 19916
rect 11888 19864 11940 19916
rect 12808 19864 12860 19916
rect 16488 19864 16540 19916
rect 16948 19864 17000 19916
rect 8760 19796 8812 19848
rect 11244 19839 11296 19848
rect 11244 19805 11253 19839
rect 11253 19805 11287 19839
rect 11287 19805 11296 19839
rect 11244 19796 11296 19805
rect 11704 19839 11756 19848
rect 11704 19805 11713 19839
rect 11713 19805 11747 19839
rect 11747 19805 11756 19839
rect 11704 19796 11756 19805
rect 12716 19839 12768 19848
rect 12716 19805 12725 19839
rect 12725 19805 12759 19839
rect 12759 19805 12768 19839
rect 12716 19796 12768 19805
rect 15752 19796 15804 19848
rect 18512 19864 18564 19916
rect 20904 19839 20956 19848
rect 4160 19728 4212 19780
rect 5448 19728 5500 19780
rect 7932 19771 7984 19780
rect 7932 19737 7941 19771
rect 7941 19737 7975 19771
rect 7975 19737 7984 19771
rect 7932 19728 7984 19737
rect 9588 19728 9640 19780
rect 10784 19728 10836 19780
rect 11152 19728 11204 19780
rect 13820 19728 13872 19780
rect 14280 19728 14332 19780
rect 17040 19771 17092 19780
rect 17040 19737 17049 19771
rect 17049 19737 17083 19771
rect 17083 19737 17092 19771
rect 17040 19728 17092 19737
rect 19340 19728 19392 19780
rect 1492 19660 1544 19712
rect 4252 19703 4304 19712
rect 4252 19669 4261 19703
rect 4261 19669 4295 19703
rect 4295 19669 4304 19703
rect 4252 19660 4304 19669
rect 4344 19660 4396 19712
rect 4712 19660 4764 19712
rect 7472 19660 7524 19712
rect 9496 19703 9548 19712
rect 9496 19669 9505 19703
rect 9505 19669 9539 19703
rect 9539 19669 9548 19703
rect 9496 19660 9548 19669
rect 9864 19660 9916 19712
rect 14004 19660 14056 19712
rect 14556 19660 14608 19712
rect 15384 19660 15436 19712
rect 16948 19703 17000 19712
rect 16948 19669 16957 19703
rect 16957 19669 16991 19703
rect 16991 19669 17000 19703
rect 16948 19660 17000 19669
rect 18604 19703 18656 19712
rect 18604 19669 18613 19703
rect 18613 19669 18647 19703
rect 18647 19669 18656 19703
rect 18604 19660 18656 19669
rect 20904 19805 20913 19839
rect 20913 19805 20947 19839
rect 20947 19805 20956 19839
rect 20904 19796 20956 19805
rect 20720 19771 20772 19780
rect 20720 19737 20729 19771
rect 20729 19737 20763 19771
rect 20763 19737 20772 19771
rect 20720 19728 20772 19737
rect 22008 19796 22060 19848
rect 24032 19839 24084 19848
rect 24032 19805 24041 19839
rect 24041 19805 24075 19839
rect 24075 19805 24084 19839
rect 24032 19796 24084 19805
rect 26332 19728 26384 19780
rect 20444 19660 20496 19712
rect 22192 19660 22244 19712
rect 23112 19660 23164 19712
rect 24952 19660 25004 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1768 19456 1820 19508
rect 2136 19456 2188 19508
rect 7564 19456 7616 19508
rect 3056 19320 3108 19372
rect 8300 19456 8352 19508
rect 9496 19456 9548 19508
rect 12716 19499 12768 19508
rect 12716 19465 12725 19499
rect 12725 19465 12759 19499
rect 12759 19465 12768 19499
rect 12716 19456 12768 19465
rect 4528 19295 4580 19304
rect 4528 19261 4562 19295
rect 4562 19261 4580 19295
rect 2504 19184 2556 19236
rect 3240 19184 3292 19236
rect 4160 19184 4212 19236
rect 4528 19252 4580 19261
rect 5264 19252 5316 19304
rect 11520 19388 11572 19440
rect 16580 19456 16632 19508
rect 16856 19499 16908 19508
rect 16856 19465 16865 19499
rect 16865 19465 16899 19499
rect 16899 19465 16908 19499
rect 16856 19456 16908 19465
rect 17408 19499 17460 19508
rect 17408 19465 17417 19499
rect 17417 19465 17451 19499
rect 17451 19465 17460 19499
rect 17408 19456 17460 19465
rect 20260 19456 20312 19508
rect 21456 19456 21508 19508
rect 24952 19499 25004 19508
rect 24952 19465 24961 19499
rect 24961 19465 24995 19499
rect 24995 19465 25004 19499
rect 24952 19456 25004 19465
rect 15108 19431 15160 19440
rect 4988 19184 5040 19236
rect 11244 19320 11296 19372
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 15108 19397 15117 19431
rect 15117 19397 15151 19431
rect 15151 19397 15160 19431
rect 15108 19388 15160 19397
rect 11888 19320 11940 19329
rect 13268 19320 13320 19372
rect 13728 19363 13780 19372
rect 13728 19329 13737 19363
rect 13737 19329 13771 19363
rect 13771 19329 13780 19363
rect 13728 19320 13780 19329
rect 14556 19320 14608 19372
rect 15752 19320 15804 19372
rect 18972 19320 19024 19372
rect 7932 19184 7984 19236
rect 1952 19116 2004 19168
rect 3608 19116 3660 19168
rect 5632 19159 5684 19168
rect 5632 19125 5641 19159
rect 5641 19125 5675 19159
rect 5675 19125 5684 19159
rect 5632 19116 5684 19125
rect 6460 19116 6512 19168
rect 6736 19116 6788 19168
rect 6920 19116 6972 19168
rect 7472 19159 7524 19168
rect 7472 19125 7481 19159
rect 7481 19125 7515 19159
rect 7515 19125 7524 19159
rect 7472 19116 7524 19125
rect 10048 19116 10100 19168
rect 10784 19252 10836 19304
rect 12716 19252 12768 19304
rect 14096 19252 14148 19304
rect 15568 19295 15620 19304
rect 15568 19261 15577 19295
rect 15577 19261 15611 19295
rect 15611 19261 15620 19295
rect 15568 19252 15620 19261
rect 16948 19295 17000 19304
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 17960 19252 18012 19304
rect 19064 19295 19116 19304
rect 19064 19261 19073 19295
rect 19073 19261 19107 19295
rect 19107 19261 19116 19295
rect 19064 19252 19116 19261
rect 20076 19388 20128 19440
rect 20720 19388 20772 19440
rect 20444 19320 20496 19372
rect 21180 19320 21232 19372
rect 23112 19388 23164 19440
rect 22652 19363 22704 19372
rect 22652 19329 22661 19363
rect 22661 19329 22695 19363
rect 22695 19329 22704 19363
rect 22652 19320 22704 19329
rect 12256 19184 12308 19236
rect 12624 19184 12676 19236
rect 11060 19116 11112 19168
rect 13820 19184 13872 19236
rect 15844 19184 15896 19236
rect 18604 19184 18656 19236
rect 19524 19252 19576 19304
rect 20996 19252 21048 19304
rect 22100 19252 22152 19304
rect 23112 19295 23164 19304
rect 23112 19261 23121 19295
rect 23121 19261 23155 19295
rect 23155 19261 23164 19295
rect 24032 19388 24084 19440
rect 25136 19388 25188 19440
rect 25596 19320 25648 19372
rect 23112 19252 23164 19261
rect 24124 19252 24176 19304
rect 25136 19252 25188 19304
rect 19340 19184 19392 19236
rect 21272 19184 21324 19236
rect 22376 19227 22428 19236
rect 22376 19193 22385 19227
rect 22385 19193 22419 19227
rect 22419 19193 22428 19227
rect 22376 19184 22428 19193
rect 13544 19159 13596 19168
rect 13544 19125 13553 19159
rect 13553 19125 13587 19159
rect 13587 19125 13596 19159
rect 13544 19116 13596 19125
rect 13636 19159 13688 19168
rect 13636 19125 13645 19159
rect 13645 19125 13679 19159
rect 13679 19125 13688 19159
rect 14556 19159 14608 19168
rect 13636 19116 13688 19125
rect 14556 19125 14565 19159
rect 14565 19125 14599 19159
rect 14599 19125 14608 19159
rect 14556 19116 14608 19125
rect 16212 19159 16264 19168
rect 16212 19125 16221 19159
rect 16221 19125 16255 19159
rect 16255 19125 16264 19159
rect 16212 19116 16264 19125
rect 16488 19116 16540 19168
rect 17132 19159 17184 19168
rect 17132 19125 17141 19159
rect 17141 19125 17175 19159
rect 17175 19125 17184 19159
rect 17132 19116 17184 19125
rect 17776 19159 17828 19168
rect 17776 19125 17785 19159
rect 17785 19125 17819 19159
rect 17819 19125 17828 19159
rect 17776 19116 17828 19125
rect 18512 19159 18564 19168
rect 18512 19125 18521 19159
rect 18521 19125 18555 19159
rect 18555 19125 18564 19159
rect 18512 19116 18564 19125
rect 18696 19159 18748 19168
rect 18696 19125 18705 19159
rect 18705 19125 18739 19159
rect 18739 19125 18748 19159
rect 18696 19116 18748 19125
rect 19248 19116 19300 19168
rect 20260 19159 20312 19168
rect 20260 19125 20269 19159
rect 20269 19125 20303 19159
rect 20303 19125 20312 19159
rect 20260 19116 20312 19125
rect 20444 19116 20496 19168
rect 20904 19116 20956 19168
rect 21548 19116 21600 19168
rect 21732 19116 21784 19168
rect 24216 19116 24268 19168
rect 25688 19116 25740 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2780 18955 2832 18964
rect 2780 18921 2789 18955
rect 2789 18921 2823 18955
rect 2823 18921 2832 18955
rect 2780 18912 2832 18921
rect 4528 18912 4580 18964
rect 5448 18912 5500 18964
rect 8024 18955 8076 18964
rect 8024 18921 8033 18955
rect 8033 18921 8067 18955
rect 8067 18921 8076 18955
rect 8024 18912 8076 18921
rect 10048 18912 10100 18964
rect 11060 18912 11112 18964
rect 12808 18955 12860 18964
rect 2504 18844 2556 18896
rect 2596 18844 2648 18896
rect 3332 18844 3384 18896
rect 5632 18887 5684 18896
rect 1584 18776 1636 18828
rect 2412 18776 2464 18828
rect 4160 18776 4212 18828
rect 5632 18853 5666 18887
rect 5666 18853 5684 18887
rect 5632 18844 5684 18853
rect 7656 18844 7708 18896
rect 4988 18776 5040 18828
rect 6460 18776 6512 18828
rect 7564 18776 7616 18828
rect 8852 18776 8904 18828
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 11244 18844 11296 18896
rect 12808 18921 12817 18955
rect 12817 18921 12851 18955
rect 12851 18921 12860 18955
rect 12808 18912 12860 18921
rect 13268 18955 13320 18964
rect 13268 18921 13277 18955
rect 13277 18921 13311 18955
rect 13311 18921 13320 18955
rect 13268 18912 13320 18921
rect 13636 18912 13688 18964
rect 15108 18912 15160 18964
rect 15476 18955 15528 18964
rect 15476 18921 15485 18955
rect 15485 18921 15519 18955
rect 15519 18921 15528 18955
rect 15476 18912 15528 18921
rect 15660 18912 15712 18964
rect 17684 18912 17736 18964
rect 20076 18912 20128 18964
rect 22008 18912 22060 18964
rect 22652 18912 22704 18964
rect 24124 18912 24176 18964
rect 25228 18912 25280 18964
rect 13360 18844 13412 18896
rect 15844 18887 15896 18896
rect 15844 18853 15853 18887
rect 15853 18853 15887 18887
rect 15887 18853 15896 18887
rect 15844 18844 15896 18853
rect 21916 18844 21968 18896
rect 22560 18844 22612 18896
rect 23112 18844 23164 18896
rect 10784 18819 10836 18828
rect 10784 18785 10793 18819
rect 10793 18785 10827 18819
rect 10827 18785 10836 18819
rect 10784 18776 10836 18785
rect 11336 18776 11388 18828
rect 13176 18776 13228 18828
rect 13452 18776 13504 18828
rect 13728 18819 13780 18828
rect 13728 18785 13737 18819
rect 13737 18785 13771 18819
rect 13771 18785 13780 18819
rect 13728 18776 13780 18785
rect 15384 18776 15436 18828
rect 17408 18776 17460 18828
rect 19064 18776 19116 18828
rect 20260 18776 20312 18828
rect 20996 18776 21048 18828
rect 2504 18640 2556 18692
rect 7104 18640 7156 18692
rect 8668 18640 8720 18692
rect 13452 18640 13504 18692
rect 14556 18708 14608 18760
rect 15844 18708 15896 18760
rect 19432 18751 19484 18760
rect 19432 18717 19441 18751
rect 19441 18717 19475 18751
rect 19475 18717 19484 18751
rect 19432 18708 19484 18717
rect 21456 18751 21508 18760
rect 21456 18717 21465 18751
rect 21465 18717 21499 18751
rect 21499 18717 21508 18751
rect 21456 18708 21508 18717
rect 20076 18640 20128 18692
rect 20628 18640 20680 18692
rect 1952 18615 2004 18624
rect 1952 18581 1961 18615
rect 1961 18581 1995 18615
rect 1995 18581 2004 18615
rect 1952 18572 2004 18581
rect 3056 18572 3108 18624
rect 3240 18572 3292 18624
rect 3976 18572 4028 18624
rect 5264 18615 5316 18624
rect 5264 18581 5273 18615
rect 5273 18581 5307 18615
rect 5307 18581 5316 18615
rect 5264 18572 5316 18581
rect 6736 18572 6788 18624
rect 7840 18572 7892 18624
rect 7932 18615 7984 18624
rect 7932 18581 7941 18615
rect 7941 18581 7975 18615
rect 7975 18581 7984 18615
rect 9036 18615 9088 18624
rect 7932 18572 7984 18581
rect 9036 18581 9045 18615
rect 9045 18581 9079 18615
rect 9079 18581 9088 18615
rect 9036 18572 9088 18581
rect 13636 18572 13688 18624
rect 14372 18615 14424 18624
rect 14372 18581 14381 18615
rect 14381 18581 14415 18615
rect 14415 18581 14424 18615
rect 14372 18572 14424 18581
rect 17960 18572 18012 18624
rect 18880 18615 18932 18624
rect 18880 18581 18889 18615
rect 18889 18581 18923 18615
rect 18923 18581 18932 18615
rect 18880 18572 18932 18581
rect 20444 18572 20496 18624
rect 21548 18572 21600 18624
rect 23020 18776 23072 18828
rect 24124 18776 24176 18828
rect 24308 18776 24360 18828
rect 24952 18819 25004 18828
rect 24952 18785 24961 18819
rect 24961 18785 24995 18819
rect 24995 18785 25004 18819
rect 24952 18776 25004 18785
rect 22744 18572 22796 18624
rect 24216 18572 24268 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2872 18368 2924 18420
rect 4160 18411 4212 18420
rect 4160 18377 4169 18411
rect 4169 18377 4203 18411
rect 4203 18377 4212 18411
rect 4160 18368 4212 18377
rect 5540 18368 5592 18420
rect 6460 18368 6512 18420
rect 7104 18411 7156 18420
rect 7104 18377 7113 18411
rect 7113 18377 7147 18411
rect 7147 18377 7156 18411
rect 7104 18368 7156 18377
rect 8392 18368 8444 18420
rect 9680 18368 9732 18420
rect 10784 18368 10836 18420
rect 11152 18368 11204 18420
rect 13360 18368 13412 18420
rect 13728 18368 13780 18420
rect 4344 18300 4396 18352
rect 7840 18300 7892 18352
rect 8760 18300 8812 18352
rect 5264 18232 5316 18284
rect 1952 18207 2004 18216
rect 1952 18173 1961 18207
rect 1961 18173 1995 18207
rect 1995 18173 2004 18207
rect 1952 18164 2004 18173
rect 8116 18275 8168 18284
rect 8116 18241 8125 18275
rect 8125 18241 8159 18275
rect 8159 18241 8168 18275
rect 8116 18232 8168 18241
rect 8208 18275 8260 18284
rect 8208 18241 8217 18275
rect 8217 18241 8251 18275
rect 8251 18241 8260 18275
rect 8208 18232 8260 18241
rect 9588 18232 9640 18284
rect 9956 18300 10008 18352
rect 6736 18164 6788 18216
rect 7656 18164 7708 18216
rect 8944 18164 8996 18216
rect 11060 18164 11112 18216
rect 11244 18232 11296 18284
rect 11520 18232 11572 18284
rect 12624 18232 12676 18284
rect 14096 18368 14148 18420
rect 15844 18368 15896 18420
rect 17408 18411 17460 18420
rect 15016 18232 15068 18284
rect 17408 18377 17417 18411
rect 17417 18377 17451 18411
rect 17451 18377 17460 18411
rect 17408 18368 17460 18377
rect 18972 18368 19024 18420
rect 19432 18368 19484 18420
rect 21640 18411 21692 18420
rect 21640 18377 21649 18411
rect 21649 18377 21683 18411
rect 21683 18377 21692 18411
rect 21640 18368 21692 18377
rect 22744 18411 22796 18420
rect 22744 18377 22753 18411
rect 22753 18377 22787 18411
rect 22787 18377 22796 18411
rect 22744 18368 22796 18377
rect 23020 18411 23072 18420
rect 23020 18377 23029 18411
rect 23029 18377 23063 18411
rect 23063 18377 23072 18411
rect 23020 18368 23072 18377
rect 24216 18368 24268 18420
rect 25504 18368 25556 18420
rect 18328 18343 18380 18352
rect 18328 18309 18337 18343
rect 18337 18309 18371 18343
rect 18371 18309 18380 18343
rect 18328 18300 18380 18309
rect 23572 18300 23624 18352
rect 24400 18300 24452 18352
rect 24952 18300 25004 18352
rect 18512 18232 18564 18284
rect 21180 18232 21232 18284
rect 21640 18232 21692 18284
rect 24032 18232 24084 18284
rect 11612 18164 11664 18216
rect 13084 18164 13136 18216
rect 13728 18164 13780 18216
rect 3608 18096 3660 18148
rect 5448 18096 5500 18148
rect 7840 18096 7892 18148
rect 9404 18096 9456 18148
rect 3332 18071 3384 18080
rect 3332 18037 3341 18071
rect 3341 18037 3375 18071
rect 3375 18037 3384 18071
rect 3332 18028 3384 18037
rect 5172 18071 5224 18080
rect 5172 18037 5181 18071
rect 5181 18037 5215 18071
rect 5215 18037 5224 18071
rect 5172 18028 5224 18037
rect 5632 18071 5684 18080
rect 5632 18037 5641 18071
rect 5641 18037 5675 18071
rect 5675 18037 5684 18071
rect 5632 18028 5684 18037
rect 7472 18071 7524 18080
rect 7472 18037 7481 18071
rect 7481 18037 7515 18071
rect 7515 18037 7524 18071
rect 7472 18028 7524 18037
rect 7656 18071 7708 18080
rect 7656 18037 7665 18071
rect 7665 18037 7699 18071
rect 7699 18037 7708 18071
rect 7656 18028 7708 18037
rect 8852 18028 8904 18080
rect 11244 18071 11296 18080
rect 11244 18037 11253 18071
rect 11253 18037 11287 18071
rect 11287 18037 11296 18071
rect 11244 18028 11296 18037
rect 11336 18028 11388 18080
rect 14004 18096 14056 18148
rect 15660 18164 15712 18216
rect 18144 18207 18196 18216
rect 18144 18173 18153 18207
rect 18153 18173 18187 18207
rect 18187 18173 18196 18207
rect 18144 18164 18196 18173
rect 19248 18164 19300 18216
rect 23020 18164 23072 18216
rect 24124 18207 24176 18216
rect 24124 18173 24133 18207
rect 24133 18173 24167 18207
rect 24167 18173 24176 18207
rect 24124 18164 24176 18173
rect 24860 18164 24912 18216
rect 17316 18096 17368 18148
rect 20996 18096 21048 18148
rect 13084 18028 13136 18080
rect 16488 18071 16540 18080
rect 16488 18037 16497 18071
rect 16497 18037 16531 18071
rect 16531 18037 16540 18071
rect 16488 18028 16540 18037
rect 20904 18028 20956 18080
rect 22192 18096 22244 18148
rect 24676 18096 24728 18148
rect 22008 18071 22060 18080
rect 22008 18037 22017 18071
rect 22017 18037 22051 18071
rect 22051 18037 22060 18071
rect 22008 18028 22060 18037
rect 22376 18028 22428 18080
rect 24124 18028 24176 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1584 17867 1636 17876
rect 1584 17833 1593 17867
rect 1593 17833 1627 17867
rect 1627 17833 1636 17867
rect 1584 17824 1636 17833
rect 2596 17824 2648 17876
rect 5448 17824 5500 17876
rect 2780 17799 2832 17808
rect 2780 17765 2789 17799
rect 2789 17765 2823 17799
rect 2823 17765 2832 17799
rect 2780 17756 2832 17765
rect 3424 17756 3476 17808
rect 3608 17756 3660 17808
rect 7656 17824 7708 17876
rect 8208 17824 8260 17876
rect 9680 17824 9732 17876
rect 10876 17867 10928 17876
rect 10876 17833 10885 17867
rect 10885 17833 10919 17867
rect 10919 17833 10928 17867
rect 10876 17824 10928 17833
rect 11152 17867 11204 17876
rect 11152 17833 11161 17867
rect 11161 17833 11195 17867
rect 11195 17833 11204 17867
rect 11152 17824 11204 17833
rect 11520 17867 11572 17876
rect 11520 17833 11529 17867
rect 11529 17833 11563 17867
rect 11563 17833 11572 17867
rect 11520 17824 11572 17833
rect 12992 17824 13044 17876
rect 13452 17867 13504 17876
rect 13452 17833 13461 17867
rect 13461 17833 13495 17867
rect 13495 17833 13504 17867
rect 13452 17824 13504 17833
rect 13820 17824 13872 17876
rect 15108 17867 15160 17876
rect 15108 17833 15117 17867
rect 15117 17833 15151 17867
rect 15151 17833 15160 17867
rect 15108 17824 15160 17833
rect 15752 17824 15804 17876
rect 16396 17824 16448 17876
rect 18236 17867 18288 17876
rect 18236 17833 18245 17867
rect 18245 17833 18279 17867
rect 18279 17833 18288 17867
rect 18236 17824 18288 17833
rect 18788 17867 18840 17876
rect 18788 17833 18797 17867
rect 18797 17833 18831 17867
rect 18831 17833 18840 17867
rect 18788 17824 18840 17833
rect 19248 17867 19300 17876
rect 19248 17833 19257 17867
rect 19257 17833 19291 17867
rect 19291 17833 19300 17867
rect 19248 17824 19300 17833
rect 19984 17824 20036 17876
rect 21456 17824 21508 17876
rect 22560 17867 22612 17876
rect 22560 17833 22569 17867
rect 22569 17833 22603 17867
rect 22603 17833 22612 17867
rect 22560 17824 22612 17833
rect 23112 17824 23164 17876
rect 23296 17824 23348 17876
rect 24216 17824 24268 17876
rect 24400 17824 24452 17876
rect 25412 17867 25464 17876
rect 25412 17833 25421 17867
rect 25421 17833 25455 17867
rect 25455 17833 25464 17867
rect 25412 17824 25464 17833
rect 6828 17799 6880 17808
rect 3056 17688 3108 17740
rect 2872 17663 2924 17672
rect 2504 17552 2556 17604
rect 2320 17484 2372 17536
rect 2872 17629 2881 17663
rect 2881 17629 2915 17663
rect 2915 17629 2924 17663
rect 2872 17620 2924 17629
rect 3240 17620 3292 17672
rect 6828 17765 6837 17799
rect 6837 17765 6871 17799
rect 6871 17765 6880 17799
rect 6828 17756 6880 17765
rect 8944 17756 8996 17808
rect 14188 17799 14240 17808
rect 14188 17765 14197 17799
rect 14197 17765 14231 17799
rect 14231 17765 14240 17799
rect 14188 17756 14240 17765
rect 15292 17756 15344 17808
rect 16488 17756 16540 17808
rect 22008 17799 22060 17808
rect 4988 17688 5040 17740
rect 5080 17620 5132 17672
rect 6920 17663 6972 17672
rect 6920 17629 6929 17663
rect 6929 17629 6963 17663
rect 6963 17629 6972 17663
rect 6920 17620 6972 17629
rect 8300 17688 8352 17740
rect 12900 17688 12952 17740
rect 13636 17688 13688 17740
rect 17500 17688 17552 17740
rect 22008 17765 22017 17799
rect 22017 17765 22051 17799
rect 22051 17765 22060 17799
rect 22008 17756 22060 17765
rect 22652 17756 22704 17808
rect 19248 17688 19300 17740
rect 21180 17688 21232 17740
rect 21916 17688 21968 17740
rect 22744 17731 22796 17740
rect 22744 17697 22753 17731
rect 22753 17697 22787 17731
rect 22787 17697 22796 17731
rect 22744 17688 22796 17697
rect 24952 17688 25004 17740
rect 8484 17663 8536 17672
rect 5540 17552 5592 17604
rect 8484 17629 8493 17663
rect 8493 17629 8527 17663
rect 8527 17629 8536 17663
rect 8484 17620 8536 17629
rect 8576 17663 8628 17672
rect 8576 17629 8585 17663
rect 8585 17629 8619 17663
rect 8619 17629 8628 17663
rect 8576 17620 8628 17629
rect 8760 17552 8812 17604
rect 4528 17484 4580 17536
rect 4804 17484 4856 17536
rect 6460 17527 6512 17536
rect 6460 17493 6469 17527
rect 6469 17493 6503 17527
rect 6503 17493 6512 17527
rect 6460 17484 6512 17493
rect 8024 17527 8076 17536
rect 8024 17493 8033 17527
rect 8033 17493 8067 17527
rect 8067 17493 8076 17527
rect 8024 17484 8076 17493
rect 9404 17527 9456 17536
rect 9404 17493 9413 17527
rect 9413 17493 9447 17527
rect 9447 17493 9456 17527
rect 11152 17620 11204 17672
rect 13452 17620 13504 17672
rect 15016 17620 15068 17672
rect 13912 17595 13964 17604
rect 13912 17561 13921 17595
rect 13921 17561 13955 17595
rect 13955 17561 13964 17595
rect 13912 17552 13964 17561
rect 9404 17484 9456 17493
rect 12348 17484 12400 17536
rect 18604 17620 18656 17672
rect 20076 17620 20128 17672
rect 20352 17620 20404 17672
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 16764 17552 16816 17604
rect 19432 17552 19484 17604
rect 15660 17484 15712 17536
rect 16672 17527 16724 17536
rect 16672 17493 16681 17527
rect 16681 17493 16715 17527
rect 16715 17493 16724 17527
rect 16672 17484 16724 17493
rect 17592 17527 17644 17536
rect 17592 17493 17601 17527
rect 17601 17493 17635 17527
rect 17635 17493 17644 17527
rect 17592 17484 17644 17493
rect 19708 17527 19760 17536
rect 19708 17493 19717 17527
rect 19717 17493 19751 17527
rect 19751 17493 19760 17527
rect 19708 17484 19760 17493
rect 19984 17527 20036 17536
rect 19984 17493 19993 17527
rect 19993 17493 20027 17527
rect 20027 17493 20036 17527
rect 19984 17484 20036 17493
rect 20444 17484 20496 17536
rect 20628 17484 20680 17536
rect 24676 17527 24728 17536
rect 24676 17493 24685 17527
rect 24685 17493 24719 17527
rect 24719 17493 24728 17527
rect 24676 17484 24728 17493
rect 24860 17484 24912 17536
rect 25412 17484 25464 17536
rect 25964 17484 26016 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2780 17280 2832 17332
rect 3792 17280 3844 17332
rect 5080 17280 5132 17332
rect 5448 17280 5500 17332
rect 6828 17280 6880 17332
rect 8576 17280 8628 17332
rect 11152 17280 11204 17332
rect 13452 17280 13504 17332
rect 15292 17323 15344 17332
rect 15292 17289 15301 17323
rect 15301 17289 15335 17323
rect 15335 17289 15344 17323
rect 15292 17280 15344 17289
rect 15660 17280 15712 17332
rect 17500 17323 17552 17332
rect 17500 17289 17509 17323
rect 17509 17289 17543 17323
rect 17543 17289 17552 17323
rect 17500 17280 17552 17289
rect 18236 17280 18288 17332
rect 19156 17323 19208 17332
rect 19156 17289 19165 17323
rect 19165 17289 19199 17323
rect 19199 17289 19208 17323
rect 19156 17280 19208 17289
rect 21364 17280 21416 17332
rect 21640 17323 21692 17332
rect 21640 17289 21649 17323
rect 21649 17289 21683 17323
rect 21683 17289 21692 17323
rect 21640 17280 21692 17289
rect 22652 17280 22704 17332
rect 22744 17280 22796 17332
rect 23480 17323 23532 17332
rect 23480 17289 23489 17323
rect 23489 17289 23523 17323
rect 23523 17289 23532 17323
rect 23480 17280 23532 17289
rect 23664 17323 23716 17332
rect 23664 17289 23673 17323
rect 23673 17289 23707 17323
rect 23707 17289 23716 17323
rect 23664 17280 23716 17289
rect 25780 17280 25832 17332
rect 1584 17212 1636 17264
rect 1860 17212 1912 17264
rect 3884 17212 3936 17264
rect 4344 17212 4396 17264
rect 9680 17255 9732 17264
rect 1308 17144 1360 17196
rect 1492 17144 1544 17196
rect 1952 17144 2004 17196
rect 2136 17076 2188 17128
rect 1860 17008 1912 17060
rect 3332 17008 3384 17060
rect 3792 17008 3844 17060
rect 9680 17221 9689 17255
rect 9689 17221 9723 17255
rect 9723 17221 9732 17255
rect 9680 17212 9732 17221
rect 11244 17255 11296 17264
rect 11244 17221 11253 17255
rect 11253 17221 11287 17255
rect 11287 17221 11296 17255
rect 11244 17212 11296 17221
rect 4988 17144 5040 17196
rect 5448 17144 5500 17196
rect 5540 17144 5592 17196
rect 8760 17187 8812 17196
rect 8760 17153 8769 17187
rect 8769 17153 8803 17187
rect 8803 17153 8812 17187
rect 8760 17144 8812 17153
rect 9496 17144 9548 17196
rect 11060 17144 11112 17196
rect 16488 17144 16540 17196
rect 8208 17076 8260 17128
rect 9036 17076 9088 17128
rect 9680 17076 9732 17128
rect 9956 17076 10008 17128
rect 14372 17119 14424 17128
rect 14372 17085 14381 17119
rect 14381 17085 14415 17119
rect 14415 17085 14424 17119
rect 14372 17076 14424 17085
rect 16764 17119 16816 17128
rect 16764 17085 16773 17119
rect 16773 17085 16807 17119
rect 16807 17085 16816 17119
rect 16764 17076 16816 17085
rect 9496 17008 9548 17060
rect 11704 17008 11756 17060
rect 12532 17008 12584 17060
rect 16580 17008 16632 17060
rect 18420 17144 18472 17196
rect 18604 17187 18656 17196
rect 18604 17153 18613 17187
rect 18613 17153 18647 17187
rect 18647 17153 18656 17187
rect 18604 17144 18656 17153
rect 21640 17144 21692 17196
rect 22468 17119 22520 17128
rect 22468 17085 22477 17119
rect 22477 17085 22511 17119
rect 22511 17085 22520 17119
rect 22468 17076 22520 17085
rect 23664 17076 23716 17128
rect 24676 17076 24728 17128
rect 26148 17280 26200 17332
rect 19156 17008 19208 17060
rect 19708 17008 19760 17060
rect 20628 17008 20680 17060
rect 21732 17008 21784 17060
rect 22560 17008 22612 17060
rect 23756 17008 23808 17060
rect 25320 17008 25372 17060
rect 26148 17008 26200 17060
rect 1308 16940 1360 16992
rect 2044 16940 2096 16992
rect 3424 16983 3476 16992
rect 3424 16949 3433 16983
rect 3433 16949 3467 16983
rect 3467 16949 3476 16983
rect 3424 16940 3476 16949
rect 4160 16940 4212 16992
rect 4988 16983 5040 16992
rect 4988 16949 4997 16983
rect 4997 16949 5031 16983
rect 5031 16949 5040 16983
rect 4988 16940 5040 16949
rect 7012 16983 7064 16992
rect 7012 16949 7021 16983
rect 7021 16949 7055 16983
rect 7055 16949 7064 16983
rect 7012 16940 7064 16949
rect 8300 16983 8352 16992
rect 8300 16949 8309 16983
rect 8309 16949 8343 16983
rect 8343 16949 8352 16983
rect 8300 16940 8352 16949
rect 13452 16940 13504 16992
rect 14924 16983 14976 16992
rect 14924 16949 14933 16983
rect 14933 16949 14967 16983
rect 14967 16949 14976 16983
rect 14924 16940 14976 16949
rect 16396 16983 16448 16992
rect 16396 16949 16405 16983
rect 16405 16949 16439 16983
rect 16439 16949 16448 16983
rect 16396 16940 16448 16949
rect 16856 16983 16908 16992
rect 16856 16949 16865 16983
rect 16865 16949 16899 16983
rect 16899 16949 16908 16983
rect 16856 16940 16908 16949
rect 18052 16983 18104 16992
rect 18052 16949 18061 16983
rect 18061 16949 18095 16983
rect 18095 16949 18104 16983
rect 18052 16940 18104 16949
rect 20720 16940 20772 16992
rect 21272 16940 21324 16992
rect 22652 16983 22704 16992
rect 22652 16949 22661 16983
rect 22661 16949 22695 16983
rect 22695 16949 22704 16983
rect 22652 16940 22704 16949
rect 23112 16940 23164 16992
rect 24952 16940 25004 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2780 16779 2832 16788
rect 2780 16745 2789 16779
rect 2789 16745 2823 16779
rect 2823 16745 2832 16779
rect 3240 16779 3292 16788
rect 2780 16736 2832 16745
rect 3240 16745 3249 16779
rect 3249 16745 3283 16779
rect 3283 16745 3292 16779
rect 3240 16736 3292 16745
rect 3792 16779 3844 16788
rect 3792 16745 3801 16779
rect 3801 16745 3835 16779
rect 3835 16745 3844 16779
rect 3792 16736 3844 16745
rect 4160 16736 4212 16788
rect 5540 16736 5592 16788
rect 8300 16736 8352 16788
rect 9496 16779 9548 16788
rect 9496 16745 9505 16779
rect 9505 16745 9539 16779
rect 9539 16745 9548 16779
rect 9496 16736 9548 16745
rect 9956 16779 10008 16788
rect 9956 16745 9965 16779
rect 9965 16745 9999 16779
rect 9999 16745 10008 16779
rect 9956 16736 10008 16745
rect 12624 16736 12676 16788
rect 12808 16736 12860 16788
rect 14556 16779 14608 16788
rect 14556 16745 14565 16779
rect 14565 16745 14599 16779
rect 14599 16745 14608 16779
rect 14556 16736 14608 16745
rect 16396 16736 16448 16788
rect 18420 16736 18472 16788
rect 19248 16779 19300 16788
rect 19248 16745 19257 16779
rect 19257 16745 19291 16779
rect 19291 16745 19300 16779
rect 19248 16736 19300 16745
rect 19432 16736 19484 16788
rect 20260 16779 20312 16788
rect 20260 16745 20269 16779
rect 20269 16745 20303 16779
rect 20303 16745 20312 16779
rect 20260 16736 20312 16745
rect 20628 16779 20680 16788
rect 20628 16745 20637 16779
rect 20637 16745 20671 16779
rect 20671 16745 20680 16779
rect 20628 16736 20680 16745
rect 21272 16779 21324 16788
rect 2136 16711 2188 16720
rect 2136 16677 2145 16711
rect 2145 16677 2179 16711
rect 2179 16677 2188 16711
rect 2136 16668 2188 16677
rect 1676 16600 1728 16652
rect 3792 16600 3844 16652
rect 6092 16711 6144 16720
rect 6092 16677 6101 16711
rect 6101 16677 6135 16711
rect 6135 16677 6144 16711
rect 6092 16668 6144 16677
rect 6736 16668 6788 16720
rect 4804 16600 4856 16652
rect 11152 16668 11204 16720
rect 12900 16668 12952 16720
rect 14832 16668 14884 16720
rect 17500 16668 17552 16720
rect 18604 16711 18656 16720
rect 10324 16643 10376 16652
rect 10324 16609 10333 16643
rect 10333 16609 10367 16643
rect 10367 16609 10376 16643
rect 10324 16600 10376 16609
rect 12532 16643 12584 16652
rect 12532 16609 12541 16643
rect 12541 16609 12575 16643
rect 12575 16609 12584 16643
rect 12532 16600 12584 16609
rect 13176 16643 13228 16652
rect 13176 16609 13185 16643
rect 13185 16609 13219 16643
rect 13219 16609 13228 16643
rect 13176 16600 13228 16609
rect 13728 16600 13780 16652
rect 15108 16643 15160 16652
rect 15108 16609 15117 16643
rect 15117 16609 15151 16643
rect 15151 16609 15160 16643
rect 15108 16600 15160 16609
rect 16028 16643 16080 16652
rect 16028 16609 16037 16643
rect 16037 16609 16071 16643
rect 16071 16609 16080 16643
rect 16028 16600 16080 16609
rect 2780 16532 2832 16584
rect 6552 16575 6604 16584
rect 3516 16464 3568 16516
rect 2412 16439 2464 16448
rect 2412 16405 2421 16439
rect 2421 16405 2455 16439
rect 2455 16405 2464 16439
rect 2412 16396 2464 16405
rect 2780 16396 2832 16448
rect 6552 16541 6561 16575
rect 6561 16541 6595 16575
rect 6595 16541 6604 16575
rect 6552 16532 6604 16541
rect 13268 16575 13320 16584
rect 13268 16541 13277 16575
rect 13277 16541 13311 16575
rect 13311 16541 13320 16575
rect 13268 16532 13320 16541
rect 13452 16575 13504 16584
rect 13452 16541 13461 16575
rect 13461 16541 13495 16575
rect 13495 16541 13504 16575
rect 13452 16532 13504 16541
rect 13912 16532 13964 16584
rect 14648 16532 14700 16584
rect 15568 16532 15620 16584
rect 16396 16532 16448 16584
rect 16856 16600 16908 16652
rect 17132 16600 17184 16652
rect 17684 16575 17736 16584
rect 17684 16541 17693 16575
rect 17693 16541 17727 16575
rect 17727 16541 17736 16575
rect 17684 16532 17736 16541
rect 18604 16677 18613 16711
rect 18613 16677 18647 16711
rect 18647 16677 18656 16711
rect 18604 16668 18656 16677
rect 21272 16745 21281 16779
rect 21281 16745 21315 16779
rect 21315 16745 21324 16779
rect 21272 16736 21324 16745
rect 21916 16779 21968 16788
rect 21916 16745 21925 16779
rect 21925 16745 21959 16779
rect 21959 16745 21968 16779
rect 21916 16736 21968 16745
rect 22468 16779 22520 16788
rect 22468 16745 22477 16779
rect 22477 16745 22511 16779
rect 22511 16745 22520 16779
rect 22468 16736 22520 16745
rect 24676 16736 24728 16788
rect 25044 16779 25096 16788
rect 25044 16745 25053 16779
rect 25053 16745 25087 16779
rect 25087 16745 25096 16779
rect 25044 16736 25096 16745
rect 25688 16736 25740 16788
rect 20996 16668 21048 16720
rect 23296 16668 23348 16720
rect 24216 16668 24268 16720
rect 18972 16600 19024 16652
rect 19156 16643 19208 16652
rect 19156 16609 19165 16643
rect 19165 16609 19199 16643
rect 19199 16609 19208 16643
rect 19156 16600 19208 16609
rect 19616 16643 19668 16652
rect 19616 16609 19625 16643
rect 19625 16609 19659 16643
rect 19659 16609 19668 16643
rect 19616 16600 19668 16609
rect 22744 16643 22796 16652
rect 22744 16609 22753 16643
rect 22753 16609 22787 16643
rect 22787 16609 22796 16643
rect 22744 16600 22796 16609
rect 23756 16600 23808 16652
rect 23940 16600 23992 16652
rect 25320 16600 25372 16652
rect 5448 16439 5500 16448
rect 5448 16405 5457 16439
rect 5457 16405 5491 16439
rect 5491 16405 5500 16439
rect 5448 16396 5500 16405
rect 17868 16464 17920 16516
rect 19340 16464 19392 16516
rect 20720 16532 20772 16584
rect 20628 16464 20680 16516
rect 21456 16464 21508 16516
rect 23940 16464 23992 16516
rect 8116 16396 8168 16448
rect 11704 16439 11756 16448
rect 11704 16405 11713 16439
rect 11713 16405 11747 16439
rect 11747 16405 11756 16439
rect 11704 16396 11756 16405
rect 12808 16439 12860 16448
rect 12808 16405 12817 16439
rect 12817 16405 12851 16439
rect 12851 16405 12860 16439
rect 12808 16396 12860 16405
rect 15660 16439 15712 16448
rect 15660 16405 15669 16439
rect 15669 16405 15703 16439
rect 15703 16405 15712 16439
rect 15660 16396 15712 16405
rect 16764 16439 16816 16448
rect 16764 16405 16773 16439
rect 16773 16405 16807 16439
rect 16807 16405 16816 16439
rect 16764 16396 16816 16405
rect 17224 16439 17276 16448
rect 17224 16405 17233 16439
rect 17233 16405 17267 16439
rect 17267 16405 17276 16439
rect 17224 16396 17276 16405
rect 22652 16396 22704 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2044 16235 2096 16244
rect 2044 16201 2053 16235
rect 2053 16201 2087 16235
rect 2087 16201 2096 16235
rect 2044 16192 2096 16201
rect 2136 16192 2188 16244
rect 3424 16235 3476 16244
rect 3424 16201 3433 16235
rect 3433 16201 3467 16235
rect 3467 16201 3476 16235
rect 3424 16192 3476 16201
rect 5540 16192 5592 16244
rect 6736 16192 6788 16244
rect 9128 16192 9180 16244
rect 9680 16235 9732 16244
rect 3792 16124 3844 16176
rect 2504 16099 2556 16108
rect 2504 16065 2513 16099
rect 2513 16065 2547 16099
rect 2547 16065 2556 16099
rect 2504 16056 2556 16065
rect 2780 16056 2832 16108
rect 3884 16056 3936 16108
rect 6092 16056 6144 16108
rect 9680 16201 9689 16235
rect 9689 16201 9723 16235
rect 9723 16201 9732 16235
rect 9680 16192 9732 16201
rect 10324 16192 10376 16244
rect 10876 16192 10928 16244
rect 11152 16235 11204 16244
rect 11152 16201 11161 16235
rect 11161 16201 11195 16235
rect 11195 16201 11204 16235
rect 11152 16192 11204 16201
rect 11888 16235 11940 16244
rect 11888 16201 11897 16235
rect 11897 16201 11931 16235
rect 11931 16201 11940 16235
rect 11888 16192 11940 16201
rect 12348 16192 12400 16244
rect 13452 16235 13504 16244
rect 13452 16201 13461 16235
rect 13461 16201 13495 16235
rect 13495 16201 13504 16235
rect 13452 16192 13504 16201
rect 13820 16192 13872 16244
rect 14280 16192 14332 16244
rect 14556 16192 14608 16244
rect 16396 16235 16448 16244
rect 16396 16201 16405 16235
rect 16405 16201 16439 16235
rect 16439 16201 16448 16235
rect 16396 16192 16448 16201
rect 19064 16192 19116 16244
rect 20628 16192 20680 16244
rect 20904 16192 20956 16244
rect 16304 16167 16356 16176
rect 16304 16133 16313 16167
rect 16313 16133 16347 16167
rect 16347 16133 16356 16167
rect 16304 16124 16356 16133
rect 17868 16167 17920 16176
rect 17868 16133 17877 16167
rect 17877 16133 17911 16167
rect 17911 16133 17920 16167
rect 17868 16124 17920 16133
rect 18512 16124 18564 16176
rect 18696 16124 18748 16176
rect 3700 15988 3752 16040
rect 6552 15988 6604 16040
rect 11704 16056 11756 16108
rect 13176 16056 13228 16108
rect 13452 16056 13504 16108
rect 13820 16056 13872 16108
rect 16764 16056 16816 16108
rect 17500 16056 17552 16108
rect 11244 16031 11296 16040
rect 11244 15997 11253 16031
rect 11253 15997 11287 16031
rect 11287 15997 11296 16031
rect 11244 15988 11296 15997
rect 12808 16031 12860 16040
rect 12808 15997 12817 16031
rect 12817 15997 12851 16031
rect 12851 15997 12860 16031
rect 12808 15988 12860 15997
rect 17040 15988 17092 16040
rect 17684 15988 17736 16040
rect 2688 15920 2740 15972
rect 10968 15920 11020 15972
rect 12440 15920 12492 15972
rect 13728 15920 13780 15972
rect 13912 15920 13964 15972
rect 14924 15920 14976 15972
rect 16304 15920 16356 15972
rect 16672 15920 16724 15972
rect 19156 15920 19208 15972
rect 19432 15920 19484 15972
rect 20076 15920 20128 15972
rect 22468 16192 22520 16244
rect 22744 16235 22796 16244
rect 22744 16201 22753 16235
rect 22753 16201 22787 16235
rect 22787 16201 22796 16235
rect 22744 16192 22796 16201
rect 22100 16056 22152 16108
rect 23296 16192 23348 16244
rect 23664 16235 23716 16244
rect 23664 16201 23673 16235
rect 23673 16201 23707 16235
rect 23707 16201 23716 16235
rect 23664 16192 23716 16201
rect 24860 16192 24912 16244
rect 25504 16192 25556 16244
rect 25780 16192 25832 16244
rect 24032 16056 24084 16108
rect 22008 16031 22060 16040
rect 22008 15997 22017 16031
rect 22017 15997 22051 16031
rect 22051 15997 22060 16031
rect 22008 15988 22060 15997
rect 24860 15988 24912 16040
rect 26240 16031 26292 16040
rect 26240 15997 26249 16031
rect 26249 15997 26283 16031
rect 26283 15997 26292 16031
rect 26240 15988 26292 15997
rect 23940 15920 23992 15972
rect 25320 15920 25372 15972
rect 25872 15920 25924 15972
rect 1768 15852 1820 15904
rect 3332 15852 3384 15904
rect 4804 15852 4856 15904
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 5632 15895 5684 15904
rect 5632 15861 5641 15895
rect 5641 15861 5675 15895
rect 5675 15861 5684 15895
rect 5632 15852 5684 15861
rect 6552 15895 6604 15904
rect 6552 15861 6561 15895
rect 6561 15861 6595 15895
rect 6595 15861 6604 15895
rect 6552 15852 6604 15861
rect 6828 15852 6880 15904
rect 13820 15895 13872 15904
rect 13820 15861 13829 15895
rect 13829 15861 13863 15895
rect 13863 15861 13872 15895
rect 13820 15852 13872 15861
rect 14372 15895 14424 15904
rect 14372 15861 14381 15895
rect 14381 15861 14415 15895
rect 14415 15861 14424 15895
rect 14372 15852 14424 15861
rect 15568 15895 15620 15904
rect 15568 15861 15577 15895
rect 15577 15861 15611 15895
rect 15611 15861 15620 15895
rect 15568 15852 15620 15861
rect 17132 15852 17184 15904
rect 18144 15852 18196 15904
rect 23296 15852 23348 15904
rect 24032 15895 24084 15904
rect 24032 15861 24041 15895
rect 24041 15861 24075 15895
rect 24075 15861 24084 15895
rect 24032 15852 24084 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2504 15648 2556 15700
rect 3424 15648 3476 15700
rect 3884 15691 3936 15700
rect 3884 15657 3893 15691
rect 3893 15657 3927 15691
rect 3927 15657 3936 15691
rect 3884 15648 3936 15657
rect 2412 15512 2464 15564
rect 2688 15512 2740 15564
rect 4068 15580 4120 15632
rect 5448 15580 5500 15632
rect 5632 15648 5684 15700
rect 12164 15691 12216 15700
rect 12164 15657 12173 15691
rect 12173 15657 12207 15691
rect 12207 15657 12216 15691
rect 12164 15648 12216 15657
rect 13084 15648 13136 15700
rect 13360 15648 13412 15700
rect 13544 15648 13596 15700
rect 13728 15648 13780 15700
rect 14280 15691 14332 15700
rect 14280 15657 14289 15691
rect 14289 15657 14323 15691
rect 14323 15657 14332 15691
rect 14280 15648 14332 15657
rect 14648 15691 14700 15700
rect 14648 15657 14657 15691
rect 14657 15657 14691 15691
rect 14691 15657 14700 15691
rect 14648 15648 14700 15657
rect 17408 15648 17460 15700
rect 18052 15648 18104 15700
rect 18420 15648 18472 15700
rect 19340 15691 19392 15700
rect 19340 15657 19349 15691
rect 19349 15657 19383 15691
rect 19383 15657 19392 15691
rect 19340 15648 19392 15657
rect 20352 15691 20404 15700
rect 20352 15657 20361 15691
rect 20361 15657 20395 15691
rect 20395 15657 20404 15691
rect 20352 15648 20404 15657
rect 20628 15691 20680 15700
rect 20628 15657 20637 15691
rect 20637 15657 20671 15691
rect 20671 15657 20680 15691
rect 20628 15648 20680 15657
rect 21272 15648 21324 15700
rect 6736 15580 6788 15632
rect 7472 15580 7524 15632
rect 8116 15580 8168 15632
rect 8392 15623 8444 15632
rect 8392 15589 8401 15623
rect 8401 15589 8435 15623
rect 8435 15589 8444 15623
rect 8392 15580 8444 15589
rect 9864 15580 9916 15632
rect 11152 15580 11204 15632
rect 13268 15580 13320 15632
rect 4344 15512 4396 15564
rect 4804 15512 4856 15564
rect 6552 15512 6604 15564
rect 8300 15512 8352 15564
rect 10692 15512 10744 15564
rect 10876 15512 10928 15564
rect 15568 15512 15620 15564
rect 16396 15512 16448 15564
rect 1584 15444 1636 15496
rect 2044 15444 2096 15496
rect 2504 15444 2556 15496
rect 2780 15376 2832 15428
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 2412 15351 2464 15360
rect 2412 15317 2421 15351
rect 2421 15317 2455 15351
rect 2455 15317 2464 15351
rect 2412 15308 2464 15317
rect 8576 15487 8628 15496
rect 8576 15453 8585 15487
rect 8585 15453 8619 15487
rect 8619 15453 8628 15487
rect 8576 15444 8628 15453
rect 13544 15444 13596 15496
rect 13912 15487 13964 15496
rect 13912 15453 13921 15487
rect 13921 15453 13955 15487
rect 13955 15453 13964 15487
rect 13912 15444 13964 15453
rect 15108 15487 15160 15496
rect 15108 15453 15117 15487
rect 15117 15453 15151 15487
rect 15151 15453 15160 15487
rect 15108 15444 15160 15453
rect 6092 15419 6144 15428
rect 6092 15385 6101 15419
rect 6101 15385 6135 15419
rect 6135 15385 6144 15419
rect 6092 15376 6144 15385
rect 7748 15419 7800 15428
rect 7748 15385 7757 15419
rect 7757 15385 7791 15419
rect 7791 15385 7800 15419
rect 7748 15376 7800 15385
rect 8484 15376 8536 15428
rect 9312 15376 9364 15428
rect 9680 15376 9732 15428
rect 19248 15580 19300 15632
rect 20996 15580 21048 15632
rect 21180 15580 21232 15632
rect 21548 15648 21600 15700
rect 22100 15648 22152 15700
rect 22192 15648 22244 15700
rect 24032 15648 24084 15700
rect 25228 15648 25280 15700
rect 25504 15623 25556 15632
rect 25504 15589 25513 15623
rect 25513 15589 25547 15623
rect 25547 15589 25556 15623
rect 25504 15580 25556 15589
rect 17960 15512 18012 15564
rect 19340 15512 19392 15564
rect 19524 15512 19576 15564
rect 21916 15512 21968 15564
rect 22376 15512 22428 15564
rect 24952 15555 25004 15564
rect 24952 15521 24961 15555
rect 24961 15521 24995 15555
rect 24995 15521 25004 15555
rect 24952 15512 25004 15521
rect 18788 15487 18840 15496
rect 18236 15419 18288 15428
rect 18236 15385 18245 15419
rect 18245 15385 18279 15419
rect 18279 15385 18288 15419
rect 18236 15376 18288 15385
rect 18788 15453 18797 15487
rect 18797 15453 18831 15487
rect 18831 15453 18840 15487
rect 18788 15444 18840 15453
rect 20628 15444 20680 15496
rect 22468 15487 22520 15496
rect 22468 15453 22477 15487
rect 22477 15453 22511 15487
rect 22511 15453 22520 15487
rect 22468 15444 22520 15453
rect 20996 15376 21048 15428
rect 3700 15308 3752 15360
rect 3976 15308 4028 15360
rect 9036 15351 9088 15360
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 14096 15308 14148 15360
rect 15476 15351 15528 15360
rect 15476 15317 15485 15351
rect 15485 15317 15519 15351
rect 15519 15317 15528 15351
rect 15476 15308 15528 15317
rect 15568 15308 15620 15360
rect 17316 15308 17368 15360
rect 17500 15308 17552 15360
rect 18604 15308 18656 15360
rect 19892 15308 19944 15360
rect 21640 15308 21692 15360
rect 21824 15308 21876 15360
rect 22836 15308 22888 15360
rect 23480 15308 23532 15360
rect 24124 15308 24176 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2688 15104 2740 15156
rect 7196 15104 7248 15156
rect 8116 15147 8168 15156
rect 8116 15113 8125 15147
rect 8125 15113 8159 15147
rect 8159 15113 8168 15147
rect 8116 15104 8168 15113
rect 8300 15104 8352 15156
rect 9312 15104 9364 15156
rect 10876 15147 10928 15156
rect 10876 15113 10885 15147
rect 10885 15113 10919 15147
rect 10919 15113 10928 15147
rect 10876 15104 10928 15113
rect 11704 15104 11756 15156
rect 13728 15104 13780 15156
rect 14464 15147 14516 15156
rect 14464 15113 14473 15147
rect 14473 15113 14507 15147
rect 14507 15113 14516 15147
rect 14464 15104 14516 15113
rect 17224 15104 17276 15156
rect 17868 15104 17920 15156
rect 20260 15104 20312 15156
rect 21916 15147 21968 15156
rect 21916 15113 21925 15147
rect 21925 15113 21959 15147
rect 21959 15113 21968 15147
rect 21916 15104 21968 15113
rect 22100 15104 22152 15156
rect 22468 15104 22520 15156
rect 22560 15104 22612 15156
rect 24952 15147 25004 15156
rect 24952 15113 24961 15147
rect 24961 15113 24995 15147
rect 24995 15113 25004 15147
rect 24952 15104 25004 15113
rect 25964 15104 26016 15156
rect 2780 15036 2832 15088
rect 1492 14968 1544 15020
rect 1768 14968 1820 15020
rect 2320 14968 2372 15020
rect 3976 15036 4028 15088
rect 6552 15036 6604 15088
rect 3608 14968 3660 15020
rect 7564 15011 7616 15020
rect 7564 14977 7573 15011
rect 7573 14977 7607 15011
rect 7607 14977 7616 15011
rect 7564 14968 7616 14977
rect 1952 14900 2004 14952
rect 3148 14900 3200 14952
rect 4620 14900 4672 14952
rect 7196 14900 7248 14952
rect 4252 14875 4304 14884
rect 4252 14841 4286 14875
rect 4286 14841 4304 14875
rect 4252 14832 4304 14841
rect 4344 14832 4396 14884
rect 7748 14900 7800 14952
rect 10140 15036 10192 15088
rect 11244 15036 11296 15088
rect 11060 15011 11112 15020
rect 11060 14977 11069 15011
rect 11069 14977 11103 15011
rect 11103 14977 11112 15011
rect 11060 14968 11112 14977
rect 9588 14900 9640 14952
rect 10140 14900 10192 14952
rect 10600 14900 10652 14952
rect 14648 15036 14700 15088
rect 15476 15011 15528 15020
rect 15476 14977 15485 15011
rect 15485 14977 15519 15011
rect 15519 14977 15528 15011
rect 15476 14968 15528 14977
rect 17408 14968 17460 15020
rect 18512 15011 18564 15020
rect 18512 14977 18521 15011
rect 18521 14977 18555 15011
rect 18555 14977 18564 15011
rect 18512 14968 18564 14977
rect 18788 15036 18840 15088
rect 22376 15079 22428 15088
rect 22376 15045 22385 15079
rect 22385 15045 22419 15079
rect 22419 15045 22428 15079
rect 22376 15036 22428 15045
rect 22744 15036 22796 15088
rect 24032 15036 24084 15088
rect 26240 15079 26292 15088
rect 24124 15011 24176 15020
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 13084 14943 13136 14952
rect 8392 14832 8444 14884
rect 9036 14832 9088 14884
rect 13084 14909 13093 14943
rect 13093 14909 13127 14943
rect 13127 14909 13136 14943
rect 13084 14900 13136 14909
rect 13452 14900 13504 14952
rect 14004 14900 14056 14952
rect 14924 14900 14976 14952
rect 17040 14900 17092 14952
rect 19892 14900 19944 14952
rect 15752 14875 15804 14884
rect 15752 14841 15786 14875
rect 15786 14841 15804 14875
rect 15752 14832 15804 14841
rect 17868 14832 17920 14884
rect 22192 14900 22244 14952
rect 23480 14943 23532 14952
rect 23480 14909 23489 14943
rect 23489 14909 23523 14943
rect 23523 14909 23532 14943
rect 26240 15045 26249 15079
rect 26249 15045 26283 15079
rect 26283 15045 26292 15079
rect 26240 15036 26292 15045
rect 23480 14900 23532 14909
rect 20260 14875 20312 14884
rect 1492 14764 1544 14816
rect 2504 14764 2556 14816
rect 2872 14764 2924 14816
rect 3700 14764 3752 14816
rect 5172 14764 5224 14816
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 5356 14764 5408 14773
rect 5448 14764 5500 14816
rect 6368 14764 6420 14816
rect 7472 14764 7524 14816
rect 10048 14764 10100 14816
rect 10692 14764 10744 14816
rect 11152 14764 11204 14816
rect 12256 14807 12308 14816
rect 12256 14773 12265 14807
rect 12265 14773 12299 14807
rect 12299 14773 12308 14807
rect 12256 14764 12308 14773
rect 12624 14764 12676 14816
rect 13176 14764 13228 14816
rect 13820 14807 13872 14816
rect 13820 14773 13829 14807
rect 13829 14773 13863 14807
rect 13863 14773 13872 14807
rect 13820 14764 13872 14773
rect 16856 14807 16908 14816
rect 16856 14773 16865 14807
rect 16865 14773 16899 14807
rect 16899 14773 16908 14807
rect 16856 14764 16908 14773
rect 18052 14807 18104 14816
rect 18052 14773 18061 14807
rect 18061 14773 18095 14807
rect 18095 14773 18104 14807
rect 18052 14764 18104 14773
rect 18604 14764 18656 14816
rect 18696 14764 18748 14816
rect 20260 14841 20294 14875
rect 20294 14841 20312 14875
rect 20260 14832 20312 14841
rect 20812 14832 20864 14884
rect 21824 14832 21876 14884
rect 20444 14764 20496 14816
rect 22652 14807 22704 14816
rect 22652 14773 22661 14807
rect 22661 14773 22695 14807
rect 22695 14773 22704 14807
rect 22652 14764 22704 14773
rect 23664 14807 23716 14816
rect 23664 14773 23673 14807
rect 23673 14773 23707 14807
rect 23707 14773 23716 14807
rect 23664 14764 23716 14773
rect 24032 14807 24084 14816
rect 24032 14773 24041 14807
rect 24041 14773 24075 14807
rect 24075 14773 24084 14807
rect 24032 14764 24084 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 2412 14603 2464 14612
rect 2412 14569 2421 14603
rect 2421 14569 2455 14603
rect 2455 14569 2464 14603
rect 2412 14560 2464 14569
rect 2780 14560 2832 14612
rect 3056 14560 3108 14612
rect 4252 14560 4304 14612
rect 6184 14603 6236 14612
rect 6184 14569 6193 14603
rect 6193 14569 6227 14603
rect 6227 14569 6236 14603
rect 6184 14560 6236 14569
rect 6920 14560 6972 14612
rect 8024 14603 8076 14612
rect 8024 14569 8033 14603
rect 8033 14569 8067 14603
rect 8067 14569 8076 14603
rect 8024 14560 8076 14569
rect 8300 14560 8352 14612
rect 10140 14560 10192 14612
rect 10876 14603 10928 14612
rect 10876 14569 10885 14603
rect 10885 14569 10919 14603
rect 10919 14569 10928 14603
rect 10876 14560 10928 14569
rect 13360 14603 13412 14612
rect 13360 14569 13369 14603
rect 13369 14569 13403 14603
rect 13403 14569 13412 14603
rect 13360 14560 13412 14569
rect 13912 14603 13964 14612
rect 13912 14569 13921 14603
rect 13921 14569 13955 14603
rect 13955 14569 13964 14603
rect 13912 14560 13964 14569
rect 14280 14603 14332 14612
rect 14280 14569 14289 14603
rect 14289 14569 14323 14603
rect 14323 14569 14332 14603
rect 14280 14560 14332 14569
rect 14372 14560 14424 14612
rect 15108 14603 15160 14612
rect 15108 14569 15117 14603
rect 15117 14569 15151 14603
rect 15151 14569 15160 14603
rect 15108 14560 15160 14569
rect 15752 14560 15804 14612
rect 16580 14560 16632 14612
rect 17868 14603 17920 14612
rect 17868 14569 17877 14603
rect 17877 14569 17911 14603
rect 17911 14569 17920 14603
rect 17868 14560 17920 14569
rect 18420 14603 18472 14612
rect 18420 14569 18429 14603
rect 18429 14569 18463 14603
rect 18463 14569 18472 14603
rect 18420 14560 18472 14569
rect 19248 14603 19300 14612
rect 19248 14569 19257 14603
rect 19257 14569 19291 14603
rect 19291 14569 19300 14603
rect 19248 14560 19300 14569
rect 19524 14560 19576 14612
rect 21088 14603 21140 14612
rect 21088 14569 21097 14603
rect 21097 14569 21131 14603
rect 21131 14569 21140 14603
rect 21088 14560 21140 14569
rect 21272 14560 21324 14612
rect 22376 14560 22428 14612
rect 23480 14560 23532 14612
rect 24124 14560 24176 14612
rect 6368 14492 6420 14544
rect 7564 14492 7616 14544
rect 1768 14424 1820 14476
rect 1952 14424 2004 14476
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 4160 14424 4212 14476
rect 5356 14424 5408 14476
rect 6736 14467 6788 14476
rect 6736 14433 6745 14467
rect 6745 14433 6779 14467
rect 6779 14433 6788 14467
rect 6736 14424 6788 14433
rect 9128 14492 9180 14544
rect 12164 14492 12216 14544
rect 14556 14492 14608 14544
rect 15936 14535 15988 14544
rect 15936 14501 15945 14535
rect 15945 14501 15979 14535
rect 15979 14501 15988 14535
rect 15936 14492 15988 14501
rect 16396 14535 16448 14544
rect 16396 14501 16405 14535
rect 16405 14501 16439 14535
rect 16439 14501 16448 14535
rect 16396 14492 16448 14501
rect 16856 14492 16908 14544
rect 21364 14492 21416 14544
rect 22100 14492 22152 14544
rect 1860 14356 1912 14408
rect 2688 14356 2740 14408
rect 4252 14399 4304 14408
rect 4252 14365 4261 14399
rect 4261 14365 4295 14399
rect 4295 14365 4304 14399
rect 4252 14356 4304 14365
rect 11704 14424 11756 14476
rect 12532 14424 12584 14476
rect 12992 14424 13044 14476
rect 15476 14424 15528 14476
rect 16488 14467 16540 14476
rect 16488 14433 16497 14467
rect 16497 14433 16531 14467
rect 16531 14433 16540 14467
rect 16488 14424 16540 14433
rect 16764 14467 16816 14476
rect 16764 14433 16798 14467
rect 16798 14433 16816 14467
rect 16764 14424 16816 14433
rect 8668 14356 8720 14408
rect 9956 14356 10008 14408
rect 3608 14288 3660 14340
rect 6920 14331 6972 14340
rect 6920 14297 6929 14331
rect 6929 14297 6963 14331
rect 6963 14297 6972 14331
rect 6920 14288 6972 14297
rect 10876 14356 10928 14408
rect 11244 14399 11296 14408
rect 11244 14365 11253 14399
rect 11253 14365 11287 14399
rect 11287 14365 11296 14399
rect 11244 14356 11296 14365
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 18604 14356 18656 14408
rect 18972 14356 19024 14408
rect 19248 14356 19300 14408
rect 20076 14424 20128 14476
rect 20720 14424 20772 14476
rect 21456 14424 21508 14476
rect 23388 14424 23440 14476
rect 25504 14424 25556 14476
rect 20628 14399 20680 14408
rect 19156 14331 19208 14340
rect 19156 14297 19165 14331
rect 19165 14297 19199 14331
rect 19199 14297 19208 14331
rect 20628 14365 20637 14399
rect 20637 14365 20671 14399
rect 20671 14365 20680 14399
rect 20628 14356 20680 14365
rect 19156 14288 19208 14297
rect 20260 14288 20312 14340
rect 20536 14288 20588 14340
rect 1768 14220 1820 14272
rect 5540 14220 5592 14272
rect 6552 14263 6604 14272
rect 6552 14229 6561 14263
rect 6561 14229 6595 14263
rect 6595 14229 6604 14263
rect 6552 14220 6604 14229
rect 9588 14220 9640 14272
rect 10600 14220 10652 14272
rect 12348 14220 12400 14272
rect 20352 14263 20404 14272
rect 20352 14229 20361 14263
rect 20361 14229 20395 14263
rect 20395 14229 20404 14263
rect 20352 14220 20404 14229
rect 24952 14356 25004 14408
rect 26240 14399 26292 14408
rect 24032 14288 24084 14340
rect 25044 14288 25096 14340
rect 26240 14365 26249 14399
rect 26249 14365 26283 14399
rect 26283 14365 26292 14399
rect 26240 14356 26292 14365
rect 22652 14220 22704 14272
rect 24124 14220 24176 14272
rect 25780 14263 25832 14272
rect 25780 14229 25789 14263
rect 25789 14229 25823 14263
rect 25823 14229 25832 14263
rect 25780 14220 25832 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2044 14016 2096 14068
rect 2688 14059 2740 14068
rect 2688 14025 2697 14059
rect 2697 14025 2731 14059
rect 2731 14025 2740 14059
rect 2688 14016 2740 14025
rect 2780 14016 2832 14068
rect 1952 13880 2004 13932
rect 2044 13880 2096 13932
rect 3608 13948 3660 14000
rect 4988 13991 5040 14000
rect 2688 13812 2740 13864
rect 4988 13957 4997 13991
rect 4997 13957 5031 13991
rect 5031 13957 5040 13991
rect 4988 13948 5040 13957
rect 5172 13948 5224 14000
rect 5448 13923 5500 13932
rect 5448 13889 5457 13923
rect 5457 13889 5491 13923
rect 5491 13889 5500 13923
rect 5448 13880 5500 13889
rect 8484 14016 8536 14068
rect 10876 14016 10928 14068
rect 12256 14016 12308 14068
rect 12532 14016 12584 14068
rect 16488 14016 16540 14068
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 17776 14059 17828 14068
rect 17776 14025 17785 14059
rect 17785 14025 17819 14059
rect 17819 14025 17828 14059
rect 17776 14016 17828 14025
rect 18512 14016 18564 14068
rect 19248 14016 19300 14068
rect 19616 14016 19668 14068
rect 20812 14059 20864 14068
rect 8392 13991 8444 14000
rect 8392 13957 8401 13991
rect 8401 13957 8435 13991
rect 8435 13957 8444 13991
rect 8392 13948 8444 13957
rect 11704 13948 11756 14000
rect 14004 13991 14056 14000
rect 14004 13957 14013 13991
rect 14013 13957 14047 13991
rect 14047 13957 14056 13991
rect 14004 13948 14056 13957
rect 15292 13948 15344 14000
rect 6552 13880 6604 13932
rect 1952 13787 2004 13796
rect 1952 13753 1961 13787
rect 1961 13753 1995 13787
rect 1995 13753 2004 13787
rect 1952 13744 2004 13753
rect 2228 13744 2280 13796
rect 1860 13676 1912 13728
rect 3148 13676 3200 13728
rect 3792 13719 3844 13728
rect 3792 13685 3801 13719
rect 3801 13685 3835 13719
rect 3835 13685 3844 13719
rect 3792 13676 3844 13685
rect 6276 13676 6328 13728
rect 7748 13812 7800 13864
rect 9128 13812 9180 13864
rect 9588 13812 9640 13864
rect 12164 13880 12216 13932
rect 14464 13923 14516 13932
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 9496 13744 9548 13796
rect 10048 13744 10100 13796
rect 14464 13889 14473 13923
rect 14473 13889 14507 13923
rect 14507 13889 14516 13923
rect 14464 13880 14516 13889
rect 13728 13812 13780 13864
rect 16764 13880 16816 13932
rect 18880 13948 18932 14000
rect 20812 14025 20821 14059
rect 20821 14025 20855 14059
rect 20855 14025 20864 14059
rect 20812 14016 20864 14025
rect 21456 14059 21508 14068
rect 21456 14025 21465 14059
rect 21465 14025 21499 14059
rect 21499 14025 21508 14059
rect 21456 14016 21508 14025
rect 22008 14016 22060 14068
rect 22744 14016 22796 14068
rect 23480 14059 23532 14068
rect 23480 14025 23489 14059
rect 23489 14025 23523 14059
rect 23523 14025 23532 14059
rect 23480 14016 23532 14025
rect 24032 14016 24084 14068
rect 25412 14059 25464 14068
rect 25412 14025 25421 14059
rect 25421 14025 25455 14059
rect 25455 14025 25464 14059
rect 25412 14016 25464 14025
rect 26608 14016 26660 14068
rect 22376 13948 22428 14000
rect 18052 13880 18104 13932
rect 15476 13812 15528 13864
rect 20628 13880 20680 13932
rect 14096 13744 14148 13796
rect 17960 13744 18012 13796
rect 18512 13744 18564 13796
rect 20444 13812 20496 13864
rect 21364 13812 21416 13864
rect 22008 13880 22060 13932
rect 24124 13923 24176 13932
rect 24124 13889 24133 13923
rect 24133 13889 24167 13923
rect 24167 13889 24176 13923
rect 24124 13880 24176 13889
rect 25044 13948 25096 14000
rect 25228 13948 25280 14000
rect 24308 13880 24360 13932
rect 25412 13880 25464 13932
rect 25872 13880 25924 13932
rect 25228 13855 25280 13864
rect 20352 13744 20404 13796
rect 10692 13676 10744 13728
rect 10968 13676 11020 13728
rect 11060 13676 11112 13728
rect 12900 13676 12952 13728
rect 15936 13676 15988 13728
rect 18788 13676 18840 13728
rect 19156 13676 19208 13728
rect 20076 13676 20128 13728
rect 22100 13744 22152 13796
rect 25228 13821 25237 13855
rect 25237 13821 25271 13855
rect 25271 13821 25280 13855
rect 25228 13812 25280 13821
rect 25872 13744 25924 13796
rect 22652 13676 22704 13728
rect 24032 13719 24084 13728
rect 24032 13685 24041 13719
rect 24041 13685 24075 13719
rect 24075 13685 24084 13719
rect 24032 13676 24084 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1860 13472 1912 13524
rect 2228 13515 2280 13524
rect 2228 13481 2237 13515
rect 2237 13481 2271 13515
rect 2271 13481 2280 13515
rect 2228 13472 2280 13481
rect 2412 13472 2464 13524
rect 3148 13472 3200 13524
rect 4804 13515 4856 13524
rect 4804 13481 4813 13515
rect 4813 13481 4847 13515
rect 4847 13481 4856 13515
rect 4804 13472 4856 13481
rect 5172 13472 5224 13524
rect 7748 13515 7800 13524
rect 7748 13481 7757 13515
rect 7757 13481 7791 13515
rect 7791 13481 7800 13515
rect 7748 13472 7800 13481
rect 8116 13472 8168 13524
rect 8300 13515 8352 13524
rect 8300 13481 8309 13515
rect 8309 13481 8343 13515
rect 8343 13481 8352 13515
rect 8300 13472 8352 13481
rect 8668 13515 8720 13524
rect 8668 13481 8677 13515
rect 8677 13481 8711 13515
rect 8711 13481 8720 13515
rect 8668 13472 8720 13481
rect 9036 13515 9088 13524
rect 9036 13481 9045 13515
rect 9045 13481 9079 13515
rect 9079 13481 9088 13515
rect 9036 13472 9088 13481
rect 9496 13515 9548 13524
rect 9496 13481 9505 13515
rect 9505 13481 9539 13515
rect 9539 13481 9548 13515
rect 9496 13472 9548 13481
rect 10140 13472 10192 13524
rect 11244 13515 11296 13524
rect 11244 13481 11253 13515
rect 11253 13481 11287 13515
rect 11287 13481 11296 13515
rect 11244 13472 11296 13481
rect 11612 13515 11664 13524
rect 11612 13481 11621 13515
rect 11621 13481 11655 13515
rect 11655 13481 11664 13515
rect 11612 13472 11664 13481
rect 13176 13515 13228 13524
rect 13176 13481 13185 13515
rect 13185 13481 13219 13515
rect 13219 13481 13228 13515
rect 13176 13472 13228 13481
rect 13912 13515 13964 13524
rect 13912 13481 13921 13515
rect 13921 13481 13955 13515
rect 13955 13481 13964 13515
rect 13912 13472 13964 13481
rect 14188 13515 14240 13524
rect 14188 13481 14197 13515
rect 14197 13481 14231 13515
rect 14231 13481 14240 13515
rect 14188 13472 14240 13481
rect 16580 13472 16632 13524
rect 17868 13472 17920 13524
rect 19064 13515 19116 13524
rect 19064 13481 19073 13515
rect 19073 13481 19107 13515
rect 19107 13481 19116 13515
rect 19064 13472 19116 13481
rect 19248 13472 19300 13524
rect 21824 13472 21876 13524
rect 22008 13472 22060 13524
rect 24032 13472 24084 13524
rect 2044 13404 2096 13456
rect 2964 13404 3016 13456
rect 4344 13447 4396 13456
rect 4344 13413 4353 13447
rect 4353 13413 4387 13447
rect 4387 13413 4396 13447
rect 4344 13404 4396 13413
rect 6276 13404 6328 13456
rect 11520 13404 11572 13456
rect 13820 13404 13872 13456
rect 17316 13447 17368 13456
rect 2688 13336 2740 13388
rect 5448 13336 5500 13388
rect 6184 13336 6236 13388
rect 7196 13336 7248 13388
rect 9312 13336 9364 13388
rect 10876 13336 10928 13388
rect 11888 13336 11940 13388
rect 14096 13336 14148 13388
rect 14740 13336 14792 13388
rect 16304 13379 16356 13388
rect 16304 13345 16313 13379
rect 16313 13345 16347 13379
rect 16347 13345 16356 13379
rect 16304 13336 16356 13345
rect 17316 13413 17325 13447
rect 17325 13413 17359 13447
rect 17359 13413 17368 13447
rect 17316 13404 17368 13413
rect 18880 13404 18932 13456
rect 19800 13404 19852 13456
rect 17868 13379 17920 13388
rect 17868 13345 17877 13379
rect 17877 13345 17911 13379
rect 17911 13345 17920 13379
rect 17868 13336 17920 13345
rect 18420 13336 18472 13388
rect 19432 13379 19484 13388
rect 19432 13345 19441 13379
rect 19441 13345 19475 13379
rect 19475 13345 19484 13379
rect 19432 13336 19484 13345
rect 20628 13336 20680 13388
rect 1860 13268 1912 13320
rect 2136 13268 2188 13320
rect 4068 13268 4120 13320
rect 4988 13268 5040 13320
rect 5356 13311 5408 13320
rect 5356 13277 5365 13311
rect 5365 13277 5399 13311
rect 5399 13277 5408 13311
rect 5356 13268 5408 13277
rect 6276 13268 6328 13320
rect 9496 13268 9548 13320
rect 4160 13200 4212 13252
rect 5080 13200 5132 13252
rect 1676 13132 1728 13184
rect 6000 13132 6052 13184
rect 6184 13175 6236 13184
rect 6184 13141 6193 13175
rect 6193 13141 6227 13175
rect 6227 13141 6236 13175
rect 6184 13132 6236 13141
rect 10048 13200 10100 13252
rect 10600 13268 10652 13320
rect 11428 13268 11480 13320
rect 12256 13268 12308 13320
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 13728 13268 13780 13320
rect 14924 13311 14976 13320
rect 14924 13277 14933 13311
rect 14933 13277 14967 13311
rect 14967 13277 14976 13311
rect 14924 13268 14976 13277
rect 15292 13268 15344 13320
rect 17592 13268 17644 13320
rect 7288 13132 7340 13184
rect 11152 13132 11204 13184
rect 12808 13175 12860 13184
rect 12808 13141 12817 13175
rect 12817 13141 12851 13175
rect 12851 13141 12860 13175
rect 12808 13132 12860 13141
rect 16764 13200 16816 13252
rect 17500 13243 17552 13252
rect 17500 13209 17509 13243
rect 17509 13209 17543 13243
rect 17543 13209 17552 13243
rect 17500 13200 17552 13209
rect 22652 13404 22704 13456
rect 21456 13336 21508 13388
rect 22744 13336 22796 13388
rect 22284 13268 22336 13320
rect 22560 13268 22612 13320
rect 23388 13268 23440 13320
rect 24308 13336 24360 13388
rect 24584 13472 24636 13524
rect 24860 13472 24912 13524
rect 25320 13472 25372 13524
rect 25872 13515 25924 13524
rect 25872 13481 25881 13515
rect 25881 13481 25915 13515
rect 25915 13481 25924 13515
rect 25872 13472 25924 13481
rect 26240 13515 26292 13524
rect 26240 13481 26249 13515
rect 26249 13481 26283 13515
rect 26283 13481 26292 13515
rect 26240 13472 26292 13481
rect 24860 13336 24912 13388
rect 25044 13336 25096 13388
rect 19156 13200 19208 13252
rect 23480 13200 23532 13252
rect 25320 13268 25372 13320
rect 13912 13132 13964 13184
rect 14648 13175 14700 13184
rect 14648 13141 14657 13175
rect 14657 13141 14691 13175
rect 14691 13141 14700 13175
rect 14648 13132 14700 13141
rect 15752 13175 15804 13184
rect 15752 13141 15761 13175
rect 15761 13141 15795 13175
rect 15795 13141 15804 13175
rect 15752 13132 15804 13141
rect 15936 13175 15988 13184
rect 15936 13141 15945 13175
rect 15945 13141 15979 13175
rect 15979 13141 15988 13175
rect 15936 13132 15988 13141
rect 20812 13132 20864 13184
rect 22284 13175 22336 13184
rect 22284 13141 22293 13175
rect 22293 13141 22327 13175
rect 22327 13141 22336 13175
rect 22284 13132 22336 13141
rect 23848 13132 23900 13184
rect 24032 13132 24084 13184
rect 24952 13132 25004 13184
rect 25504 13175 25556 13184
rect 25504 13141 25513 13175
rect 25513 13141 25547 13175
rect 25547 13141 25556 13175
rect 25504 13132 25556 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1860 12971 1912 12980
rect 1860 12937 1869 12971
rect 1869 12937 1903 12971
rect 1903 12937 1912 12971
rect 1860 12928 1912 12937
rect 2044 12971 2096 12980
rect 2044 12937 2053 12971
rect 2053 12937 2087 12971
rect 2087 12937 2096 12971
rect 2044 12928 2096 12937
rect 2780 12928 2832 12980
rect 5356 12928 5408 12980
rect 8944 12928 8996 12980
rect 9496 12971 9548 12980
rect 9496 12937 9505 12971
rect 9505 12937 9539 12971
rect 9539 12937 9548 12971
rect 9496 12928 9548 12937
rect 10232 12928 10284 12980
rect 10692 12928 10744 12980
rect 11244 12928 11296 12980
rect 11612 12971 11664 12980
rect 11612 12937 11621 12971
rect 11621 12937 11655 12971
rect 11655 12937 11664 12971
rect 11612 12928 11664 12937
rect 12532 12928 12584 12980
rect 13268 12928 13320 12980
rect 14372 12971 14424 12980
rect 14372 12937 14381 12971
rect 14381 12937 14415 12971
rect 14415 12937 14424 12971
rect 14372 12928 14424 12937
rect 16120 12971 16172 12980
rect 16120 12937 16129 12971
rect 16129 12937 16163 12971
rect 16163 12937 16172 12971
rect 16120 12928 16172 12937
rect 16488 12928 16540 12980
rect 18420 12971 18472 12980
rect 2136 12860 2188 12912
rect 5448 12860 5500 12912
rect 4068 12792 4120 12844
rect 7012 12860 7064 12912
rect 8392 12903 8444 12912
rect 8392 12869 8401 12903
rect 8401 12869 8435 12903
rect 8435 12869 8444 12903
rect 8392 12860 8444 12869
rect 3792 12724 3844 12776
rect 4068 12699 4120 12708
rect 4068 12665 4077 12699
rect 4077 12665 4111 12699
rect 4111 12665 4120 12699
rect 4068 12656 4120 12665
rect 2412 12631 2464 12640
rect 2412 12597 2421 12631
rect 2421 12597 2455 12631
rect 2455 12597 2464 12631
rect 2412 12588 2464 12597
rect 2688 12588 2740 12640
rect 3608 12588 3660 12640
rect 6000 12792 6052 12844
rect 8484 12792 8536 12844
rect 5356 12724 5408 12776
rect 6092 12724 6144 12776
rect 6552 12724 6604 12776
rect 7288 12724 7340 12776
rect 8392 12724 8444 12776
rect 16304 12860 16356 12912
rect 10600 12835 10652 12844
rect 10600 12801 10609 12835
rect 10609 12801 10643 12835
rect 10643 12801 10652 12835
rect 10600 12792 10652 12801
rect 12808 12792 12860 12844
rect 9956 12724 10008 12776
rect 11244 12724 11296 12776
rect 13268 12724 13320 12776
rect 13912 12792 13964 12844
rect 14648 12792 14700 12844
rect 18420 12937 18429 12971
rect 18429 12937 18463 12971
rect 18463 12937 18472 12971
rect 18420 12928 18472 12937
rect 18880 12928 18932 12980
rect 19248 12928 19300 12980
rect 19800 12928 19852 12980
rect 20536 12928 20588 12980
rect 20720 12928 20772 12980
rect 20904 12928 20956 12980
rect 22744 12971 22796 12980
rect 22744 12937 22753 12971
rect 22753 12937 22787 12971
rect 22787 12937 22796 12971
rect 22744 12928 22796 12937
rect 23388 12928 23440 12980
rect 24124 12928 24176 12980
rect 24860 12928 24912 12980
rect 17500 12903 17552 12912
rect 17500 12869 17509 12903
rect 17509 12869 17543 12903
rect 17543 12869 17552 12903
rect 17500 12860 17552 12869
rect 17592 12860 17644 12912
rect 18328 12860 18380 12912
rect 21548 12860 21600 12912
rect 22008 12860 22060 12912
rect 22376 12860 22428 12912
rect 23296 12860 23348 12912
rect 23848 12860 23900 12912
rect 16764 12835 16816 12844
rect 16764 12801 16773 12835
rect 16773 12801 16807 12835
rect 16807 12801 16816 12835
rect 16764 12792 16816 12801
rect 19984 12792 20036 12844
rect 20260 12792 20312 12844
rect 20812 12792 20864 12844
rect 14372 12724 14424 12776
rect 16580 12767 16632 12776
rect 16580 12733 16589 12767
rect 16589 12733 16623 12767
rect 16623 12733 16632 12767
rect 16580 12724 16632 12733
rect 18972 12724 19024 12776
rect 19432 12724 19484 12776
rect 20168 12724 20220 12776
rect 20904 12724 20956 12776
rect 21180 12724 21232 12776
rect 22836 12792 22888 12844
rect 24492 12860 24544 12912
rect 25044 12903 25096 12912
rect 25044 12869 25053 12903
rect 25053 12869 25087 12903
rect 25087 12869 25096 12903
rect 25044 12860 25096 12869
rect 23112 12724 23164 12776
rect 23296 12724 23348 12776
rect 24032 12724 24084 12776
rect 5448 12588 5500 12640
rect 11888 12656 11940 12708
rect 5724 12588 5776 12640
rect 6276 12588 6328 12640
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 8852 12631 8904 12640
rect 8852 12597 8861 12631
rect 8861 12597 8895 12631
rect 8895 12597 8904 12631
rect 8852 12588 8904 12597
rect 10048 12588 10100 12640
rect 13452 12656 13504 12708
rect 14924 12699 14976 12708
rect 14924 12665 14933 12699
rect 14933 12665 14967 12699
rect 14967 12665 14976 12699
rect 14924 12656 14976 12665
rect 15568 12656 15620 12708
rect 19156 12699 19208 12708
rect 19156 12665 19190 12699
rect 19190 12665 19208 12699
rect 19156 12656 19208 12665
rect 19616 12656 19668 12708
rect 21732 12699 21784 12708
rect 21732 12665 21741 12699
rect 21741 12665 21775 12699
rect 21775 12665 21784 12699
rect 21732 12656 21784 12665
rect 22100 12656 22152 12708
rect 23480 12656 23532 12708
rect 24308 12724 24360 12776
rect 25044 12724 25096 12776
rect 13360 12631 13412 12640
rect 13360 12597 13369 12631
rect 13369 12597 13403 12631
rect 13403 12597 13412 12631
rect 13360 12588 13412 12597
rect 14556 12631 14608 12640
rect 14556 12597 14565 12631
rect 14565 12597 14599 12631
rect 14599 12597 14608 12631
rect 14556 12588 14608 12597
rect 16212 12631 16264 12640
rect 16212 12597 16221 12631
rect 16221 12597 16255 12631
rect 16255 12597 16264 12631
rect 16212 12588 16264 12597
rect 16304 12588 16356 12640
rect 16948 12588 17000 12640
rect 18420 12588 18472 12640
rect 20168 12588 20220 12640
rect 20720 12588 20772 12640
rect 20812 12588 20864 12640
rect 21088 12588 21140 12640
rect 25320 12588 25372 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2136 12427 2188 12436
rect 2136 12393 2145 12427
rect 2145 12393 2179 12427
rect 2179 12393 2188 12427
rect 2136 12384 2188 12393
rect 4252 12427 4304 12436
rect 4252 12393 4261 12427
rect 4261 12393 4295 12427
rect 4295 12393 4304 12427
rect 4252 12384 4304 12393
rect 5448 12384 5500 12436
rect 848 12316 900 12368
rect 2044 12316 2096 12368
rect 1768 12248 1820 12300
rect 3792 12316 3844 12368
rect 3148 12248 3200 12300
rect 5540 12316 5592 12368
rect 4068 12291 4120 12300
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 6000 12384 6052 12436
rect 6736 12384 6788 12436
rect 7012 12427 7064 12436
rect 7012 12393 7021 12427
rect 7021 12393 7055 12427
rect 7055 12393 7064 12427
rect 7012 12384 7064 12393
rect 6920 12316 6972 12368
rect 8208 12384 8260 12436
rect 9036 12427 9088 12436
rect 9036 12393 9045 12427
rect 9045 12393 9079 12427
rect 9079 12393 9088 12427
rect 9036 12384 9088 12393
rect 9312 12384 9364 12436
rect 9680 12384 9732 12436
rect 10048 12427 10100 12436
rect 10048 12393 10057 12427
rect 10057 12393 10091 12427
rect 10091 12393 10100 12427
rect 10048 12384 10100 12393
rect 11060 12384 11112 12436
rect 11428 12427 11480 12436
rect 11428 12393 11437 12427
rect 11437 12393 11471 12427
rect 11471 12393 11480 12427
rect 11428 12384 11480 12393
rect 11704 12427 11756 12436
rect 11704 12393 11713 12427
rect 11713 12393 11747 12427
rect 11747 12393 11756 12427
rect 11704 12384 11756 12393
rect 12256 12384 12308 12436
rect 14924 12384 14976 12436
rect 15200 12384 15252 12436
rect 15752 12384 15804 12436
rect 17868 12384 17920 12436
rect 18972 12427 19024 12436
rect 18972 12393 18981 12427
rect 18981 12393 19015 12427
rect 19015 12393 19024 12427
rect 18972 12384 19024 12393
rect 7564 12316 7616 12368
rect 19340 12384 19392 12436
rect 19432 12427 19484 12436
rect 19432 12393 19441 12427
rect 19441 12393 19475 12427
rect 19475 12393 19484 12427
rect 19432 12384 19484 12393
rect 21180 12384 21232 12436
rect 4068 12248 4120 12257
rect 2320 12180 2372 12232
rect 2596 12180 2648 12232
rect 3424 12180 3476 12232
rect 3884 12180 3936 12232
rect 4344 12180 4396 12232
rect 4620 12180 4672 12232
rect 2412 12155 2464 12164
rect 2412 12121 2421 12155
rect 2421 12121 2455 12155
rect 2455 12121 2464 12155
rect 2412 12112 2464 12121
rect 5356 12180 5408 12232
rect 1400 12044 1452 12096
rect 5448 12155 5500 12164
rect 5448 12121 5457 12155
rect 5457 12121 5491 12155
rect 5491 12121 5500 12155
rect 5448 12112 5500 12121
rect 6092 12248 6144 12300
rect 6828 12248 6880 12300
rect 7012 12248 7064 12300
rect 7288 12248 7340 12300
rect 6184 12180 6236 12232
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 4620 12087 4672 12096
rect 4620 12053 4629 12087
rect 4629 12053 4663 12087
rect 4663 12053 4672 12087
rect 4620 12044 4672 12053
rect 6460 12044 6512 12096
rect 7012 12044 7064 12096
rect 7288 12112 7340 12164
rect 7748 12248 7800 12300
rect 7932 12248 7984 12300
rect 8760 12248 8812 12300
rect 9404 12248 9456 12300
rect 9588 12248 9640 12300
rect 9864 12248 9916 12300
rect 10048 12248 10100 12300
rect 10876 12248 10928 12300
rect 12164 12291 12216 12300
rect 8208 12180 8260 12232
rect 8484 12180 8536 12232
rect 9312 12180 9364 12232
rect 10784 12223 10836 12232
rect 10784 12189 10793 12223
rect 10793 12189 10827 12223
rect 10827 12189 10836 12223
rect 10784 12180 10836 12189
rect 12164 12257 12198 12291
rect 12198 12257 12216 12291
rect 16580 12291 16632 12300
rect 12164 12248 12216 12257
rect 16580 12257 16589 12291
rect 16589 12257 16623 12291
rect 16623 12257 16632 12291
rect 16580 12248 16632 12257
rect 19064 12248 19116 12300
rect 20720 12359 20772 12368
rect 20720 12325 20729 12359
rect 20729 12325 20763 12359
rect 20763 12325 20772 12359
rect 20720 12316 20772 12325
rect 22100 12384 22152 12436
rect 23388 12427 23440 12436
rect 23388 12393 23397 12427
rect 23397 12393 23431 12427
rect 23431 12393 23440 12427
rect 23388 12384 23440 12393
rect 23756 12427 23808 12436
rect 23756 12393 23765 12427
rect 23765 12393 23799 12427
rect 23799 12393 23808 12427
rect 23756 12384 23808 12393
rect 23848 12427 23900 12436
rect 23848 12393 23857 12427
rect 23857 12393 23891 12427
rect 23891 12393 23900 12427
rect 24492 12427 24544 12436
rect 23848 12384 23900 12393
rect 24492 12393 24501 12427
rect 24501 12393 24535 12427
rect 24535 12393 24544 12427
rect 24492 12384 24544 12393
rect 24860 12384 24912 12436
rect 22652 12316 22704 12368
rect 23480 12316 23532 12368
rect 19432 12248 19484 12300
rect 21732 12248 21784 12300
rect 24952 12291 25004 12300
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 16672 12223 16724 12232
rect 16672 12189 16681 12223
rect 16681 12189 16715 12223
rect 16715 12189 16724 12223
rect 16672 12180 16724 12189
rect 17408 12180 17460 12232
rect 18052 12223 18104 12232
rect 18052 12189 18061 12223
rect 18061 12189 18095 12223
rect 18095 12189 18104 12223
rect 18052 12180 18104 12189
rect 18420 12180 18472 12232
rect 19248 12180 19300 12232
rect 19616 12180 19668 12232
rect 22284 12223 22336 12232
rect 9404 12112 9456 12164
rect 9956 12112 10008 12164
rect 19156 12112 19208 12164
rect 8024 12087 8076 12096
rect 8024 12053 8033 12087
rect 8033 12053 8067 12087
rect 8067 12053 8076 12087
rect 8024 12044 8076 12053
rect 13176 12044 13228 12096
rect 14188 12087 14240 12096
rect 14188 12053 14197 12087
rect 14197 12053 14231 12087
rect 14231 12053 14240 12087
rect 14188 12044 14240 12053
rect 15568 12087 15620 12096
rect 15568 12053 15577 12087
rect 15577 12053 15611 12087
rect 15611 12053 15620 12087
rect 15568 12044 15620 12053
rect 16212 12087 16264 12096
rect 16212 12053 16221 12087
rect 16221 12053 16255 12087
rect 16255 12053 16264 12087
rect 16212 12044 16264 12053
rect 19248 12044 19300 12096
rect 21088 12112 21140 12164
rect 21364 12112 21416 12164
rect 22284 12189 22293 12223
rect 22293 12189 22327 12223
rect 22327 12189 22336 12223
rect 22284 12180 22336 12189
rect 23480 12180 23532 12232
rect 24952 12257 24961 12291
rect 24961 12257 24995 12291
rect 24995 12257 25004 12291
rect 24952 12248 25004 12257
rect 25596 12291 25648 12300
rect 25596 12257 25605 12291
rect 25605 12257 25639 12291
rect 25639 12257 25648 12291
rect 25596 12248 25648 12257
rect 24032 12223 24084 12232
rect 24032 12189 24041 12223
rect 24041 12189 24075 12223
rect 24075 12189 24084 12223
rect 24032 12180 24084 12189
rect 25780 12180 25832 12232
rect 21824 12044 21876 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2596 11883 2648 11892
rect 2596 11849 2605 11883
rect 2605 11849 2639 11883
rect 2639 11849 2648 11883
rect 2596 11840 2648 11849
rect 3148 11840 3200 11892
rect 3516 11840 3568 11892
rect 1400 11636 1452 11688
rect 1952 11679 2004 11688
rect 1952 11645 1961 11679
rect 1961 11645 1995 11679
rect 1995 11645 2004 11679
rect 1952 11636 2004 11645
rect 2412 11636 2464 11688
rect 5540 11840 5592 11892
rect 6736 11840 6788 11892
rect 7012 11840 7064 11892
rect 8208 11883 8260 11892
rect 8208 11849 8217 11883
rect 8217 11849 8251 11883
rect 8251 11849 8260 11883
rect 8208 11840 8260 11849
rect 8576 11840 8628 11892
rect 9128 11883 9180 11892
rect 9128 11849 9137 11883
rect 9137 11849 9171 11883
rect 9171 11849 9180 11883
rect 9128 11840 9180 11849
rect 13912 11840 13964 11892
rect 15292 11883 15344 11892
rect 15292 11849 15301 11883
rect 15301 11849 15335 11883
rect 15335 11849 15344 11883
rect 15292 11840 15344 11849
rect 5356 11772 5408 11824
rect 6092 11772 6144 11824
rect 6276 11772 6328 11824
rect 3884 11568 3936 11620
rect 6276 11636 6328 11688
rect 9496 11704 9548 11756
rect 18972 11840 19024 11892
rect 21640 11840 21692 11892
rect 21824 11883 21876 11892
rect 21824 11849 21833 11883
rect 21833 11849 21867 11883
rect 21867 11849 21876 11883
rect 21824 11840 21876 11849
rect 22284 11840 22336 11892
rect 24032 11840 24084 11892
rect 24952 11883 25004 11892
rect 24952 11849 24961 11883
rect 24961 11849 24995 11883
rect 24995 11849 25004 11883
rect 24952 11840 25004 11849
rect 25412 11883 25464 11892
rect 25412 11849 25421 11883
rect 25421 11849 25455 11883
rect 25455 11849 25464 11883
rect 25412 11840 25464 11849
rect 4252 11568 4304 11620
rect 4804 11568 4856 11620
rect 7012 11568 7064 11620
rect 1768 11500 1820 11552
rect 4528 11543 4580 11552
rect 4528 11509 4537 11543
rect 4537 11509 4571 11543
rect 4571 11509 4580 11543
rect 4528 11500 4580 11509
rect 6184 11543 6236 11552
rect 6184 11509 6193 11543
rect 6193 11509 6227 11543
rect 6227 11509 6236 11543
rect 6184 11500 6236 11509
rect 7196 11500 7248 11552
rect 7748 11500 7800 11552
rect 10876 11500 10928 11552
rect 11888 11500 11940 11552
rect 14648 11636 14700 11688
rect 19524 11704 19576 11756
rect 19984 11704 20036 11756
rect 20904 11704 20956 11756
rect 21272 11747 21324 11756
rect 21272 11713 21281 11747
rect 21281 11713 21315 11747
rect 21315 11713 21324 11747
rect 21272 11704 21324 11713
rect 21456 11704 21508 11756
rect 16212 11636 16264 11688
rect 20720 11679 20772 11688
rect 20720 11645 20729 11679
rect 20729 11645 20763 11679
rect 20763 11645 20772 11679
rect 20720 11636 20772 11645
rect 13176 11568 13228 11620
rect 15568 11568 15620 11620
rect 19248 11568 19300 11620
rect 19616 11568 19668 11620
rect 13820 11500 13872 11552
rect 14188 11500 14240 11552
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 16856 11500 16908 11509
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 19156 11500 19208 11552
rect 19432 11543 19484 11552
rect 19432 11509 19441 11543
rect 19441 11509 19475 11543
rect 19475 11509 19484 11543
rect 19432 11500 19484 11509
rect 22100 11704 22152 11756
rect 22376 11747 22428 11756
rect 22376 11713 22385 11747
rect 22385 11713 22419 11747
rect 22419 11713 22428 11747
rect 22376 11704 22428 11713
rect 23480 11704 23532 11756
rect 26056 11840 26108 11892
rect 26240 11815 26292 11824
rect 26240 11781 26249 11815
rect 26249 11781 26283 11815
rect 26283 11781 26292 11815
rect 26240 11772 26292 11781
rect 23388 11500 23440 11552
rect 24032 11543 24084 11552
rect 24032 11509 24041 11543
rect 24041 11509 24075 11543
rect 24075 11509 24084 11543
rect 24032 11500 24084 11509
rect 24400 11500 24452 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1952 11339 2004 11348
rect 1952 11305 1961 11339
rect 1961 11305 1995 11339
rect 1995 11305 2004 11339
rect 1952 11296 2004 11305
rect 2044 11296 2096 11348
rect 2872 11339 2924 11348
rect 2872 11305 2881 11339
rect 2881 11305 2915 11339
rect 2915 11305 2924 11339
rect 2872 11296 2924 11305
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 4068 11296 4120 11348
rect 5356 11296 5408 11348
rect 6276 11296 6328 11348
rect 6828 11296 6880 11348
rect 7012 11296 7064 11348
rect 8208 11339 8260 11348
rect 1308 11228 1360 11280
rect 1860 11228 1912 11280
rect 4252 11160 4304 11212
rect 4528 11160 4580 11212
rect 5448 11160 5500 11212
rect 6460 11228 6512 11280
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 3148 11092 3200 11144
rect 6184 11092 6236 11144
rect 8208 11305 8217 11339
rect 8217 11305 8251 11339
rect 8251 11305 8260 11339
rect 8208 11296 8260 11305
rect 8300 11296 8352 11348
rect 9496 11296 9548 11348
rect 11612 11296 11664 11348
rect 12164 11296 12216 11348
rect 12716 11339 12768 11348
rect 12716 11305 12725 11339
rect 12725 11305 12759 11339
rect 12759 11305 12768 11339
rect 12716 11296 12768 11305
rect 13268 11296 13320 11348
rect 13544 11296 13596 11348
rect 14280 11296 14332 11348
rect 15660 11296 15712 11348
rect 17408 11296 17460 11348
rect 19156 11296 19208 11348
rect 20720 11296 20772 11348
rect 20904 11339 20956 11348
rect 20904 11305 20913 11339
rect 20913 11305 20947 11339
rect 20947 11305 20956 11339
rect 20904 11296 20956 11305
rect 21272 11339 21324 11348
rect 21272 11305 21281 11339
rect 21281 11305 21315 11339
rect 21315 11305 21324 11339
rect 21272 11296 21324 11305
rect 22008 11339 22060 11348
rect 22008 11305 22017 11339
rect 22017 11305 22051 11339
rect 22051 11305 22060 11339
rect 22008 11296 22060 11305
rect 22468 11339 22520 11348
rect 22468 11305 22477 11339
rect 22477 11305 22511 11339
rect 22511 11305 22520 11339
rect 22468 11296 22520 11305
rect 23848 11296 23900 11348
rect 24216 11296 24268 11348
rect 24860 11296 24912 11348
rect 10876 11228 10928 11280
rect 15936 11271 15988 11280
rect 15936 11237 15945 11271
rect 15945 11237 15979 11271
rect 15979 11237 15988 11271
rect 15936 11228 15988 11237
rect 16856 11228 16908 11280
rect 19432 11228 19484 11280
rect 22376 11271 22428 11280
rect 7380 11160 7432 11212
rect 8208 11160 8260 11212
rect 10416 11203 10468 11212
rect 10416 11169 10425 11203
rect 10425 11169 10459 11203
rect 10459 11169 10468 11203
rect 10416 11160 10468 11169
rect 11888 11160 11940 11212
rect 15292 11203 15344 11212
rect 15292 11169 15301 11203
rect 15301 11169 15335 11203
rect 15335 11169 15344 11203
rect 15292 11160 15344 11169
rect 15476 11160 15528 11212
rect 16304 11160 16356 11212
rect 18972 11160 19024 11212
rect 19708 11160 19760 11212
rect 19892 11160 19944 11212
rect 20352 11160 20404 11212
rect 22376 11237 22385 11271
rect 22385 11237 22419 11271
rect 22419 11237 22428 11271
rect 22376 11228 22428 11237
rect 23572 11228 23624 11280
rect 12992 11092 13044 11144
rect 14740 11135 14792 11144
rect 2136 11024 2188 11076
rect 6092 11024 6144 11076
rect 8116 11024 8168 11076
rect 3792 10999 3844 11008
rect 3792 10965 3801 10999
rect 3801 10965 3835 10999
rect 3835 10965 3844 10999
rect 3792 10956 3844 10965
rect 9036 10999 9088 11008
rect 9036 10965 9045 10999
rect 9045 10965 9079 10999
rect 9079 10965 9088 10999
rect 9036 10956 9088 10965
rect 12164 10956 12216 11008
rect 12440 10956 12492 11008
rect 14740 11101 14749 11135
rect 14749 11101 14783 11135
rect 14783 11101 14792 11135
rect 14740 11092 14792 11101
rect 16212 11092 16264 11144
rect 16396 11092 16448 11144
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 18880 11067 18932 11076
rect 18880 11033 18889 11067
rect 18889 11033 18923 11067
rect 18923 11033 18932 11067
rect 21088 11092 21140 11144
rect 22744 11160 22796 11212
rect 24216 11160 24268 11212
rect 22008 11092 22060 11144
rect 22928 11135 22980 11144
rect 22928 11101 22937 11135
rect 22937 11101 22971 11135
rect 22971 11101 22980 11135
rect 22928 11092 22980 11101
rect 23204 11092 23256 11144
rect 23480 11092 23532 11144
rect 24032 11092 24084 11144
rect 18880 11024 18932 11033
rect 21824 11024 21876 11076
rect 24400 11024 24452 11076
rect 14188 10956 14240 11008
rect 18420 10999 18472 11008
rect 18420 10965 18429 10999
rect 18429 10965 18463 10999
rect 18463 10965 18472 10999
rect 18420 10956 18472 10965
rect 19800 10956 19852 11008
rect 20628 10956 20680 11008
rect 23112 10956 23164 11008
rect 23480 10956 23532 11008
rect 24032 10956 24084 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 4252 10752 4304 10804
rect 4988 10795 5040 10804
rect 4988 10761 4997 10795
rect 4997 10761 5031 10795
rect 5031 10761 5040 10795
rect 4988 10752 5040 10761
rect 5540 10752 5592 10804
rect 6828 10752 6880 10804
rect 7288 10795 7340 10804
rect 5172 10727 5224 10736
rect 5172 10693 5181 10727
rect 5181 10693 5215 10727
rect 5215 10693 5224 10727
rect 5172 10684 5224 10693
rect 5356 10684 5408 10736
rect 7012 10684 7064 10736
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 7288 10761 7297 10795
rect 7297 10761 7331 10795
rect 7331 10761 7340 10795
rect 7288 10752 7340 10761
rect 10416 10795 10468 10804
rect 10416 10761 10425 10795
rect 10425 10761 10459 10795
rect 10459 10761 10468 10795
rect 10416 10752 10468 10761
rect 11612 10795 11664 10804
rect 11612 10761 11621 10795
rect 11621 10761 11655 10795
rect 11655 10761 11664 10795
rect 11612 10752 11664 10761
rect 11888 10795 11940 10804
rect 11888 10761 11897 10795
rect 11897 10761 11931 10795
rect 11931 10761 11940 10795
rect 11888 10752 11940 10761
rect 12992 10795 13044 10804
rect 12992 10761 13001 10795
rect 13001 10761 13035 10795
rect 13035 10761 13044 10795
rect 12992 10752 13044 10761
rect 13544 10752 13596 10804
rect 18972 10752 19024 10804
rect 19432 10795 19484 10804
rect 19432 10761 19441 10795
rect 19441 10761 19475 10795
rect 19475 10761 19484 10795
rect 19432 10752 19484 10761
rect 20168 10752 20220 10804
rect 8024 10616 8076 10668
rect 9036 10616 9088 10668
rect 10968 10659 11020 10668
rect 3792 10548 3844 10600
rect 4712 10548 4764 10600
rect 7932 10548 7984 10600
rect 10968 10625 10977 10659
rect 10977 10625 11011 10659
rect 11011 10625 11020 10659
rect 10968 10616 11020 10625
rect 17868 10684 17920 10736
rect 22100 10752 22152 10804
rect 22560 10752 22612 10804
rect 22652 10752 22704 10804
rect 23204 10752 23256 10804
rect 23756 10752 23808 10804
rect 24768 10795 24820 10804
rect 24768 10761 24777 10795
rect 24777 10761 24811 10795
rect 24811 10761 24820 10795
rect 24768 10752 24820 10761
rect 25596 10795 25648 10804
rect 25596 10761 25605 10795
rect 25605 10761 25639 10795
rect 25639 10761 25648 10795
rect 25596 10752 25648 10761
rect 20444 10684 20496 10736
rect 24584 10684 24636 10736
rect 13820 10659 13872 10668
rect 13820 10625 13829 10659
rect 13829 10625 13863 10659
rect 13863 10625 13872 10659
rect 13820 10616 13872 10625
rect 15568 10616 15620 10668
rect 17408 10659 17460 10668
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 18420 10616 18472 10668
rect 19892 10616 19944 10668
rect 20168 10616 20220 10668
rect 20628 10616 20680 10668
rect 21456 10616 21508 10668
rect 21548 10616 21600 10668
rect 22008 10616 22060 10668
rect 22376 10616 22428 10668
rect 22744 10616 22796 10668
rect 10876 10548 10928 10600
rect 16212 10591 16264 10600
rect 16212 10557 16221 10591
rect 16221 10557 16255 10591
rect 16255 10557 16264 10591
rect 16212 10548 16264 10557
rect 17776 10548 17828 10600
rect 18236 10548 18288 10600
rect 2044 10523 2096 10532
rect 2044 10489 2053 10523
rect 2053 10489 2087 10523
rect 2087 10489 2096 10523
rect 2044 10480 2096 10489
rect 2780 10480 2832 10532
rect 3240 10480 3292 10532
rect 4804 10480 4856 10532
rect 3884 10412 3936 10464
rect 5724 10412 5776 10464
rect 6368 10412 6420 10464
rect 7288 10412 7340 10464
rect 8208 10412 8260 10464
rect 8484 10412 8536 10464
rect 8760 10455 8812 10464
rect 8760 10421 8769 10455
rect 8769 10421 8803 10455
rect 8803 10421 8812 10455
rect 8760 10412 8812 10421
rect 9588 10412 9640 10464
rect 12348 10480 12400 10532
rect 14188 10523 14240 10532
rect 14188 10489 14222 10523
rect 14222 10489 14240 10523
rect 14188 10480 14240 10489
rect 16764 10523 16816 10532
rect 16764 10489 16773 10523
rect 16773 10489 16807 10523
rect 16807 10489 16816 10523
rect 16764 10480 16816 10489
rect 18144 10480 18196 10532
rect 18788 10480 18840 10532
rect 20904 10480 20956 10532
rect 21088 10480 21140 10532
rect 10876 10455 10928 10464
rect 10876 10421 10885 10455
rect 10885 10421 10919 10455
rect 10919 10421 10928 10455
rect 10876 10412 10928 10421
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 14740 10412 14792 10464
rect 15568 10412 15620 10464
rect 16304 10412 16356 10464
rect 18052 10455 18104 10464
rect 18052 10421 18061 10455
rect 18061 10421 18095 10455
rect 18095 10421 18104 10455
rect 18052 10412 18104 10421
rect 18236 10412 18288 10464
rect 18420 10455 18472 10464
rect 18420 10421 18429 10455
rect 18429 10421 18463 10455
rect 18463 10421 18472 10455
rect 18420 10412 18472 10421
rect 19248 10412 19300 10464
rect 19432 10412 19484 10464
rect 19984 10455 20036 10464
rect 19984 10421 19993 10455
rect 19993 10421 20027 10455
rect 20027 10421 20036 10455
rect 19984 10412 20036 10421
rect 21640 10480 21692 10532
rect 22560 10548 22612 10600
rect 22928 10591 22980 10600
rect 22928 10557 22937 10591
rect 22937 10557 22971 10591
rect 22971 10557 22980 10591
rect 22928 10548 22980 10557
rect 24768 10548 24820 10600
rect 24032 10480 24084 10532
rect 22284 10412 22336 10464
rect 23848 10412 23900 10464
rect 24216 10412 24268 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 2688 10208 2740 10260
rect 2872 10208 2924 10260
rect 3332 10208 3384 10260
rect 4712 10208 4764 10260
rect 5908 10251 5960 10260
rect 5908 10217 5917 10251
rect 5917 10217 5951 10251
rect 5951 10217 5960 10251
rect 5908 10208 5960 10217
rect 6460 10251 6512 10260
rect 6460 10217 6469 10251
rect 6469 10217 6503 10251
rect 6503 10217 6512 10251
rect 6460 10208 6512 10217
rect 9496 10208 9548 10260
rect 9680 10208 9732 10260
rect 10876 10208 10928 10260
rect 11152 10208 11204 10260
rect 11980 10208 12032 10260
rect 13452 10251 13504 10260
rect 13452 10217 13461 10251
rect 13461 10217 13495 10251
rect 13495 10217 13504 10251
rect 13452 10208 13504 10217
rect 13820 10208 13872 10260
rect 15384 10208 15436 10260
rect 15752 10251 15804 10260
rect 15752 10217 15761 10251
rect 15761 10217 15795 10251
rect 15795 10217 15804 10251
rect 15752 10208 15804 10217
rect 16396 10208 16448 10260
rect 16580 10208 16632 10260
rect 19432 10208 19484 10260
rect 19984 10251 20036 10260
rect 19984 10217 19993 10251
rect 19993 10217 20027 10251
rect 20027 10217 20036 10251
rect 19984 10208 20036 10217
rect 20812 10208 20864 10260
rect 21272 10208 21324 10260
rect 21548 10208 21600 10260
rect 22008 10208 22060 10260
rect 22468 10251 22520 10260
rect 22468 10217 22477 10251
rect 22477 10217 22511 10251
rect 22511 10217 22520 10251
rect 22468 10208 22520 10217
rect 23756 10251 23808 10260
rect 23756 10217 23765 10251
rect 23765 10217 23799 10251
rect 23799 10217 23808 10251
rect 23756 10208 23808 10217
rect 24032 10208 24084 10260
rect 24768 10251 24820 10260
rect 24768 10217 24777 10251
rect 24777 10217 24811 10251
rect 24811 10217 24820 10251
rect 24768 10208 24820 10217
rect 25044 10251 25096 10260
rect 25044 10217 25053 10251
rect 25053 10217 25087 10251
rect 25087 10217 25096 10251
rect 25044 10208 25096 10217
rect 25780 10251 25832 10260
rect 25780 10217 25789 10251
rect 25789 10217 25823 10251
rect 25823 10217 25832 10251
rect 25780 10208 25832 10217
rect 3148 10140 3200 10192
rect 2688 10072 2740 10124
rect 3148 10004 3200 10056
rect 2964 9936 3016 9988
rect 3332 9936 3384 9988
rect 5080 10140 5132 10192
rect 5540 10140 5592 10192
rect 11060 10140 11112 10192
rect 12900 10140 12952 10192
rect 13728 10140 13780 10192
rect 17960 10140 18012 10192
rect 4712 10072 4764 10124
rect 5816 10072 5868 10124
rect 7932 10072 7984 10124
rect 9220 10072 9272 10124
rect 10324 10072 10376 10124
rect 10600 10072 10652 10124
rect 6368 10004 6420 10056
rect 4344 9936 4396 9988
rect 5724 9936 5776 9988
rect 6276 9936 6328 9988
rect 7380 10004 7432 10056
rect 7656 9979 7708 9988
rect 7656 9945 7665 9979
rect 7665 9945 7699 9979
rect 7699 9945 7708 9979
rect 7656 9936 7708 9945
rect 8024 9936 8076 9988
rect 8576 10004 8628 10056
rect 10968 10047 11020 10056
rect 10968 10013 10977 10047
rect 10977 10013 11011 10047
rect 11011 10013 11020 10047
rect 10968 10004 11020 10013
rect 12992 10072 13044 10124
rect 13820 10115 13872 10124
rect 12348 10004 12400 10056
rect 12532 10047 12584 10056
rect 12532 10013 12541 10047
rect 12541 10013 12575 10047
rect 12575 10013 12584 10047
rect 12532 10004 12584 10013
rect 13176 10004 13228 10056
rect 13820 10081 13829 10115
rect 13829 10081 13863 10115
rect 13863 10081 13872 10115
rect 13820 10072 13872 10081
rect 16856 10072 16908 10124
rect 17224 10115 17276 10124
rect 17224 10081 17233 10115
rect 17233 10081 17267 10115
rect 17267 10081 17276 10115
rect 17224 10072 17276 10081
rect 18788 10115 18840 10124
rect 18788 10081 18797 10115
rect 18797 10081 18831 10115
rect 18831 10081 18840 10115
rect 18788 10072 18840 10081
rect 20168 10140 20220 10192
rect 22928 10183 22980 10192
rect 22928 10149 22937 10183
rect 22937 10149 22971 10183
rect 22971 10149 22980 10183
rect 22928 10140 22980 10149
rect 24216 10140 24268 10192
rect 24952 10140 25004 10192
rect 20444 10072 20496 10124
rect 22284 10072 22336 10124
rect 23664 10072 23716 10124
rect 24584 10115 24636 10124
rect 24584 10081 24593 10115
rect 24593 10081 24627 10115
rect 24627 10081 24636 10115
rect 24584 10072 24636 10081
rect 24768 10072 24820 10124
rect 15936 10047 15988 10056
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 17408 10047 17460 10056
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 18972 10047 19024 10056
rect 17408 10004 17460 10013
rect 18972 10013 18981 10047
rect 18981 10013 19015 10047
rect 19015 10013 19024 10047
rect 18972 10004 19024 10013
rect 19064 10004 19116 10056
rect 20628 10004 20680 10056
rect 21456 10004 21508 10056
rect 22652 10004 22704 10056
rect 23296 10047 23348 10056
rect 23296 10013 23305 10047
rect 23305 10013 23339 10047
rect 23339 10013 23348 10047
rect 23296 10004 23348 10013
rect 2596 9868 2648 9920
rect 4068 9911 4120 9920
rect 4068 9877 4077 9911
rect 4077 9877 4111 9911
rect 4111 9877 4120 9911
rect 4068 9868 4120 9877
rect 7288 9868 7340 9920
rect 7564 9868 7616 9920
rect 8208 9868 8260 9920
rect 9496 9936 9548 9988
rect 11336 9979 11388 9988
rect 11336 9945 11345 9979
rect 11345 9945 11379 9979
rect 11379 9945 11388 9979
rect 11336 9936 11388 9945
rect 14188 9936 14240 9988
rect 18880 9936 18932 9988
rect 21640 9936 21692 9988
rect 23204 9936 23256 9988
rect 9588 9868 9640 9920
rect 10324 9868 10376 9920
rect 12256 9868 12308 9920
rect 16856 9911 16908 9920
rect 16856 9877 16865 9911
rect 16865 9877 16899 9911
rect 16899 9877 16908 9911
rect 16856 9868 16908 9877
rect 17960 9868 18012 9920
rect 18236 9868 18288 9920
rect 18420 9911 18472 9920
rect 18420 9877 18429 9911
rect 18429 9877 18463 9911
rect 18463 9877 18472 9911
rect 18420 9868 18472 9877
rect 24032 9911 24084 9920
rect 24032 9877 24041 9911
rect 24041 9877 24075 9911
rect 24075 9877 24084 9911
rect 24032 9868 24084 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2872 9707 2924 9716
rect 2872 9673 2881 9707
rect 2881 9673 2915 9707
rect 2915 9673 2924 9707
rect 2872 9664 2924 9673
rect 1768 9639 1820 9648
rect 1768 9605 1777 9639
rect 1777 9605 1811 9639
rect 1811 9605 1820 9639
rect 1768 9596 1820 9605
rect 2780 9528 2832 9580
rect 3056 9664 3108 9716
rect 5080 9664 5132 9716
rect 6276 9664 6328 9716
rect 6460 9707 6512 9716
rect 6460 9673 6469 9707
rect 6469 9673 6503 9707
rect 6503 9673 6512 9707
rect 6460 9664 6512 9673
rect 9496 9664 9548 9716
rect 10876 9664 10928 9716
rect 4344 9528 4396 9580
rect 8392 9596 8444 9648
rect 11060 9664 11112 9716
rect 12532 9664 12584 9716
rect 12716 9664 12768 9716
rect 14188 9664 14240 9716
rect 17776 9707 17828 9716
rect 11336 9596 11388 9648
rect 11520 9639 11572 9648
rect 11520 9605 11529 9639
rect 11529 9605 11563 9639
rect 11563 9605 11572 9639
rect 11520 9596 11572 9605
rect 12900 9639 12952 9648
rect 12900 9605 12909 9639
rect 12909 9605 12943 9639
rect 12943 9605 12952 9639
rect 12900 9596 12952 9605
rect 14556 9596 14608 9648
rect 16028 9596 16080 9648
rect 17776 9673 17785 9707
rect 17785 9673 17819 9707
rect 17819 9673 17828 9707
rect 17776 9664 17828 9673
rect 19064 9707 19116 9716
rect 19064 9673 19073 9707
rect 19073 9673 19107 9707
rect 19107 9673 19116 9707
rect 19064 9664 19116 9673
rect 20444 9664 20496 9716
rect 20628 9664 20680 9716
rect 22284 9707 22336 9716
rect 22284 9673 22293 9707
rect 22293 9673 22327 9707
rect 22327 9673 22336 9707
rect 22284 9664 22336 9673
rect 22652 9707 22704 9716
rect 22652 9673 22661 9707
rect 22661 9673 22695 9707
rect 22695 9673 22704 9707
rect 22652 9664 22704 9673
rect 23664 9664 23716 9716
rect 23848 9707 23900 9716
rect 23848 9673 23857 9707
rect 23857 9673 23891 9707
rect 23891 9673 23900 9707
rect 23848 9664 23900 9673
rect 24768 9664 24820 9716
rect 20536 9596 20588 9648
rect 22928 9639 22980 9648
rect 22928 9605 22937 9639
rect 22937 9605 22971 9639
rect 22971 9605 22980 9639
rect 22928 9596 22980 9605
rect 6736 9528 6788 9580
rect 7012 9528 7064 9580
rect 7932 9528 7984 9580
rect 8208 9571 8260 9580
rect 8208 9537 8217 9571
rect 8217 9537 8251 9571
rect 8251 9537 8260 9571
rect 8208 9528 8260 9537
rect 2688 9460 2740 9512
rect 8024 9503 8076 9512
rect 8024 9469 8033 9503
rect 8033 9469 8067 9503
rect 8067 9469 8076 9503
rect 8024 9460 8076 9469
rect 8944 9460 8996 9512
rect 9036 9460 9088 9512
rect 9496 9503 9548 9512
rect 9496 9469 9530 9503
rect 9530 9469 9548 9503
rect 9496 9460 9548 9469
rect 2136 9435 2188 9444
rect 2136 9401 2145 9435
rect 2145 9401 2179 9435
rect 2179 9401 2188 9435
rect 2136 9392 2188 9401
rect 3148 9392 3200 9444
rect 4252 9392 4304 9444
rect 6736 9392 6788 9444
rect 7748 9392 7800 9444
rect 9404 9392 9456 9444
rect 9680 9392 9732 9444
rect 10324 9392 10376 9444
rect 11060 9392 11112 9444
rect 1584 9324 1636 9376
rect 5908 9324 5960 9376
rect 6368 9324 6420 9376
rect 7380 9324 7432 9376
rect 7656 9367 7708 9376
rect 7656 9333 7665 9367
rect 7665 9333 7699 9367
rect 7699 9333 7708 9367
rect 7656 9324 7708 9333
rect 9036 9367 9088 9376
rect 9036 9333 9045 9367
rect 9045 9333 9079 9367
rect 9079 9333 9088 9367
rect 9036 9324 9088 9333
rect 12440 9367 12492 9376
rect 12440 9333 12449 9367
rect 12449 9333 12483 9367
rect 12483 9333 12492 9367
rect 12440 9324 12492 9333
rect 12992 9324 13044 9376
rect 15108 9528 15160 9580
rect 15936 9528 15988 9580
rect 18604 9571 18656 9580
rect 18604 9537 18613 9571
rect 18613 9537 18647 9571
rect 18647 9537 18656 9571
rect 18604 9528 18656 9537
rect 18972 9528 19024 9580
rect 20260 9571 20312 9580
rect 20260 9537 20269 9571
rect 20269 9537 20303 9571
rect 20303 9537 20312 9571
rect 20260 9528 20312 9537
rect 20628 9528 20680 9580
rect 21180 9528 21232 9580
rect 21364 9528 21416 9580
rect 21916 9528 21968 9580
rect 23848 9528 23900 9580
rect 16396 9503 16448 9512
rect 16396 9469 16405 9503
rect 16405 9469 16439 9503
rect 16439 9469 16448 9503
rect 16396 9460 16448 9469
rect 17776 9460 17828 9512
rect 20536 9460 20588 9512
rect 20812 9460 20864 9512
rect 21640 9503 21692 9512
rect 21640 9469 21649 9503
rect 21649 9469 21683 9503
rect 21683 9469 21692 9503
rect 21640 9460 21692 9469
rect 23664 9503 23716 9512
rect 15752 9392 15804 9444
rect 17960 9392 18012 9444
rect 21548 9435 21600 9444
rect 13452 9324 13504 9376
rect 14648 9324 14700 9376
rect 16120 9324 16172 9376
rect 16304 9367 16356 9376
rect 16304 9333 16313 9367
rect 16313 9333 16347 9367
rect 16347 9333 16356 9367
rect 16304 9324 16356 9333
rect 17224 9324 17276 9376
rect 18328 9324 18380 9376
rect 18972 9324 19024 9376
rect 20812 9324 20864 9376
rect 21548 9401 21557 9435
rect 21557 9401 21591 9435
rect 21591 9401 21600 9435
rect 23664 9469 23673 9503
rect 23673 9469 23707 9503
rect 23707 9469 23716 9503
rect 23664 9460 23716 9469
rect 24860 9460 24912 9512
rect 21548 9392 21600 9401
rect 24308 9392 24360 9444
rect 23020 9324 23072 9376
rect 23388 9324 23440 9376
rect 26056 9367 26108 9376
rect 26056 9333 26065 9367
rect 26065 9333 26099 9367
rect 26099 9333 26108 9367
rect 26056 9324 26108 9333
rect 26424 9367 26476 9376
rect 26424 9333 26433 9367
rect 26433 9333 26467 9367
rect 26467 9333 26476 9367
rect 26424 9324 26476 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2412 9163 2464 9172
rect 2412 9129 2421 9163
rect 2421 9129 2455 9163
rect 2455 9129 2464 9163
rect 2412 9120 2464 9129
rect 4712 9120 4764 9172
rect 4896 9163 4948 9172
rect 4896 9129 4905 9163
rect 4905 9129 4939 9163
rect 4939 9129 4948 9163
rect 4896 9120 4948 9129
rect 7748 9120 7800 9172
rect 7932 9120 7984 9172
rect 8944 9120 8996 9172
rect 9496 9120 9548 9172
rect 9772 9120 9824 9172
rect 10140 9120 10192 9172
rect 10968 9120 11020 9172
rect 13176 9163 13228 9172
rect 13176 9129 13185 9163
rect 13185 9129 13219 9163
rect 13219 9129 13228 9163
rect 13176 9120 13228 9129
rect 13728 9120 13780 9172
rect 14004 9163 14056 9172
rect 14004 9129 14013 9163
rect 14013 9129 14047 9163
rect 14047 9129 14056 9163
rect 14004 9120 14056 9129
rect 4804 9095 4856 9104
rect 4804 9061 4813 9095
rect 4813 9061 4847 9095
rect 4847 9061 4856 9095
rect 4804 9052 4856 9061
rect 5816 9095 5868 9104
rect 5816 9061 5825 9095
rect 5825 9061 5859 9095
rect 5859 9061 5868 9095
rect 5816 9052 5868 9061
rect 2228 8984 2280 9036
rect 4252 8984 4304 9036
rect 7012 9052 7064 9104
rect 8576 9052 8628 9104
rect 11796 9052 11848 9104
rect 13360 9052 13412 9104
rect 14924 9120 14976 9172
rect 15108 9163 15160 9172
rect 15108 9129 15117 9163
rect 15117 9129 15151 9163
rect 15151 9129 15160 9163
rect 15108 9120 15160 9129
rect 17408 9120 17460 9172
rect 18788 9163 18840 9172
rect 18788 9129 18797 9163
rect 18797 9129 18831 9163
rect 18831 9129 18840 9163
rect 18788 9120 18840 9129
rect 20260 9163 20312 9172
rect 20260 9129 20269 9163
rect 20269 9129 20303 9163
rect 20303 9129 20312 9163
rect 20260 9120 20312 9129
rect 20720 9163 20772 9172
rect 20720 9129 20729 9163
rect 20729 9129 20763 9163
rect 20763 9129 20772 9163
rect 20720 9120 20772 9129
rect 20904 9120 20956 9172
rect 21916 9163 21968 9172
rect 15292 9052 15344 9104
rect 15844 9052 15896 9104
rect 19432 9052 19484 9104
rect 21364 9052 21416 9104
rect 21916 9129 21925 9163
rect 21925 9129 21959 9163
rect 21959 9129 21968 9163
rect 21916 9120 21968 9129
rect 23296 9163 23348 9172
rect 23296 9129 23305 9163
rect 23305 9129 23339 9163
rect 23339 9129 23348 9163
rect 23296 9120 23348 9129
rect 23480 9120 23532 9172
rect 24308 9163 24360 9172
rect 24308 9129 24317 9163
rect 24317 9129 24351 9163
rect 24351 9129 24360 9163
rect 24308 9120 24360 9129
rect 25044 9163 25096 9172
rect 25044 9129 25053 9163
rect 25053 9129 25087 9163
rect 25087 9129 25096 9163
rect 25044 9120 25096 9129
rect 25412 9163 25464 9172
rect 25412 9129 25421 9163
rect 25421 9129 25455 9163
rect 25455 9129 25464 9163
rect 25412 9120 25464 9129
rect 25780 9163 25832 9172
rect 25780 9129 25789 9163
rect 25789 9129 25823 9163
rect 25823 9129 25832 9163
rect 25780 9120 25832 9129
rect 26240 9163 26292 9172
rect 26240 9129 26249 9163
rect 26249 9129 26283 9163
rect 26283 9129 26292 9163
rect 26240 9120 26292 9129
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 3148 8916 3200 8968
rect 3700 8916 3752 8968
rect 5448 8916 5500 8968
rect 6368 8984 6420 9036
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 11980 8984 12032 9036
rect 17960 8984 18012 9036
rect 18052 8984 18104 9036
rect 20168 8984 20220 9036
rect 20812 8984 20864 9036
rect 21732 8984 21784 9036
rect 9036 8916 9088 8968
rect 9772 8916 9824 8968
rect 14188 8959 14240 8968
rect 14188 8925 14197 8959
rect 14197 8925 14231 8959
rect 14231 8925 14240 8959
rect 14188 8916 14240 8925
rect 14740 8916 14792 8968
rect 13544 8848 13596 8900
rect 5172 8780 5224 8832
rect 5540 8823 5592 8832
rect 5540 8789 5549 8823
rect 5549 8789 5583 8823
rect 5583 8789 5592 8823
rect 5540 8780 5592 8789
rect 6460 8780 6512 8832
rect 7932 8780 7984 8832
rect 12164 8780 12216 8832
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 14740 8823 14792 8832
rect 14740 8789 14749 8823
rect 14749 8789 14783 8823
rect 14783 8789 14792 8823
rect 14740 8780 14792 8789
rect 16304 8916 16356 8968
rect 17224 8916 17276 8968
rect 18236 8959 18288 8968
rect 18236 8925 18245 8959
rect 18245 8925 18279 8959
rect 18279 8925 18288 8959
rect 18236 8916 18288 8925
rect 16580 8848 16632 8900
rect 18604 8916 18656 8968
rect 19984 8916 20036 8968
rect 20628 8916 20680 8968
rect 21364 8959 21416 8968
rect 21364 8925 21373 8959
rect 21373 8925 21407 8959
rect 21407 8925 21416 8959
rect 21364 8916 21416 8925
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 21456 8916 21508 8925
rect 19616 8891 19668 8900
rect 15568 8780 15620 8832
rect 17224 8780 17276 8832
rect 17408 8780 17460 8832
rect 19616 8857 19625 8891
rect 19625 8857 19659 8891
rect 19659 8857 19668 8891
rect 19616 8848 19668 8857
rect 20996 8848 21048 8900
rect 21916 8848 21968 8900
rect 22100 8984 22152 9036
rect 23020 8984 23072 9036
rect 23940 8984 23992 9036
rect 26056 8916 26108 8968
rect 23572 8848 23624 8900
rect 20628 8780 20680 8832
rect 20904 8823 20956 8832
rect 20904 8789 20913 8823
rect 20913 8789 20947 8823
rect 20947 8789 20956 8823
rect 20904 8780 20956 8789
rect 21364 8780 21416 8832
rect 22284 8823 22336 8832
rect 22284 8789 22293 8823
rect 22293 8789 22327 8823
rect 22327 8789 22336 8823
rect 22284 8780 22336 8789
rect 22652 8823 22704 8832
rect 22652 8789 22661 8823
rect 22661 8789 22695 8823
rect 22695 8789 22704 8823
rect 22652 8780 22704 8789
rect 22928 8823 22980 8832
rect 22928 8789 22937 8823
rect 22937 8789 22971 8823
rect 22971 8789 22980 8823
rect 22928 8780 22980 8789
rect 23664 8823 23716 8832
rect 23664 8789 23673 8823
rect 23673 8789 23707 8823
rect 23707 8789 23716 8823
rect 23664 8780 23716 8789
rect 23940 8823 23992 8832
rect 23940 8789 23949 8823
rect 23949 8789 23983 8823
rect 23983 8789 23992 8823
rect 23940 8780 23992 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2044 8576 2096 8628
rect 2320 8576 2372 8628
rect 4896 8576 4948 8628
rect 2872 8508 2924 8560
rect 1768 8440 1820 8492
rect 3700 8483 3752 8492
rect 1860 8415 1912 8424
rect 1860 8381 1869 8415
rect 1869 8381 1903 8415
rect 1903 8381 1912 8415
rect 1860 8372 1912 8381
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 3332 8372 3384 8424
rect 2964 8236 3016 8288
rect 3700 8304 3752 8356
rect 5264 8508 5316 8560
rect 4804 8440 4856 8492
rect 5448 8440 5500 8492
rect 9496 8576 9548 8628
rect 10048 8576 10100 8628
rect 12072 8619 12124 8628
rect 12072 8585 12081 8619
rect 12081 8585 12115 8619
rect 12115 8585 12124 8619
rect 12072 8576 12124 8585
rect 14464 8576 14516 8628
rect 15752 8619 15804 8628
rect 15752 8585 15761 8619
rect 15761 8585 15795 8619
rect 15795 8585 15804 8619
rect 15752 8576 15804 8585
rect 20168 8576 20220 8628
rect 20536 8619 20588 8628
rect 20536 8585 20545 8619
rect 20545 8585 20579 8619
rect 20579 8585 20588 8619
rect 20536 8576 20588 8585
rect 21456 8576 21508 8628
rect 7012 8440 7064 8492
rect 10048 8440 10100 8492
rect 10600 8440 10652 8492
rect 16028 8508 16080 8560
rect 4712 8372 4764 8424
rect 6184 8372 6236 8424
rect 5632 8304 5684 8356
rect 3884 8236 3936 8288
rect 4988 8236 5040 8288
rect 6184 8236 6236 8288
rect 9036 8372 9088 8424
rect 10968 8440 11020 8492
rect 12992 8440 13044 8492
rect 16212 8483 16264 8492
rect 16212 8449 16221 8483
rect 16221 8449 16255 8483
rect 16255 8449 16264 8483
rect 16212 8440 16264 8449
rect 19064 8508 19116 8560
rect 20996 8483 21048 8492
rect 20996 8449 21005 8483
rect 21005 8449 21039 8483
rect 21039 8449 21048 8483
rect 20996 8440 21048 8449
rect 7932 8304 7984 8356
rect 10784 8304 10836 8356
rect 15844 8372 15896 8424
rect 16672 8372 16724 8424
rect 13636 8304 13688 8356
rect 7012 8279 7064 8288
rect 7012 8245 7021 8279
rect 7021 8245 7055 8279
rect 7055 8245 7064 8279
rect 7012 8236 7064 8245
rect 9772 8236 9824 8288
rect 11520 8236 11572 8288
rect 11796 8236 11848 8288
rect 12440 8236 12492 8288
rect 15476 8304 15528 8356
rect 15292 8236 15344 8288
rect 15568 8236 15620 8288
rect 20720 8372 20772 8424
rect 20444 8304 20496 8356
rect 21732 8372 21784 8424
rect 22836 8576 22888 8628
rect 23020 8619 23072 8628
rect 23020 8585 23029 8619
rect 23029 8585 23063 8619
rect 23063 8585 23072 8619
rect 23020 8576 23072 8585
rect 23480 8619 23532 8628
rect 23480 8585 23489 8619
rect 23489 8585 23523 8619
rect 23523 8585 23532 8619
rect 23480 8576 23532 8585
rect 24032 8576 24084 8628
rect 25136 8576 25188 8628
rect 25688 8619 25740 8628
rect 25688 8585 25697 8619
rect 25697 8585 25731 8619
rect 25731 8585 25740 8619
rect 25688 8576 25740 8585
rect 25964 8619 26016 8628
rect 25964 8585 25973 8619
rect 25973 8585 26007 8619
rect 26007 8585 26016 8619
rect 25964 8576 26016 8585
rect 26332 8619 26384 8628
rect 26332 8585 26341 8619
rect 26341 8585 26375 8619
rect 26375 8585 26384 8619
rect 26332 8576 26384 8585
rect 23204 8508 23256 8560
rect 26148 8508 26200 8560
rect 22192 8440 22244 8492
rect 23480 8440 23532 8492
rect 23664 8415 23716 8424
rect 23664 8381 23673 8415
rect 23673 8381 23707 8415
rect 23707 8381 23716 8415
rect 23664 8372 23716 8381
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 21272 8236 21324 8288
rect 21640 8236 21692 8288
rect 22744 8236 22796 8288
rect 23848 8279 23900 8288
rect 23848 8245 23857 8279
rect 23857 8245 23891 8279
rect 23891 8245 23900 8279
rect 23848 8236 23900 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2228 8075 2280 8084
rect 2228 8041 2237 8075
rect 2237 8041 2271 8075
rect 2271 8041 2280 8075
rect 2228 8032 2280 8041
rect 2412 8032 2464 8084
rect 4160 8032 4212 8084
rect 4712 8075 4764 8084
rect 4712 8041 4721 8075
rect 4721 8041 4755 8075
rect 4755 8041 4764 8075
rect 4712 8032 4764 8041
rect 4988 8032 5040 8084
rect 8668 8032 8720 8084
rect 10692 8032 10744 8084
rect 11152 8032 11204 8084
rect 12348 8032 12400 8084
rect 14188 8032 14240 8084
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 18236 8032 18288 8084
rect 20996 8032 21048 8084
rect 22836 8032 22888 8084
rect 24124 8032 24176 8084
rect 25044 8075 25096 8084
rect 25044 8041 25053 8075
rect 25053 8041 25087 8075
rect 25087 8041 25096 8075
rect 25044 8032 25096 8041
rect 2964 7964 3016 8016
rect 6092 7964 6144 8016
rect 8576 7964 8628 8016
rect 10784 7964 10836 8016
rect 10968 7964 11020 8016
rect 14648 7964 14700 8016
rect 16120 7964 16172 8016
rect 3608 7896 3660 7948
rect 6184 7896 6236 7948
rect 8392 7939 8444 7948
rect 8392 7905 8401 7939
rect 8401 7905 8435 7939
rect 8435 7905 8444 7939
rect 8392 7896 8444 7905
rect 3056 7828 3108 7880
rect 3700 7828 3752 7880
rect 7932 7828 7984 7880
rect 8208 7828 8260 7880
rect 9772 7828 9824 7880
rect 10876 7828 10928 7880
rect 12164 7896 12216 7948
rect 15292 7871 15344 7880
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 3884 7735 3936 7744
rect 3884 7701 3893 7735
rect 3893 7701 3927 7735
rect 3927 7701 3936 7735
rect 3884 7692 3936 7701
rect 4620 7692 4672 7744
rect 5540 7692 5592 7744
rect 6368 7692 6420 7744
rect 7012 7692 7064 7744
rect 8024 7735 8076 7744
rect 8024 7701 8033 7735
rect 8033 7701 8067 7735
rect 8067 7701 8076 7735
rect 8024 7692 8076 7701
rect 9588 7692 9640 7744
rect 11520 7692 11572 7744
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 18236 7871 18288 7880
rect 18236 7837 18245 7871
rect 18245 7837 18279 7871
rect 18279 7837 18288 7871
rect 18236 7828 18288 7837
rect 18512 7964 18564 8016
rect 21916 7964 21968 8016
rect 19340 7939 19392 7948
rect 19340 7905 19349 7939
rect 19349 7905 19383 7939
rect 19383 7905 19392 7939
rect 19340 7896 19392 7905
rect 22376 7896 22428 7948
rect 22744 7896 22796 7948
rect 23480 7896 23532 7948
rect 24032 7939 24084 7948
rect 24032 7905 24041 7939
rect 24041 7905 24075 7939
rect 24075 7905 24084 7939
rect 24032 7896 24084 7905
rect 25228 7896 25280 7948
rect 18604 7828 18656 7880
rect 19248 7828 19300 7880
rect 18512 7760 18564 7812
rect 19892 7803 19944 7812
rect 19892 7769 19901 7803
rect 19901 7769 19935 7803
rect 19935 7769 19944 7803
rect 19892 7760 19944 7769
rect 12992 7692 13044 7744
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 14464 7735 14516 7744
rect 14464 7701 14473 7735
rect 14473 7701 14507 7735
rect 14507 7701 14516 7735
rect 14464 7692 14516 7701
rect 16028 7692 16080 7744
rect 17408 7692 17460 7744
rect 18236 7692 18288 7744
rect 20444 7760 20496 7812
rect 21732 7828 21784 7880
rect 23020 7871 23072 7880
rect 23020 7837 23029 7871
rect 23029 7837 23063 7871
rect 23063 7837 23072 7871
rect 23020 7828 23072 7837
rect 26056 7871 26108 7880
rect 26056 7837 26065 7871
rect 26065 7837 26099 7871
rect 26099 7837 26108 7871
rect 26056 7828 26108 7837
rect 23388 7760 23440 7812
rect 21548 7692 21600 7744
rect 21916 7735 21968 7744
rect 21916 7701 21925 7735
rect 21925 7701 21959 7735
rect 21959 7701 21968 7735
rect 21916 7692 21968 7701
rect 22376 7735 22428 7744
rect 22376 7701 22385 7735
rect 22385 7701 22419 7735
rect 22419 7701 22428 7735
rect 22376 7692 22428 7701
rect 23480 7735 23532 7744
rect 23480 7701 23489 7735
rect 23489 7701 23523 7735
rect 23523 7701 23532 7735
rect 23480 7692 23532 7701
rect 23572 7692 23624 7744
rect 25136 7692 25188 7744
rect 25320 7735 25372 7744
rect 25320 7701 25329 7735
rect 25329 7701 25363 7735
rect 25363 7701 25372 7735
rect 25320 7692 25372 7701
rect 25688 7735 25740 7744
rect 25688 7701 25697 7735
rect 25697 7701 25731 7735
rect 25731 7701 25740 7735
rect 25688 7692 25740 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 3148 7531 3200 7540
rect 3148 7497 3157 7531
rect 3157 7497 3191 7531
rect 3191 7497 3200 7531
rect 3148 7488 3200 7497
rect 6092 7531 6144 7540
rect 6092 7497 6101 7531
rect 6101 7497 6135 7531
rect 6135 7497 6144 7531
rect 6092 7488 6144 7497
rect 8208 7531 8260 7540
rect 8208 7497 8217 7531
rect 8217 7497 8251 7531
rect 8251 7497 8260 7531
rect 8208 7488 8260 7497
rect 8392 7488 8444 7540
rect 10876 7488 10928 7540
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 18052 7531 18104 7540
rect 18052 7497 18061 7531
rect 18061 7497 18095 7531
rect 18095 7497 18104 7531
rect 18052 7488 18104 7497
rect 19340 7531 19392 7540
rect 19340 7497 19349 7531
rect 19349 7497 19383 7531
rect 19383 7497 19392 7531
rect 19340 7488 19392 7497
rect 20812 7488 20864 7540
rect 21180 7531 21232 7540
rect 21180 7497 21189 7531
rect 21189 7497 21223 7531
rect 21223 7497 21232 7531
rect 21180 7488 21232 7497
rect 22928 7531 22980 7540
rect 22928 7497 22937 7531
rect 22937 7497 22971 7531
rect 22971 7497 22980 7531
rect 22928 7488 22980 7497
rect 24032 7488 24084 7540
rect 25228 7488 25280 7540
rect 25504 7488 25556 7540
rect 3056 7463 3108 7472
rect 3056 7429 3065 7463
rect 3065 7429 3099 7463
rect 3099 7429 3108 7463
rect 3056 7420 3108 7429
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 7104 7463 7156 7472
rect 2228 7352 2280 7361
rect 1952 7327 2004 7336
rect 1952 7293 1961 7327
rect 1961 7293 1995 7327
rect 1995 7293 2004 7327
rect 1952 7284 2004 7293
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 7104 7429 7113 7463
rect 7113 7429 7147 7463
rect 7147 7429 7156 7463
rect 7104 7420 7156 7429
rect 8576 7463 8628 7472
rect 8576 7429 8585 7463
rect 8585 7429 8619 7463
rect 8619 7429 8628 7463
rect 8576 7420 8628 7429
rect 12440 7463 12492 7472
rect 12440 7429 12449 7463
rect 12449 7429 12483 7463
rect 12483 7429 12492 7463
rect 12440 7420 12492 7429
rect 17592 7420 17644 7472
rect 18512 7420 18564 7472
rect 7932 7352 7984 7404
rect 9772 7395 9824 7404
rect 9772 7361 9781 7395
rect 9781 7361 9815 7395
rect 9815 7361 9824 7395
rect 9772 7352 9824 7361
rect 11796 7352 11848 7404
rect 13544 7352 13596 7404
rect 14004 7352 14056 7404
rect 16120 7395 16172 7404
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 19892 7352 19944 7404
rect 20260 7352 20312 7404
rect 20720 7420 20772 7472
rect 20904 7352 20956 7404
rect 21640 7395 21692 7404
rect 21640 7361 21649 7395
rect 21649 7361 21683 7395
rect 21683 7361 21692 7395
rect 21640 7352 21692 7361
rect 22560 7352 22612 7404
rect 3792 7284 3844 7336
rect 5540 7284 5592 7336
rect 6184 7284 6236 7336
rect 7564 7327 7616 7336
rect 7564 7293 7573 7327
rect 7573 7293 7607 7327
rect 7607 7293 7616 7327
rect 7564 7284 7616 7293
rect 11152 7327 11204 7336
rect 11152 7293 11161 7327
rect 11161 7293 11195 7327
rect 11195 7293 11204 7327
rect 11152 7284 11204 7293
rect 13820 7284 13872 7336
rect 14464 7327 14516 7336
rect 14464 7293 14473 7327
rect 14473 7293 14507 7327
rect 14507 7293 14516 7327
rect 14464 7284 14516 7293
rect 15660 7284 15712 7336
rect 19984 7284 20036 7336
rect 21548 7327 21600 7336
rect 21548 7293 21557 7327
rect 21557 7293 21591 7327
rect 21591 7293 21600 7327
rect 21548 7284 21600 7293
rect 23848 7284 23900 7336
rect 24768 7327 24820 7336
rect 24768 7293 24777 7327
rect 24777 7293 24811 7327
rect 24811 7293 24820 7327
rect 24768 7284 24820 7293
rect 5264 7216 5316 7268
rect 7380 7216 7432 7268
rect 9588 7259 9640 7268
rect 9588 7225 9597 7259
rect 9597 7225 9631 7259
rect 9631 7225 9640 7259
rect 9588 7216 9640 7225
rect 10968 7216 11020 7268
rect 11060 7216 11112 7268
rect 15752 7216 15804 7268
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 2780 7148 2832 7200
rect 3516 7191 3568 7200
rect 3516 7157 3525 7191
rect 3525 7157 3559 7191
rect 3559 7157 3568 7191
rect 3516 7148 3568 7157
rect 4160 7191 4212 7200
rect 4160 7157 4169 7191
rect 4169 7157 4203 7191
rect 4203 7157 4212 7191
rect 4160 7148 4212 7157
rect 4712 7191 4764 7200
rect 4712 7157 4721 7191
rect 4721 7157 4755 7191
rect 4755 7157 4764 7191
rect 4712 7148 4764 7157
rect 7564 7148 7616 7200
rect 7748 7148 7800 7200
rect 9220 7191 9272 7200
rect 9220 7157 9229 7191
rect 9229 7157 9263 7191
rect 9263 7157 9272 7191
rect 9220 7148 9272 7157
rect 9680 7191 9732 7200
rect 9680 7157 9689 7191
rect 9689 7157 9723 7191
rect 9723 7157 9732 7191
rect 9680 7148 9732 7157
rect 11336 7148 11388 7200
rect 12532 7148 12584 7200
rect 12992 7148 13044 7200
rect 13544 7148 13596 7200
rect 13912 7148 13964 7200
rect 14280 7148 14332 7200
rect 15568 7191 15620 7200
rect 15568 7157 15577 7191
rect 15577 7157 15611 7191
rect 15611 7157 15620 7191
rect 15568 7148 15620 7157
rect 18420 7191 18472 7200
rect 18420 7157 18429 7191
rect 18429 7157 18463 7191
rect 18463 7157 18472 7191
rect 18420 7148 18472 7157
rect 19340 7216 19392 7268
rect 20168 7216 20220 7268
rect 22744 7216 22796 7268
rect 23940 7216 23992 7268
rect 18788 7148 18840 7200
rect 19432 7148 19484 7200
rect 20812 7148 20864 7200
rect 21732 7148 21784 7200
rect 22008 7148 22060 7200
rect 22100 7148 22152 7200
rect 23020 7148 23072 7200
rect 23296 7191 23348 7200
rect 23296 7157 23305 7191
rect 23305 7157 23339 7191
rect 23339 7157 23348 7191
rect 23296 7148 23348 7157
rect 24124 7148 24176 7200
rect 25964 7148 26016 7200
rect 26148 7191 26200 7200
rect 26148 7157 26157 7191
rect 26157 7157 26191 7191
rect 26191 7157 26200 7191
rect 26148 7148 26200 7157
rect 26424 7191 26476 7200
rect 26424 7157 26433 7191
rect 26433 7157 26467 7191
rect 26467 7157 26476 7191
rect 26424 7148 26476 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1952 6944 2004 6996
rect 4068 6987 4120 6996
rect 4068 6953 4077 6987
rect 4077 6953 4111 6987
rect 4111 6953 4120 6987
rect 4068 6944 4120 6953
rect 4436 6987 4488 6996
rect 4436 6953 4445 6987
rect 4445 6953 4479 6987
rect 4479 6953 4488 6987
rect 4436 6944 4488 6953
rect 6276 6944 6328 6996
rect 7104 6944 7156 6996
rect 9772 6944 9824 6996
rect 11796 6987 11848 6996
rect 11796 6953 11805 6987
rect 11805 6953 11839 6987
rect 11839 6953 11848 6987
rect 11796 6944 11848 6953
rect 12532 6987 12584 6996
rect 12532 6953 12541 6987
rect 12541 6953 12575 6987
rect 12575 6953 12584 6987
rect 12532 6944 12584 6953
rect 14004 6987 14056 6996
rect 14004 6953 14013 6987
rect 14013 6953 14047 6987
rect 14047 6953 14056 6987
rect 14004 6944 14056 6953
rect 18696 6944 18748 6996
rect 19340 6944 19392 6996
rect 21272 6987 21324 6996
rect 21272 6953 21281 6987
rect 21281 6953 21315 6987
rect 21315 6953 21324 6987
rect 21272 6944 21324 6953
rect 22376 6944 22428 6996
rect 22836 6987 22888 6996
rect 22836 6953 22845 6987
rect 22845 6953 22879 6987
rect 22879 6953 22888 6987
rect 22836 6944 22888 6953
rect 2320 6876 2372 6928
rect 3148 6876 3200 6928
rect 3700 6876 3752 6928
rect 6184 6876 6236 6928
rect 4712 6808 4764 6860
rect 6276 6808 6328 6860
rect 10416 6876 10468 6928
rect 11612 6876 11664 6928
rect 13268 6919 13320 6928
rect 13268 6885 13277 6919
rect 13277 6885 13311 6919
rect 13311 6885 13320 6919
rect 13268 6876 13320 6885
rect 18604 6876 18656 6928
rect 18972 6876 19024 6928
rect 3240 6740 3292 6792
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 5264 6783 5316 6792
rect 5264 6749 5273 6783
rect 5273 6749 5307 6783
rect 5307 6749 5316 6783
rect 5264 6740 5316 6749
rect 6000 6740 6052 6792
rect 7748 6808 7800 6860
rect 8116 6851 8168 6860
rect 8116 6817 8125 6851
rect 8125 6817 8159 6851
rect 8159 6817 8168 6851
rect 8116 6808 8168 6817
rect 8208 6851 8260 6860
rect 8208 6817 8217 6851
rect 8217 6817 8251 6851
rect 8251 6817 8260 6851
rect 8208 6808 8260 6817
rect 11152 6808 11204 6860
rect 8668 6740 8720 6792
rect 9036 6740 9088 6792
rect 9220 6740 9272 6792
rect 2412 6715 2464 6724
rect 2412 6681 2421 6715
rect 2421 6681 2455 6715
rect 2455 6681 2464 6715
rect 2412 6672 2464 6681
rect 3056 6672 3108 6724
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 2780 6604 2832 6656
rect 3700 6604 3752 6656
rect 6092 6715 6144 6724
rect 6092 6681 6101 6715
rect 6101 6681 6135 6715
rect 6135 6681 6144 6715
rect 6092 6672 6144 6681
rect 8944 6672 8996 6724
rect 9496 6672 9548 6724
rect 4896 6604 4948 6656
rect 6552 6604 6604 6656
rect 7380 6604 7432 6656
rect 9772 6604 9824 6656
rect 9956 6604 10008 6656
rect 10140 6604 10192 6656
rect 11796 6672 11848 6724
rect 12716 6672 12768 6724
rect 14648 6808 14700 6860
rect 15476 6851 15528 6860
rect 15476 6817 15485 6851
rect 15485 6817 15519 6851
rect 15519 6817 15528 6851
rect 15476 6808 15528 6817
rect 16488 6851 16540 6860
rect 16488 6817 16497 6851
rect 16497 6817 16531 6851
rect 16531 6817 16540 6851
rect 16488 6808 16540 6817
rect 16672 6808 16724 6860
rect 17868 6808 17920 6860
rect 17960 6808 18012 6860
rect 19156 6808 19208 6860
rect 23664 6944 23716 6996
rect 24032 6944 24084 6996
rect 24768 6987 24820 6996
rect 24768 6953 24777 6987
rect 24777 6953 24811 6987
rect 24811 6953 24820 6987
rect 24768 6944 24820 6953
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 15292 6740 15344 6792
rect 16120 6740 16172 6792
rect 18236 6740 18288 6792
rect 19616 6740 19668 6792
rect 22376 6808 22428 6860
rect 22744 6808 22796 6860
rect 24032 6851 24084 6860
rect 24032 6817 24041 6851
rect 24041 6817 24075 6851
rect 24075 6817 24084 6851
rect 24032 6808 24084 6817
rect 14740 6672 14792 6724
rect 12532 6604 12584 6656
rect 13728 6604 13780 6656
rect 15660 6647 15712 6656
rect 15660 6613 15669 6647
rect 15669 6613 15703 6647
rect 15703 6613 15712 6647
rect 15660 6604 15712 6613
rect 16120 6647 16172 6656
rect 16120 6613 16129 6647
rect 16129 6613 16163 6647
rect 16163 6613 16172 6647
rect 16120 6604 16172 6613
rect 21180 6740 21232 6792
rect 21364 6783 21416 6792
rect 21364 6749 21373 6783
rect 21373 6749 21407 6783
rect 21407 6749 21416 6783
rect 21364 6740 21416 6749
rect 20904 6715 20956 6724
rect 20904 6681 20913 6715
rect 20913 6681 20947 6715
rect 20947 6681 20956 6715
rect 20904 6672 20956 6681
rect 22560 6740 22612 6792
rect 23296 6740 23348 6792
rect 23756 6740 23808 6792
rect 22008 6672 22060 6724
rect 25228 6740 25280 6792
rect 25780 6672 25832 6724
rect 17960 6647 18012 6656
rect 17960 6613 17969 6647
rect 17969 6613 18003 6647
rect 18003 6613 18012 6647
rect 17960 6604 18012 6613
rect 19064 6647 19116 6656
rect 19064 6613 19073 6647
rect 19073 6613 19107 6647
rect 19107 6613 19116 6647
rect 19064 6604 19116 6613
rect 19340 6604 19392 6656
rect 20168 6647 20220 6656
rect 20168 6613 20177 6647
rect 20177 6613 20211 6647
rect 20211 6613 20220 6647
rect 20168 6604 20220 6613
rect 20996 6604 21048 6656
rect 22284 6647 22336 6656
rect 22284 6613 22293 6647
rect 22293 6613 22327 6647
rect 22327 6613 22336 6647
rect 22284 6604 22336 6613
rect 23756 6647 23808 6656
rect 23756 6613 23765 6647
rect 23765 6613 23799 6647
rect 23799 6613 23808 6647
rect 23756 6604 23808 6613
rect 23848 6604 23900 6656
rect 24860 6604 24912 6656
rect 26056 6647 26108 6656
rect 26056 6613 26065 6647
rect 26065 6613 26099 6647
rect 26099 6613 26108 6647
rect 26056 6604 26108 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2504 6400 2556 6452
rect 3240 6443 3292 6452
rect 3240 6409 3249 6443
rect 3249 6409 3283 6443
rect 3283 6409 3292 6443
rect 3240 6400 3292 6409
rect 6000 6400 6052 6452
rect 7104 6400 7156 6452
rect 8116 6400 8168 6452
rect 9956 6400 10008 6452
rect 10600 6443 10652 6452
rect 6184 6332 6236 6384
rect 2228 6264 2280 6316
rect 2320 6264 2372 6316
rect 6828 6307 6880 6316
rect 2596 6239 2648 6248
rect 2596 6205 2605 6239
rect 2605 6205 2639 6239
rect 2639 6205 2648 6239
rect 2596 6196 2648 6205
rect 3240 6196 3292 6248
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 4068 6239 4120 6248
rect 4068 6205 4102 6239
rect 4102 6205 4120 6239
rect 4068 6196 4120 6205
rect 7748 6196 7800 6248
rect 4252 6128 4304 6180
rect 7380 6128 7432 6180
rect 8300 6128 8352 6180
rect 10600 6409 10609 6443
rect 10609 6409 10643 6443
rect 10643 6409 10652 6443
rect 10600 6400 10652 6409
rect 13268 6400 13320 6452
rect 15568 6400 15620 6452
rect 15936 6400 15988 6452
rect 16856 6400 16908 6452
rect 21088 6400 21140 6452
rect 22560 6443 22612 6452
rect 22560 6409 22569 6443
rect 22569 6409 22603 6443
rect 22603 6409 22612 6443
rect 22560 6400 22612 6409
rect 22836 6443 22888 6452
rect 22836 6409 22845 6443
rect 22845 6409 22879 6443
rect 22879 6409 22888 6443
rect 22836 6400 22888 6409
rect 24032 6400 24084 6452
rect 25044 6443 25096 6452
rect 25044 6409 25053 6443
rect 25053 6409 25087 6443
rect 25087 6409 25096 6443
rect 25044 6400 25096 6409
rect 25780 6443 25832 6452
rect 25780 6409 25789 6443
rect 25789 6409 25823 6443
rect 25823 6409 25832 6443
rect 25780 6400 25832 6409
rect 10508 6375 10560 6384
rect 10508 6341 10517 6375
rect 10517 6341 10551 6375
rect 10551 6341 10560 6375
rect 10508 6332 10560 6341
rect 14556 6332 14608 6384
rect 17868 6375 17920 6384
rect 17868 6341 17877 6375
rect 17877 6341 17911 6375
rect 17911 6341 17920 6375
rect 17868 6332 17920 6341
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 17132 6264 17184 6316
rect 17960 6264 18012 6316
rect 18236 6264 18288 6316
rect 18972 6264 19024 6316
rect 19616 6332 19668 6384
rect 21272 6332 21324 6384
rect 3148 6060 3200 6112
rect 5448 6060 5500 6112
rect 8208 6060 8260 6112
rect 9956 6060 10008 6112
rect 11796 6060 11848 6112
rect 12992 6196 13044 6248
rect 14096 6196 14148 6248
rect 16856 6239 16908 6248
rect 16856 6205 16865 6239
rect 16865 6205 16899 6239
rect 16899 6205 16908 6239
rect 16856 6196 16908 6205
rect 18420 6239 18472 6248
rect 18420 6205 18429 6239
rect 18429 6205 18463 6239
rect 18463 6205 18472 6239
rect 18420 6196 18472 6205
rect 19248 6196 19300 6248
rect 16764 6171 16816 6180
rect 16764 6137 16773 6171
rect 16773 6137 16807 6171
rect 16807 6137 16816 6171
rect 16764 6128 16816 6137
rect 18052 6128 18104 6180
rect 19524 6264 19576 6316
rect 19984 6264 20036 6316
rect 20168 6264 20220 6316
rect 20536 6264 20588 6316
rect 21088 6264 21140 6316
rect 23756 6264 23808 6316
rect 24032 6264 24084 6316
rect 19432 6196 19484 6248
rect 21548 6239 21600 6248
rect 21548 6205 21557 6239
rect 21557 6205 21591 6239
rect 21591 6205 21600 6239
rect 21548 6196 21600 6205
rect 22560 6196 22612 6248
rect 23664 6196 23716 6248
rect 24308 6196 24360 6248
rect 24768 6196 24820 6248
rect 25044 6196 25096 6248
rect 23296 6128 23348 6180
rect 23756 6128 23808 6180
rect 15476 6103 15528 6112
rect 15476 6069 15485 6103
rect 15485 6069 15519 6103
rect 15519 6069 15528 6103
rect 15476 6060 15528 6069
rect 17408 6103 17460 6112
rect 17408 6069 17417 6103
rect 17417 6069 17451 6103
rect 17451 6069 17460 6103
rect 17408 6060 17460 6069
rect 19432 6103 19484 6112
rect 19432 6069 19441 6103
rect 19441 6069 19475 6103
rect 19475 6069 19484 6103
rect 19432 6060 19484 6069
rect 19524 6060 19576 6112
rect 21180 6103 21232 6112
rect 21180 6069 21189 6103
rect 21189 6069 21223 6103
rect 21223 6069 21232 6103
rect 21180 6060 21232 6069
rect 22468 6060 22520 6112
rect 23664 6103 23716 6112
rect 23664 6069 23673 6103
rect 23673 6069 23707 6103
rect 23707 6069 23716 6103
rect 23664 6060 23716 6069
rect 25688 6060 25740 6112
rect 26240 6103 26292 6112
rect 26240 6069 26249 6103
rect 26249 6069 26283 6103
rect 26283 6069 26292 6103
rect 26240 6060 26292 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 2136 5856 2188 5908
rect 2964 5856 3016 5908
rect 3332 5856 3384 5908
rect 3976 5856 4028 5908
rect 4620 5899 4672 5908
rect 4620 5865 4629 5899
rect 4629 5865 4663 5899
rect 4663 5865 4672 5899
rect 4620 5856 4672 5865
rect 5356 5899 5408 5908
rect 5356 5865 5365 5899
rect 5365 5865 5399 5899
rect 5399 5865 5408 5899
rect 5356 5856 5408 5865
rect 6092 5856 6144 5908
rect 7104 5856 7156 5908
rect 8300 5899 8352 5908
rect 1400 5788 1452 5840
rect 3056 5720 3108 5772
rect 3608 5720 3660 5772
rect 6552 5788 6604 5840
rect 6920 5788 6972 5840
rect 7196 5831 7248 5840
rect 7196 5797 7230 5831
rect 7230 5797 7248 5831
rect 7196 5788 7248 5797
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 8852 5899 8904 5908
rect 8852 5865 8861 5899
rect 8861 5865 8895 5899
rect 8895 5865 8904 5899
rect 8852 5856 8904 5865
rect 11152 5856 11204 5908
rect 12716 5856 12768 5908
rect 12808 5856 12860 5908
rect 13360 5856 13412 5908
rect 14096 5899 14148 5908
rect 14096 5865 14105 5899
rect 14105 5865 14139 5899
rect 14139 5865 14148 5899
rect 14096 5856 14148 5865
rect 14280 5856 14332 5908
rect 15292 5899 15344 5908
rect 15292 5865 15301 5899
rect 15301 5865 15335 5899
rect 15335 5865 15344 5899
rect 15292 5856 15344 5865
rect 15568 5856 15620 5908
rect 16672 5899 16724 5908
rect 16672 5865 16681 5899
rect 16681 5865 16715 5899
rect 16715 5865 16724 5899
rect 16672 5856 16724 5865
rect 19156 5899 19208 5908
rect 19156 5865 19165 5899
rect 19165 5865 19199 5899
rect 19199 5865 19208 5899
rect 19156 5856 19208 5865
rect 19524 5856 19576 5908
rect 21364 5899 21416 5908
rect 21364 5865 21373 5899
rect 21373 5865 21407 5899
rect 21407 5865 21416 5899
rect 21364 5856 21416 5865
rect 21548 5856 21600 5908
rect 22468 5899 22520 5908
rect 22468 5865 22477 5899
rect 22477 5865 22511 5899
rect 22511 5865 22520 5899
rect 22468 5856 22520 5865
rect 22928 5899 22980 5908
rect 22928 5865 22937 5899
rect 22937 5865 22971 5899
rect 22971 5865 22980 5899
rect 22928 5856 22980 5865
rect 23664 5856 23716 5908
rect 9956 5831 10008 5840
rect 3516 5695 3568 5704
rect 3516 5661 3525 5695
rect 3525 5661 3559 5695
rect 3559 5661 3568 5695
rect 3516 5652 3568 5661
rect 5448 5652 5500 5704
rect 2688 5584 2740 5636
rect 5356 5584 5408 5636
rect 5540 5584 5592 5636
rect 6092 5720 6144 5772
rect 6828 5720 6880 5772
rect 9956 5797 9990 5831
rect 9990 5797 10008 5831
rect 9956 5788 10008 5797
rect 11888 5831 11940 5840
rect 11888 5797 11897 5831
rect 11897 5797 11931 5831
rect 11931 5797 11940 5831
rect 11888 5788 11940 5797
rect 17132 5831 17184 5840
rect 17132 5797 17166 5831
rect 17166 5797 17184 5831
rect 17132 5788 17184 5797
rect 19984 5831 20036 5840
rect 19984 5797 19993 5831
rect 19993 5797 20027 5831
rect 20027 5797 20036 5831
rect 19984 5788 20036 5797
rect 21272 5831 21324 5840
rect 21272 5797 21281 5831
rect 21281 5797 21315 5831
rect 21315 5797 21324 5831
rect 21272 5788 21324 5797
rect 23572 5788 23624 5840
rect 24308 5788 24360 5840
rect 26240 5831 26292 5840
rect 26240 5797 26249 5831
rect 26249 5797 26283 5831
rect 26283 5797 26292 5831
rect 26240 5788 26292 5797
rect 11980 5720 12032 5772
rect 12992 5763 13044 5772
rect 12992 5729 13026 5763
rect 13026 5729 13044 5763
rect 12992 5720 13044 5729
rect 15476 5720 15528 5772
rect 16120 5720 16172 5772
rect 17408 5720 17460 5772
rect 19524 5720 19576 5772
rect 20260 5763 20312 5772
rect 20260 5729 20269 5763
rect 20269 5729 20303 5763
rect 20303 5729 20312 5763
rect 20260 5720 20312 5729
rect 6552 5652 6604 5704
rect 9220 5652 9272 5704
rect 11796 5652 11848 5704
rect 12716 5695 12768 5704
rect 12716 5661 12725 5695
rect 12725 5661 12759 5695
rect 12759 5661 12768 5695
rect 12716 5652 12768 5661
rect 15292 5652 15344 5704
rect 16028 5652 16080 5704
rect 22744 5720 22796 5772
rect 23388 5720 23440 5772
rect 25044 5720 25096 5772
rect 25412 5720 25464 5772
rect 25780 5720 25832 5772
rect 21732 5652 21784 5704
rect 23020 5695 23072 5704
rect 23020 5661 23029 5695
rect 23029 5661 23063 5695
rect 23063 5661 23072 5695
rect 23020 5652 23072 5661
rect 1768 5559 1820 5568
rect 1768 5525 1777 5559
rect 1777 5525 1811 5559
rect 1811 5525 1820 5559
rect 1768 5516 1820 5525
rect 1860 5516 1912 5568
rect 3976 5516 4028 5568
rect 6368 5559 6420 5568
rect 6368 5525 6377 5559
rect 6377 5525 6411 5559
rect 6411 5525 6420 5559
rect 6368 5516 6420 5525
rect 9128 5584 9180 5636
rect 9220 5559 9272 5568
rect 9220 5525 9229 5559
rect 9229 5525 9263 5559
rect 9263 5525 9272 5559
rect 9220 5516 9272 5525
rect 13820 5584 13872 5636
rect 15384 5584 15436 5636
rect 18236 5627 18288 5636
rect 18236 5593 18245 5627
rect 18245 5593 18279 5627
rect 18279 5593 18288 5627
rect 18236 5584 18288 5593
rect 21548 5584 21600 5636
rect 22008 5584 22060 5636
rect 23940 5652 23992 5704
rect 24584 5695 24636 5704
rect 24584 5661 24593 5695
rect 24593 5661 24627 5695
rect 24627 5661 24636 5695
rect 24584 5652 24636 5661
rect 24768 5652 24820 5704
rect 18052 5516 18104 5568
rect 19340 5516 19392 5568
rect 21456 5516 21508 5568
rect 21824 5516 21876 5568
rect 23480 5584 23532 5636
rect 24952 5584 25004 5636
rect 25412 5559 25464 5568
rect 25412 5525 25421 5559
rect 25421 5525 25455 5559
rect 25455 5525 25464 5559
rect 25412 5516 25464 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2964 5312 3016 5364
rect 3240 5312 3292 5364
rect 6828 5312 6880 5364
rect 7012 5312 7064 5364
rect 2136 5244 2188 5296
rect 2688 5244 2740 5296
rect 1768 5176 1820 5228
rect 5724 5219 5776 5228
rect 2044 5151 2096 5160
rect 2044 5117 2053 5151
rect 2053 5117 2087 5151
rect 2087 5117 2096 5151
rect 2044 5108 2096 5117
rect 2504 5108 2556 5160
rect 3240 5151 3292 5160
rect 3240 5117 3249 5151
rect 3249 5117 3283 5151
rect 3283 5117 3292 5151
rect 3240 5108 3292 5117
rect 5724 5185 5733 5219
rect 5733 5185 5767 5219
rect 5767 5185 5776 5219
rect 5724 5176 5776 5185
rect 3516 5151 3568 5160
rect 3516 5117 3550 5151
rect 3550 5117 3568 5151
rect 3516 5108 3568 5117
rect 7840 5312 7892 5364
rect 8668 5355 8720 5364
rect 7932 5244 7984 5296
rect 8668 5321 8677 5355
rect 8677 5321 8711 5355
rect 8711 5321 8720 5355
rect 8668 5312 8720 5321
rect 10508 5355 10560 5364
rect 10508 5321 10517 5355
rect 10517 5321 10551 5355
rect 10551 5321 10560 5355
rect 10508 5312 10560 5321
rect 12624 5312 12676 5364
rect 13912 5355 13964 5364
rect 13912 5321 13921 5355
rect 13921 5321 13955 5355
rect 13955 5321 13964 5355
rect 13912 5312 13964 5321
rect 15292 5312 15344 5364
rect 17132 5312 17184 5364
rect 17684 5312 17736 5364
rect 16120 5244 16172 5296
rect 18328 5244 18380 5296
rect 10876 5176 10928 5228
rect 11152 5219 11204 5228
rect 11152 5185 11161 5219
rect 11161 5185 11195 5219
rect 11195 5185 11204 5219
rect 11152 5176 11204 5185
rect 13452 5176 13504 5228
rect 16028 5219 16080 5228
rect 16028 5185 16037 5219
rect 16037 5185 16071 5219
rect 16071 5185 16080 5219
rect 16028 5176 16080 5185
rect 19524 5312 19576 5364
rect 19984 5312 20036 5364
rect 20536 5312 20588 5364
rect 20996 5355 21048 5364
rect 20996 5321 21005 5355
rect 21005 5321 21039 5355
rect 21039 5321 21048 5355
rect 20996 5312 21048 5321
rect 20168 5219 20220 5228
rect 8024 5151 8076 5160
rect 8024 5117 8033 5151
rect 8033 5117 8067 5151
rect 8067 5117 8076 5151
rect 8024 5108 8076 5117
rect 10324 5040 10376 5092
rect 11888 5108 11940 5160
rect 13728 5108 13780 5160
rect 14280 5108 14332 5160
rect 15384 5108 15436 5160
rect 18420 5108 18472 5160
rect 20168 5185 20177 5219
rect 20177 5185 20211 5219
rect 20211 5185 20220 5219
rect 20168 5176 20220 5185
rect 21640 5219 21692 5228
rect 21640 5185 21649 5219
rect 21649 5185 21683 5219
rect 21683 5185 21692 5219
rect 21640 5176 21692 5185
rect 22744 5312 22796 5364
rect 22928 5355 22980 5364
rect 22928 5321 22937 5355
rect 22937 5321 22971 5355
rect 22971 5321 22980 5355
rect 22928 5312 22980 5321
rect 23664 5355 23716 5364
rect 23664 5321 23673 5355
rect 23673 5321 23707 5355
rect 23707 5321 23716 5355
rect 23664 5312 23716 5321
rect 24768 5355 24820 5364
rect 24768 5321 24777 5355
rect 24777 5321 24811 5355
rect 24811 5321 24820 5355
rect 24768 5312 24820 5321
rect 25044 5355 25096 5364
rect 25044 5321 25053 5355
rect 25053 5321 25087 5355
rect 25087 5321 25096 5355
rect 25044 5312 25096 5321
rect 25872 5355 25924 5364
rect 25872 5321 25881 5355
rect 25881 5321 25915 5355
rect 25915 5321 25924 5355
rect 25872 5312 25924 5321
rect 22192 5244 22244 5296
rect 25228 5244 25280 5296
rect 22100 5176 22152 5228
rect 19064 5108 19116 5160
rect 21548 5151 21600 5160
rect 4620 5015 4672 5024
rect 4620 4981 4629 5015
rect 4629 4981 4663 5015
rect 4663 4981 4672 5015
rect 4620 4972 4672 4981
rect 5356 4972 5408 5024
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 6552 4972 6604 4981
rect 7748 4972 7800 5024
rect 9496 5015 9548 5024
rect 9496 4981 9505 5015
rect 9505 4981 9539 5015
rect 9539 4981 9548 5015
rect 9496 4972 9548 4981
rect 11520 5040 11572 5092
rect 15108 5040 15160 5092
rect 11336 4972 11388 5024
rect 12716 4972 12768 5024
rect 12992 4972 13044 5024
rect 14004 4972 14056 5024
rect 14556 5015 14608 5024
rect 14556 4981 14565 5015
rect 14565 4981 14599 5015
rect 14599 4981 14608 5015
rect 14556 4972 14608 4981
rect 15384 5015 15436 5024
rect 15384 4981 15393 5015
rect 15393 4981 15427 5015
rect 15427 4981 15436 5015
rect 15384 4972 15436 4981
rect 16488 4972 16540 5024
rect 20168 5040 20220 5092
rect 18328 4972 18380 5024
rect 21180 5015 21232 5024
rect 21180 4981 21189 5015
rect 21189 4981 21223 5015
rect 21223 4981 21232 5015
rect 21180 4972 21232 4981
rect 21548 5117 21557 5151
rect 21557 5117 21591 5151
rect 21591 5117 21600 5151
rect 21548 5108 21600 5117
rect 21456 5040 21508 5092
rect 22652 5040 22704 5092
rect 23940 5176 23992 5228
rect 24308 5219 24360 5228
rect 24308 5185 24317 5219
rect 24317 5185 24351 5219
rect 24351 5185 24360 5219
rect 24308 5176 24360 5185
rect 24032 5151 24084 5160
rect 24032 5117 24041 5151
rect 24041 5117 24075 5151
rect 24075 5117 24084 5151
rect 24032 5108 24084 5117
rect 25872 5108 25924 5160
rect 25228 4972 25280 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 2320 4811 2372 4820
rect 2320 4777 2329 4811
rect 2329 4777 2363 4811
rect 2363 4777 2372 4811
rect 2320 4768 2372 4777
rect 2688 4768 2740 4820
rect 4068 4768 4120 4820
rect 4804 4768 4856 4820
rect 8944 4811 8996 4820
rect 8944 4777 8953 4811
rect 8953 4777 8987 4811
rect 8987 4777 8996 4811
rect 8944 4768 8996 4777
rect 9680 4768 9732 4820
rect 10876 4811 10928 4820
rect 10876 4777 10885 4811
rect 10885 4777 10919 4811
rect 10919 4777 10928 4811
rect 10876 4768 10928 4777
rect 11520 4811 11572 4820
rect 11520 4777 11529 4811
rect 11529 4777 11563 4811
rect 11563 4777 11572 4811
rect 11520 4768 11572 4777
rect 13820 4768 13872 4820
rect 14372 4768 14424 4820
rect 15108 4811 15160 4820
rect 15108 4777 15117 4811
rect 15117 4777 15151 4811
rect 15151 4777 15160 4811
rect 15108 4768 15160 4777
rect 18880 4768 18932 4820
rect 20720 4811 20772 4820
rect 20720 4777 20729 4811
rect 20729 4777 20763 4811
rect 20763 4777 20772 4811
rect 20720 4768 20772 4777
rect 21732 4768 21784 4820
rect 23020 4768 23072 4820
rect 24032 4768 24084 4820
rect 24308 4768 24360 4820
rect 4620 4700 4672 4752
rect 6000 4700 6052 4752
rect 8300 4700 8352 4752
rect 9956 4743 10008 4752
rect 9956 4709 9965 4743
rect 9965 4709 9999 4743
rect 9999 4709 10008 4743
rect 9956 4700 10008 4709
rect 13176 4743 13228 4752
rect 13176 4709 13185 4743
rect 13185 4709 13219 4743
rect 13219 4709 13228 4743
rect 13176 4700 13228 4709
rect 17868 4700 17920 4752
rect 18604 4700 18656 4752
rect 2320 4632 2372 4684
rect 3424 4632 3476 4684
rect 2964 4564 3016 4616
rect 3516 4564 3568 4616
rect 3240 4496 3292 4548
rect 10784 4675 10836 4684
rect 10784 4641 10793 4675
rect 10793 4641 10827 4675
rect 10827 4641 10836 4675
rect 10784 4632 10836 4641
rect 12440 4675 12492 4684
rect 12440 4641 12449 4675
rect 12449 4641 12483 4675
rect 12483 4641 12492 4675
rect 12440 4632 12492 4641
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 11152 4564 11204 4616
rect 12532 4607 12584 4616
rect 12532 4573 12541 4607
rect 12541 4573 12575 4607
rect 12575 4573 12584 4607
rect 12532 4564 12584 4573
rect 13728 4632 13780 4684
rect 14096 4607 14148 4616
rect 3976 4428 4028 4480
rect 4252 4428 4304 4480
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 14096 4564 14148 4573
rect 17224 4632 17276 4684
rect 18420 4675 18472 4684
rect 18420 4641 18429 4675
rect 18429 4641 18463 4675
rect 18463 4641 18472 4675
rect 18420 4632 18472 4641
rect 18972 4675 19024 4684
rect 18972 4641 18981 4675
rect 18981 4641 19015 4675
rect 19015 4641 19024 4675
rect 18972 4632 19024 4641
rect 21272 4675 21324 4684
rect 21272 4641 21281 4675
rect 21281 4641 21315 4675
rect 21315 4641 21324 4675
rect 21272 4632 21324 4641
rect 15660 4564 15712 4616
rect 16120 4607 16172 4616
rect 16120 4573 16129 4607
rect 16129 4573 16163 4607
rect 16163 4573 16172 4607
rect 16120 4564 16172 4573
rect 19156 4607 19208 4616
rect 19156 4573 19165 4607
rect 19165 4573 19199 4607
rect 19199 4573 19208 4607
rect 19156 4564 19208 4573
rect 20720 4564 20772 4616
rect 23112 4700 23164 4752
rect 25044 4743 25096 4752
rect 25044 4709 25053 4743
rect 25053 4709 25087 4743
rect 25087 4709 25096 4743
rect 25044 4700 25096 4709
rect 22836 4675 22888 4684
rect 22836 4641 22845 4675
rect 22845 4641 22879 4675
rect 22879 4641 22888 4675
rect 22836 4632 22888 4641
rect 24676 4632 24728 4684
rect 23020 4607 23072 4616
rect 23020 4573 23029 4607
rect 23029 4573 23063 4607
rect 23063 4573 23072 4607
rect 23020 4564 23072 4573
rect 23664 4564 23716 4616
rect 24216 4564 24268 4616
rect 18788 4496 18840 4548
rect 23296 4496 23348 4548
rect 23388 4496 23440 4548
rect 8852 4428 8904 4480
rect 9496 4428 9548 4480
rect 10324 4471 10376 4480
rect 10324 4437 10333 4471
rect 10333 4437 10367 4471
rect 10367 4437 10376 4471
rect 10324 4428 10376 4437
rect 12072 4471 12124 4480
rect 12072 4437 12081 4471
rect 12081 4437 12115 4471
rect 12115 4437 12124 4471
rect 12072 4428 12124 4437
rect 14740 4471 14792 4480
rect 14740 4437 14749 4471
rect 14749 4437 14783 4471
rect 14783 4437 14792 4471
rect 14740 4428 14792 4437
rect 16028 4471 16080 4480
rect 16028 4437 16037 4471
rect 16037 4437 16071 4471
rect 16071 4437 16080 4471
rect 16028 4428 16080 4437
rect 16856 4428 16908 4480
rect 18696 4428 18748 4480
rect 19984 4471 20036 4480
rect 19984 4437 19993 4471
rect 19993 4437 20027 4471
rect 20027 4437 20036 4471
rect 19984 4428 20036 4437
rect 21916 4428 21968 4480
rect 23572 4428 23624 4480
rect 24216 4428 24268 4480
rect 24768 4428 24820 4480
rect 26240 4471 26292 4480
rect 26240 4437 26249 4471
rect 26249 4437 26283 4471
rect 26283 4437 26292 4471
rect 26240 4428 26292 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 2964 4267 3016 4276
rect 2964 4233 2973 4267
rect 2973 4233 3007 4267
rect 3007 4233 3016 4267
rect 2964 4224 3016 4233
rect 3424 4267 3476 4276
rect 3424 4233 3433 4267
rect 3433 4233 3467 4267
rect 3467 4233 3476 4267
rect 3424 4224 3476 4233
rect 5356 4224 5408 4276
rect 2320 4156 2372 4208
rect 5448 4156 5500 4208
rect 6092 4156 6144 4208
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 4988 4131 5040 4140
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 2136 4020 2188 4072
rect 2688 4020 2740 4072
rect 9496 4156 9548 4208
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 13544 4156 13596 4208
rect 9128 4088 9180 4097
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 12348 4088 12400 4140
rect 12440 4088 12492 4140
rect 13176 4131 13228 4140
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13176 4088 13228 4097
rect 13452 4088 13504 4140
rect 18972 4224 19024 4276
rect 20168 4224 20220 4276
rect 23112 4224 23164 4276
rect 24676 4267 24728 4276
rect 24676 4233 24685 4267
rect 24685 4233 24719 4267
rect 24719 4233 24728 4267
rect 24676 4224 24728 4233
rect 25228 4224 25280 4276
rect 14096 4156 14148 4208
rect 15016 4156 15068 4208
rect 15384 4156 15436 4208
rect 14924 4131 14976 4140
rect 6092 4020 6144 4072
rect 6184 4020 6236 4072
rect 6368 4020 6420 4072
rect 2504 3952 2556 4004
rect 3884 3995 3936 4004
rect 3884 3961 3893 3995
rect 3893 3961 3927 3995
rect 3927 3961 3936 3995
rect 3884 3952 3936 3961
rect 4160 3952 4212 4004
rect 5264 3952 5316 4004
rect 9312 4020 9364 4072
rect 11060 4020 11112 4072
rect 14924 4097 14933 4131
rect 14933 4097 14967 4131
rect 14967 4097 14976 4131
rect 14924 4088 14976 4097
rect 15292 4131 15344 4140
rect 15292 4097 15301 4131
rect 15301 4097 15335 4131
rect 15335 4097 15344 4131
rect 15292 4088 15344 4097
rect 16396 4088 16448 4140
rect 16856 4131 16908 4140
rect 16856 4097 16865 4131
rect 16865 4097 16899 4131
rect 16899 4097 16908 4131
rect 16856 4088 16908 4097
rect 18420 4156 18472 4208
rect 18696 4156 18748 4208
rect 19984 4156 20036 4208
rect 14372 4020 14424 4072
rect 14648 4063 14700 4072
rect 14648 4029 14657 4063
rect 14657 4029 14691 4063
rect 14691 4029 14700 4063
rect 14648 4020 14700 4029
rect 17224 4020 17276 4072
rect 18236 4020 18288 4072
rect 18880 4020 18932 4072
rect 20260 4020 20312 4072
rect 20352 4020 20404 4072
rect 26240 4156 26292 4208
rect 21732 4131 21784 4140
rect 21732 4097 21741 4131
rect 21741 4097 21775 4131
rect 21775 4097 21784 4131
rect 21732 4088 21784 4097
rect 23480 4088 23532 4140
rect 24952 4088 25004 4140
rect 20996 4020 21048 4072
rect 22560 4020 22612 4072
rect 23756 4020 23808 4072
rect 7472 3952 7524 4004
rect 14740 3995 14792 4004
rect 2688 3884 2740 3936
rect 3792 3927 3844 3936
rect 3792 3893 3801 3927
rect 3801 3893 3835 3927
rect 3835 3893 3844 3927
rect 3792 3884 3844 3893
rect 4620 3884 4672 3936
rect 5080 3884 5132 3936
rect 6184 3927 6236 3936
rect 6184 3893 6193 3927
rect 6193 3893 6227 3927
rect 6227 3893 6236 3927
rect 6552 3927 6604 3936
rect 6184 3884 6236 3893
rect 6552 3893 6561 3927
rect 6561 3893 6595 3927
rect 6595 3893 6604 3927
rect 6552 3884 6604 3893
rect 6920 3884 6972 3936
rect 8852 3927 8904 3936
rect 8852 3893 8861 3927
rect 8861 3893 8895 3927
rect 8895 3893 8904 3927
rect 8852 3884 8904 3893
rect 9404 3884 9456 3936
rect 10784 3884 10836 3936
rect 10968 3884 11020 3936
rect 11980 3884 12032 3936
rect 12532 3884 12584 3936
rect 14740 3961 14749 3995
rect 14749 3961 14783 3995
rect 14783 3961 14792 3995
rect 14740 3952 14792 3961
rect 20168 3952 20220 4004
rect 22100 3952 22152 4004
rect 22192 3952 22244 4004
rect 25044 4063 25096 4072
rect 25044 4029 25053 4063
rect 25053 4029 25087 4063
rect 25087 4029 25096 4063
rect 25044 4020 25096 4029
rect 23940 3952 23992 4004
rect 14280 3927 14332 3936
rect 14280 3893 14289 3927
rect 14289 3893 14323 3927
rect 14323 3893 14332 3927
rect 14280 3884 14332 3893
rect 15292 3884 15344 3936
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 16212 3927 16264 3936
rect 16212 3893 16221 3927
rect 16221 3893 16255 3927
rect 16255 3893 16264 3927
rect 16212 3884 16264 3893
rect 18052 3927 18104 3936
rect 18052 3893 18061 3927
rect 18061 3893 18095 3927
rect 18095 3893 18104 3927
rect 18052 3884 18104 3893
rect 19432 3927 19484 3936
rect 19432 3893 19441 3927
rect 19441 3893 19475 3927
rect 19475 3893 19484 3927
rect 19432 3884 19484 3893
rect 20996 3884 21048 3936
rect 21180 3927 21232 3936
rect 21180 3893 21189 3927
rect 21189 3893 21223 3927
rect 21223 3893 21232 3927
rect 21180 3884 21232 3893
rect 22836 3927 22888 3936
rect 22836 3893 22845 3927
rect 22845 3893 22879 3927
rect 22879 3893 22888 3927
rect 22836 3884 22888 3893
rect 23388 3927 23440 3936
rect 23388 3893 23397 3927
rect 23397 3893 23431 3927
rect 23431 3893 23440 3927
rect 23388 3884 23440 3893
rect 23756 3884 23808 3936
rect 24032 3927 24084 3936
rect 24032 3893 24041 3927
rect 24041 3893 24075 3927
rect 24075 3893 24084 3927
rect 24032 3884 24084 3893
rect 25412 3927 25464 3936
rect 25412 3893 25421 3927
rect 25421 3893 25455 3927
rect 25455 3893 25464 3927
rect 25412 3884 25464 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 2688 3680 2740 3732
rect 3792 3680 3844 3732
rect 4068 3723 4120 3732
rect 4068 3689 4077 3723
rect 4077 3689 4111 3723
rect 4111 3689 4120 3723
rect 4068 3680 4120 3689
rect 4528 3723 4580 3732
rect 4528 3689 4537 3723
rect 4537 3689 4571 3723
rect 4571 3689 4580 3723
rect 4528 3680 4580 3689
rect 5264 3723 5316 3732
rect 5264 3689 5273 3723
rect 5273 3689 5307 3723
rect 5307 3689 5316 3723
rect 5264 3680 5316 3689
rect 9312 3723 9364 3732
rect 9312 3689 9321 3723
rect 9321 3689 9355 3723
rect 9355 3689 9364 3723
rect 9312 3680 9364 3689
rect 9680 3723 9732 3732
rect 9680 3689 9689 3723
rect 9689 3689 9723 3723
rect 9723 3689 9732 3723
rect 10140 3723 10192 3732
rect 9680 3680 9732 3689
rect 10140 3689 10149 3723
rect 10149 3689 10183 3723
rect 10183 3689 10192 3723
rect 10140 3680 10192 3689
rect 10876 3680 10928 3732
rect 11152 3680 11204 3732
rect 13084 3723 13136 3732
rect 13084 3689 13093 3723
rect 13093 3689 13127 3723
rect 13127 3689 13136 3723
rect 13084 3680 13136 3689
rect 13728 3723 13780 3732
rect 13728 3689 13737 3723
rect 13737 3689 13771 3723
rect 13771 3689 13780 3723
rect 13728 3680 13780 3689
rect 14188 3723 14240 3732
rect 14188 3689 14197 3723
rect 14197 3689 14231 3723
rect 14231 3689 14240 3723
rect 14188 3680 14240 3689
rect 14648 3680 14700 3732
rect 15476 3680 15528 3732
rect 16304 3723 16356 3732
rect 16304 3689 16313 3723
rect 16313 3689 16347 3723
rect 16347 3689 16356 3723
rect 16304 3680 16356 3689
rect 16488 3680 16540 3732
rect 18604 3723 18656 3732
rect 18604 3689 18613 3723
rect 18613 3689 18647 3723
rect 18647 3689 18656 3723
rect 18604 3680 18656 3689
rect 19064 3680 19116 3732
rect 20352 3680 20404 3732
rect 21364 3723 21416 3732
rect 2320 3655 2372 3664
rect 2320 3621 2329 3655
rect 2329 3621 2363 3655
rect 2363 3621 2372 3655
rect 2320 3612 2372 3621
rect 2044 3544 2096 3596
rect 2228 3476 2280 3528
rect 4620 3612 4672 3664
rect 4436 3587 4488 3596
rect 4436 3553 4445 3587
rect 4445 3553 4479 3587
rect 4479 3553 4488 3587
rect 4436 3544 4488 3553
rect 6184 3612 6236 3664
rect 8852 3612 8904 3664
rect 3976 3476 4028 3528
rect 5172 3476 5224 3528
rect 4804 3340 4856 3392
rect 5908 3544 5960 3596
rect 8576 3587 8628 3596
rect 8576 3553 8585 3587
rect 8585 3553 8619 3587
rect 8619 3553 8628 3587
rect 8576 3544 8628 3553
rect 9864 3544 9916 3596
rect 11612 3612 11664 3664
rect 16764 3612 16816 3664
rect 17592 3612 17644 3664
rect 17776 3655 17828 3664
rect 17776 3621 17785 3655
rect 17785 3621 17819 3655
rect 17819 3621 17828 3655
rect 17776 3612 17828 3621
rect 11244 3544 11296 3596
rect 12256 3544 12308 3596
rect 17040 3544 17092 3596
rect 11612 3476 11664 3528
rect 14924 3476 14976 3528
rect 15384 3476 15436 3528
rect 16856 3476 16908 3528
rect 17224 3476 17276 3528
rect 17960 3519 18012 3528
rect 17960 3485 17969 3519
rect 17969 3485 18003 3519
rect 18003 3485 18012 3519
rect 17960 3476 18012 3485
rect 7840 3408 7892 3460
rect 14464 3408 14516 3460
rect 19524 3612 19576 3664
rect 21364 3689 21373 3723
rect 21373 3689 21407 3723
rect 21407 3689 21416 3723
rect 21364 3680 21416 3689
rect 23572 3680 23624 3732
rect 24768 3680 24820 3732
rect 21456 3612 21508 3664
rect 23480 3655 23532 3664
rect 23480 3621 23489 3655
rect 23489 3621 23523 3655
rect 23523 3621 23532 3655
rect 23480 3612 23532 3621
rect 21272 3587 21324 3596
rect 21272 3553 21281 3587
rect 21281 3553 21315 3587
rect 21315 3553 21324 3587
rect 21272 3544 21324 3553
rect 22100 3544 22152 3596
rect 19984 3476 20036 3528
rect 7288 3340 7340 3392
rect 8668 3340 8720 3392
rect 8760 3383 8812 3392
rect 8760 3349 8769 3383
rect 8769 3349 8803 3383
rect 8803 3349 8812 3383
rect 15568 3383 15620 3392
rect 8760 3340 8812 3349
rect 15568 3349 15577 3383
rect 15577 3349 15611 3383
rect 15611 3349 15620 3383
rect 15568 3340 15620 3349
rect 15844 3383 15896 3392
rect 15844 3349 15853 3383
rect 15853 3349 15887 3383
rect 15887 3349 15896 3383
rect 15844 3340 15896 3349
rect 17408 3383 17460 3392
rect 17408 3349 17417 3383
rect 17417 3349 17451 3383
rect 17451 3349 17460 3383
rect 17408 3340 17460 3349
rect 19984 3383 20036 3392
rect 19984 3349 19993 3383
rect 19993 3349 20027 3383
rect 20027 3349 20036 3383
rect 21732 3476 21784 3528
rect 22008 3476 22060 3528
rect 22928 3519 22980 3528
rect 22928 3485 22937 3519
rect 22937 3485 22971 3519
rect 22971 3485 22980 3519
rect 22928 3476 22980 3485
rect 23020 3408 23072 3460
rect 23664 3476 23716 3528
rect 24676 3519 24728 3528
rect 24676 3485 24685 3519
rect 24685 3485 24719 3519
rect 24719 3485 24728 3519
rect 24676 3476 24728 3485
rect 24032 3451 24084 3460
rect 24032 3417 24041 3451
rect 24041 3417 24075 3451
rect 24075 3417 24084 3451
rect 24032 3408 24084 3417
rect 19984 3340 20036 3349
rect 23480 3340 23532 3392
rect 23848 3383 23900 3392
rect 23848 3349 23857 3383
rect 23857 3349 23891 3383
rect 23891 3349 23900 3383
rect 23848 3340 23900 3349
rect 24768 3340 24820 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 1768 3068 1820 3120
rect 2688 3068 2740 3120
rect 2964 3000 3016 3052
rect 2504 2975 2556 2984
rect 2504 2941 2513 2975
rect 2513 2941 2547 2975
rect 2547 2941 2556 2975
rect 2504 2932 2556 2941
rect 3700 3136 3752 3188
rect 4436 3136 4488 3188
rect 4988 3179 5040 3188
rect 4988 3145 4997 3179
rect 4997 3145 5031 3179
rect 5031 3145 5040 3179
rect 4988 3136 5040 3145
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 6184 3136 6236 3188
rect 7196 3136 7248 3188
rect 9864 3136 9916 3188
rect 10876 3136 10928 3188
rect 11152 3179 11204 3188
rect 11152 3145 11161 3179
rect 11161 3145 11195 3179
rect 11195 3145 11204 3179
rect 11152 3136 11204 3145
rect 12256 3179 12308 3188
rect 12256 3145 12265 3179
rect 12265 3145 12299 3179
rect 12299 3145 12308 3179
rect 12256 3136 12308 3145
rect 15476 3136 15528 3188
rect 15568 3136 15620 3188
rect 3516 3068 3568 3120
rect 4528 3068 4580 3120
rect 6828 3111 6880 3120
rect 6828 3077 6837 3111
rect 6837 3077 6871 3111
rect 6871 3077 6880 3111
rect 6828 3068 6880 3077
rect 10140 3068 10192 3120
rect 12164 3068 12216 3120
rect 3976 3000 4028 3052
rect 5540 3000 5592 3052
rect 7288 3000 7340 3052
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 11152 3000 11204 3052
rect 11428 3000 11480 3052
rect 12256 3000 12308 3052
rect 13728 3000 13780 3052
rect 6000 2932 6052 2984
rect 7196 2975 7248 2984
rect 7196 2941 7205 2975
rect 7205 2941 7239 2975
rect 7239 2941 7248 2975
rect 7196 2932 7248 2941
rect 8116 2932 8168 2984
rect 8208 2932 8260 2984
rect 8668 2975 8720 2984
rect 8668 2941 8702 2975
rect 8702 2941 8720 2975
rect 8668 2932 8720 2941
rect 9772 2932 9824 2984
rect 11244 2975 11296 2984
rect 11244 2941 11253 2975
rect 11253 2941 11287 2975
rect 11287 2941 11296 2975
rect 11244 2932 11296 2941
rect 2688 2864 2740 2916
rect 6368 2864 6420 2916
rect 1216 2796 1268 2848
rect 3700 2796 3752 2848
rect 7104 2864 7156 2916
rect 14004 2864 14056 2916
rect 7932 2839 7984 2848
rect 7932 2805 7941 2839
rect 7941 2805 7975 2839
rect 7975 2805 7984 2839
rect 7932 2796 7984 2805
rect 8208 2839 8260 2848
rect 8208 2805 8217 2839
rect 8217 2805 8251 2839
rect 8251 2805 8260 2839
rect 8208 2796 8260 2805
rect 9772 2839 9824 2848
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 9772 2796 9824 2805
rect 11428 2839 11480 2848
rect 11428 2805 11437 2839
rect 11437 2805 11471 2839
rect 11471 2805 11480 2839
rect 11428 2796 11480 2805
rect 11612 2796 11664 2848
rect 11796 2839 11848 2848
rect 11796 2805 11805 2839
rect 11805 2805 11839 2839
rect 11839 2805 11848 2839
rect 11796 2796 11848 2805
rect 13268 2839 13320 2848
rect 13268 2805 13277 2839
rect 13277 2805 13311 2839
rect 13311 2805 13320 2839
rect 13268 2796 13320 2805
rect 13636 2839 13688 2848
rect 13636 2805 13645 2839
rect 13645 2805 13679 2839
rect 13679 2805 13688 2839
rect 13636 2796 13688 2805
rect 14464 2796 14516 2848
rect 14924 2932 14976 2984
rect 15384 2932 15436 2984
rect 15568 2932 15620 2984
rect 17960 3136 18012 3188
rect 18788 3136 18840 3188
rect 19248 3136 19300 3188
rect 20720 3136 20772 3188
rect 22008 3136 22060 3188
rect 22284 3179 22336 3188
rect 22284 3145 22293 3179
rect 22293 3145 22327 3179
rect 22327 3145 22336 3179
rect 22284 3136 22336 3145
rect 23664 3179 23716 3188
rect 23664 3145 23673 3179
rect 23673 3145 23707 3179
rect 23707 3145 23716 3179
rect 23664 3136 23716 3145
rect 24676 3179 24728 3188
rect 24676 3145 24685 3179
rect 24685 3145 24719 3179
rect 24719 3145 24728 3179
rect 24676 3136 24728 3145
rect 16856 3068 16908 3120
rect 19984 3068 20036 3120
rect 20076 3043 20128 3052
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20076 3000 20128 3009
rect 23572 3068 23624 3120
rect 24216 3068 24268 3120
rect 21732 3043 21784 3052
rect 21732 3009 21741 3043
rect 21741 3009 21775 3043
rect 21775 3009 21784 3043
rect 21732 3000 21784 3009
rect 24032 3000 24084 3052
rect 24308 3043 24360 3052
rect 24308 3009 24317 3043
rect 24317 3009 24351 3043
rect 24351 3009 24360 3043
rect 24308 3000 24360 3009
rect 26240 3043 26292 3052
rect 26240 3009 26249 3043
rect 26249 3009 26283 3043
rect 26283 3009 26292 3043
rect 26240 3000 26292 3009
rect 17040 2932 17092 2984
rect 17592 2932 17644 2984
rect 18144 2932 18196 2984
rect 18420 2975 18472 2984
rect 18420 2941 18429 2975
rect 18429 2941 18463 2975
rect 18463 2941 18472 2975
rect 18420 2932 18472 2941
rect 18512 2975 18564 2984
rect 18512 2941 18521 2975
rect 18521 2941 18555 2975
rect 18555 2941 18564 2975
rect 18512 2932 18564 2941
rect 20812 2932 20864 2984
rect 18604 2864 18656 2916
rect 20720 2907 20772 2916
rect 20720 2873 20729 2907
rect 20729 2873 20763 2907
rect 20763 2873 20772 2907
rect 21272 2932 21324 2984
rect 22284 2932 22336 2984
rect 22468 2932 22520 2984
rect 23572 2932 23624 2984
rect 23756 2932 23808 2984
rect 24676 2932 24728 2984
rect 25780 2975 25832 2984
rect 25780 2941 25789 2975
rect 25789 2941 25823 2975
rect 25823 2941 25832 2975
rect 25780 2932 25832 2941
rect 20720 2864 20772 2873
rect 20996 2864 21048 2916
rect 25688 2864 25740 2916
rect 18052 2839 18104 2848
rect 18052 2805 18061 2839
rect 18061 2805 18095 2839
rect 18095 2805 18104 2839
rect 18052 2796 18104 2805
rect 21364 2796 21416 2848
rect 23112 2796 23164 2848
rect 23756 2796 23808 2848
rect 24216 2796 24268 2848
rect 25044 2839 25096 2848
rect 25044 2805 25053 2839
rect 25053 2805 25087 2839
rect 25087 2805 25096 2839
rect 25044 2796 25096 2805
rect 25136 2796 25188 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 2228 2592 2280 2644
rect 2872 2635 2924 2644
rect 2872 2601 2881 2635
rect 2881 2601 2915 2635
rect 2915 2601 2924 2635
rect 2872 2592 2924 2601
rect 5540 2592 5592 2644
rect 6552 2592 6604 2644
rect 8300 2635 8352 2644
rect 2780 2567 2832 2576
rect 2780 2533 2789 2567
rect 2789 2533 2823 2567
rect 2823 2533 2832 2567
rect 3700 2567 3752 2576
rect 2780 2524 2832 2533
rect 3700 2533 3709 2567
rect 3709 2533 3743 2567
rect 3743 2533 3752 2567
rect 3700 2524 3752 2533
rect 1952 2456 2004 2508
rect 4436 2456 4488 2508
rect 5080 2456 5132 2508
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 14556 2592 14608 2644
rect 14924 2635 14976 2644
rect 14924 2601 14933 2635
rect 14933 2601 14967 2635
rect 14967 2601 14976 2635
rect 14924 2592 14976 2601
rect 18972 2592 19024 2644
rect 22008 2592 22060 2644
rect 22284 2635 22336 2644
rect 22284 2601 22293 2635
rect 22293 2601 22327 2635
rect 22327 2601 22336 2635
rect 22284 2592 22336 2601
rect 23940 2592 23992 2644
rect 7932 2524 7984 2576
rect 10876 2524 10928 2576
rect 13728 2524 13780 2576
rect 15568 2524 15620 2576
rect 18144 2524 18196 2576
rect 8208 2456 8260 2508
rect 11796 2456 11848 2508
rect 12992 2456 13044 2508
rect 14464 2456 14516 2508
rect 15292 2456 15344 2508
rect 4252 2388 4304 2440
rect 20904 2524 20956 2576
rect 22560 2524 22612 2576
rect 23480 2524 23532 2576
rect 24768 2524 24820 2576
rect 20076 2456 20128 2508
rect 22744 2499 22796 2508
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 1952 2295 2004 2304
rect 1952 2261 1961 2295
rect 1961 2261 1995 2295
rect 1995 2261 2004 2295
rect 1952 2252 2004 2261
rect 11244 2252 11296 2304
rect 14556 2252 14608 2304
rect 18696 2320 18748 2372
rect 20536 2363 20588 2372
rect 20536 2329 20545 2363
rect 20545 2329 20579 2363
rect 20579 2329 20588 2363
rect 22744 2465 22753 2499
rect 22753 2465 22787 2499
rect 22787 2465 22796 2499
rect 22744 2456 22796 2465
rect 23020 2456 23072 2508
rect 24308 2456 24360 2508
rect 24492 2499 24544 2508
rect 24492 2465 24501 2499
rect 24501 2465 24535 2499
rect 24535 2465 24544 2499
rect 24492 2456 24544 2465
rect 24676 2456 24728 2508
rect 26424 2499 26476 2508
rect 26424 2465 26433 2499
rect 26433 2465 26467 2499
rect 26467 2465 26476 2499
rect 26424 2456 26476 2465
rect 21732 2431 21784 2440
rect 21732 2397 21741 2431
rect 21741 2397 21775 2431
rect 21775 2397 21784 2431
rect 21732 2388 21784 2397
rect 22928 2388 22980 2440
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 20536 2320 20588 2329
rect 16856 2295 16908 2304
rect 16856 2261 16865 2295
rect 16865 2261 16899 2295
rect 16899 2261 16908 2295
rect 16856 2252 16908 2261
rect 18328 2295 18380 2304
rect 18328 2261 18337 2295
rect 18337 2261 18371 2295
rect 18371 2261 18380 2295
rect 18328 2252 18380 2261
rect 19892 2252 19944 2304
rect 20904 2295 20956 2304
rect 20904 2261 20913 2295
rect 20913 2261 20947 2295
rect 20947 2261 20956 2295
rect 20904 2252 20956 2261
rect 22928 2295 22980 2304
rect 22928 2261 22937 2295
rect 22937 2261 22971 2295
rect 22971 2261 22980 2295
rect 22928 2252 22980 2261
rect 24768 2252 24820 2304
rect 25504 2252 25556 2304
rect 25780 2295 25832 2304
rect 25780 2261 25789 2295
rect 25789 2261 25823 2295
rect 25823 2261 25832 2295
rect 25780 2252 25832 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 11336 2048 11388 2100
rect 17408 2048 17460 2100
rect 14648 1844 14700 1896
rect 17500 1844 17552 1896
rect 5632 1640 5684 1692
rect 6644 1640 6696 1692
rect 15108 1572 15160 1624
rect 17960 1572 18012 1624
rect 24952 552 25004 604
rect 25412 552 25464 604
rect 14832 212 14884 264
rect 18144 212 18196 264
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1122 27704 1178 27713
rect 1122 27639 1178 27648
rect 308 24834 336 27520
rect 662 27160 718 27169
rect 662 27095 718 27104
rect 572 25152 624 25158
rect 572 25094 624 25100
rect 32 24806 336 24834
rect 32 12345 60 24806
rect 584 20097 612 25094
rect 676 24449 704 27095
rect 662 24440 718 24449
rect 662 24375 718 24384
rect 676 21486 704 24375
rect 664 21480 716 21486
rect 664 21422 716 21428
rect 570 20088 626 20097
rect 570 20023 626 20032
rect 860 12374 888 27520
rect 1030 25936 1086 25945
rect 1030 25871 1086 25880
rect 938 24848 994 24857
rect 938 24783 994 24792
rect 952 20058 980 24783
rect 1044 22098 1072 25871
rect 1136 24342 1164 27639
rect 1398 27520 1454 28000
rect 2042 27520 2098 28000
rect 2594 27520 2650 28000
rect 3146 27520 3202 28000
rect 3790 27520 3846 28000
rect 4342 27520 4398 28000
rect 4894 27520 4950 28000
rect 5538 27520 5594 28000
rect 6090 27520 6146 28000
rect 6642 27520 6698 28000
rect 7286 27520 7342 28000
rect 7838 27520 7894 28000
rect 8390 27520 8446 28000
rect 9034 27520 9090 28000
rect 9586 27520 9642 28000
rect 10138 27520 10194 28000
rect 10782 27520 10838 28000
rect 11334 27520 11390 28000
rect 11886 27520 11942 28000
rect 12530 27520 12586 28000
rect 13082 27520 13138 28000
rect 13634 27520 13690 28000
rect 14278 27520 14334 28000
rect 14830 27520 14886 28000
rect 15382 27520 15438 28000
rect 16026 27520 16082 28000
rect 16578 27520 16634 28000
rect 17130 27520 17186 28000
rect 17774 27520 17830 28000
rect 18326 27520 18382 28000
rect 18878 27520 18934 28000
rect 19522 27520 19578 28000
rect 20074 27520 20130 28000
rect 20626 27520 20682 28000
rect 21270 27520 21326 28000
rect 21822 27520 21878 28000
rect 22374 27520 22430 28000
rect 23018 27520 23074 28000
rect 23570 27520 23626 28000
rect 23754 27704 23810 27713
rect 23754 27639 23810 27648
rect 1306 26616 1362 26625
rect 1306 26551 1362 26560
rect 1124 24336 1176 24342
rect 1124 24278 1176 24284
rect 1032 22092 1084 22098
rect 1032 22034 1084 22040
rect 1136 22030 1164 24278
rect 1214 24168 1270 24177
rect 1214 24103 1270 24112
rect 1124 22024 1176 22030
rect 1124 21966 1176 21972
rect 1136 21146 1164 21966
rect 1124 21140 1176 21146
rect 1124 21082 1176 21088
rect 1228 20602 1256 24103
rect 1320 21690 1348 26551
rect 1412 25514 1440 27520
rect 1412 25486 1716 25514
rect 1492 25424 1544 25430
rect 1492 25366 1544 25372
rect 1400 24608 1452 24614
rect 1400 24550 1452 24556
rect 1308 21684 1360 21690
rect 1308 21626 1360 21632
rect 1216 20596 1268 20602
rect 1216 20538 1268 20544
rect 940 20052 992 20058
rect 940 19994 992 20000
rect 1412 19009 1440 24550
rect 1504 22438 1532 25366
rect 1584 24744 1636 24750
rect 1584 24686 1636 24692
rect 1596 23322 1624 24686
rect 1584 23316 1636 23322
rect 1584 23258 1636 23264
rect 1492 22432 1544 22438
rect 1492 22374 1544 22380
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1492 22092 1544 22098
rect 1492 22034 1544 22040
rect 1504 21010 1532 22034
rect 1492 21004 1544 21010
rect 1492 20946 1544 20952
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1398 19000 1454 19009
rect 1398 18935 1454 18944
rect 1504 17490 1532 19654
rect 1596 18834 1624 22374
rect 1584 18828 1636 18834
rect 1584 18770 1636 18776
rect 1582 18320 1638 18329
rect 1582 18255 1638 18264
rect 1596 17882 1624 18255
rect 1584 17876 1636 17882
rect 1584 17818 1636 17824
rect 1320 17462 1532 17490
rect 1320 17202 1348 17462
rect 1688 17354 1716 25486
rect 2056 25242 2084 27520
rect 2136 25356 2188 25362
rect 2136 25298 2188 25304
rect 2504 25356 2556 25362
rect 2504 25298 2556 25304
rect 1780 25214 2084 25242
rect 1780 19514 1808 25214
rect 2044 25152 2096 25158
rect 2044 25094 2096 25100
rect 1860 24268 1912 24274
rect 1860 24210 1912 24216
rect 1872 23338 1900 24210
rect 1952 24200 2004 24206
rect 1952 24142 2004 24148
rect 1964 23769 1992 24142
rect 1950 23760 2006 23769
rect 2056 23730 2084 25094
rect 2148 24614 2176 25298
rect 2228 25288 2280 25294
rect 2228 25230 2280 25236
rect 2136 24608 2188 24614
rect 2134 24576 2136 24585
rect 2188 24576 2190 24585
rect 2134 24511 2190 24520
rect 2240 24426 2268 25230
rect 2320 25152 2372 25158
rect 2320 25094 2372 25100
rect 2148 24398 2268 24426
rect 2148 24206 2176 24398
rect 2226 24304 2282 24313
rect 2226 24239 2228 24248
rect 2280 24239 2282 24248
rect 2228 24210 2280 24216
rect 2136 24200 2188 24206
rect 2136 24142 2188 24148
rect 2228 24064 2280 24070
rect 2228 24006 2280 24012
rect 1950 23695 2006 23704
rect 2044 23724 2096 23730
rect 2044 23666 2096 23672
rect 2056 23610 2084 23666
rect 2056 23582 2176 23610
rect 1952 23520 2004 23526
rect 2004 23480 2084 23508
rect 1952 23462 2004 23468
rect 1872 23310 1992 23338
rect 1860 22976 1912 22982
rect 1860 22918 1912 22924
rect 1872 22234 1900 22918
rect 1860 22228 1912 22234
rect 1860 22170 1912 22176
rect 1858 22128 1914 22137
rect 1858 22063 1914 22072
rect 1872 21690 1900 22063
rect 1964 21962 1992 23310
rect 1952 21956 2004 21962
rect 1952 21898 2004 21904
rect 1860 21684 1912 21690
rect 1860 21626 1912 21632
rect 2056 21434 2084 23480
rect 1872 21406 2084 21434
rect 1768 19508 1820 19514
rect 1768 19450 1820 19456
rect 1412 17326 1716 17354
rect 1308 17196 1360 17202
rect 1308 17138 1360 17144
rect 1308 16992 1360 16998
rect 1308 16934 1360 16940
rect 848 12368 900 12374
rect 18 12336 74 12345
rect 848 12310 900 12316
rect 18 12271 74 12280
rect 1320 11286 1348 16934
rect 1412 12102 1440 17326
rect 1872 17270 1900 21406
rect 2044 21344 2096 21350
rect 2044 21286 2096 21292
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 1964 18630 1992 19110
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 1964 18222 1992 18566
rect 1952 18216 2004 18222
rect 1952 18158 2004 18164
rect 1584 17264 1636 17270
rect 1584 17206 1636 17212
rect 1860 17264 1912 17270
rect 1860 17206 1912 17212
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 1504 15026 1532 17138
rect 1596 15502 1624 17206
rect 1964 17202 1992 18158
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 1950 17096 2006 17105
rect 1860 17060 1912 17066
rect 1950 17031 2006 17040
rect 1860 17002 1912 17008
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1584 15360 1636 15366
rect 1688 15337 1716 16594
rect 1766 16144 1822 16153
rect 1766 16079 1822 16088
rect 1780 15910 1808 16079
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1584 15302 1636 15308
rect 1674 15328 1730 15337
rect 1596 15065 1624 15302
rect 1674 15263 1730 15272
rect 1582 15056 1638 15065
rect 1492 15020 1544 15026
rect 1582 14991 1638 15000
rect 1492 14962 1544 14968
rect 1582 14920 1638 14929
rect 1582 14855 1638 14864
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1400 12096 1452 12102
rect 1400 12038 1452 12044
rect 1412 11694 1440 12038
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1308 11280 1360 11286
rect 1308 11222 1360 11228
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10033 1440 11086
rect 1504 10985 1532 14758
rect 1490 10976 1546 10985
rect 1490 10911 1546 10920
rect 1596 10810 1624 14855
rect 1688 13190 1716 15263
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1780 14482 1808 14962
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1872 14414 1900 17002
rect 1964 14958 1992 17031
rect 2056 16998 2084 21286
rect 2148 20602 2176 23582
rect 2136 20596 2188 20602
rect 2136 20538 2188 20544
rect 2136 19508 2188 19514
rect 2136 19450 2188 19456
rect 2148 17377 2176 19450
rect 2134 17368 2190 17377
rect 2134 17303 2190 17312
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 2044 16992 2096 16998
rect 2044 16934 2096 16940
rect 2148 16726 2176 17070
rect 2136 16720 2188 16726
rect 2136 16662 2188 16668
rect 2042 16552 2098 16561
rect 2042 16487 2098 16496
rect 2056 16250 2084 16487
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 1952 14952 2004 14958
rect 1952 14894 2004 14900
rect 1964 14618 1992 14894
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1952 14476 2004 14482
rect 1952 14418 2004 14424
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1780 12866 1808 14214
rect 1964 13938 1992 14418
rect 2056 14074 2084 15438
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 1952 13796 2004 13802
rect 1952 13738 2004 13744
rect 1860 13728 1912 13734
rect 1860 13670 1912 13676
rect 1872 13530 1900 13670
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1872 12986 1900 13262
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1780 12838 1900 12866
rect 1766 12336 1822 12345
rect 1766 12271 1768 12280
rect 1820 12271 1822 12280
rect 1768 12242 1820 12248
rect 1872 11665 1900 12838
rect 1964 12073 1992 13738
rect 2056 13462 2084 13874
rect 2044 13456 2096 13462
rect 2044 13398 2096 13404
rect 2148 13326 2176 16186
rect 2240 13802 2268 24006
rect 2332 23594 2360 25094
rect 2412 24744 2464 24750
rect 2410 24712 2412 24721
rect 2464 24712 2466 24721
rect 2410 24647 2466 24656
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2320 23588 2372 23594
rect 2320 23530 2372 23536
rect 2332 21146 2360 23530
rect 2320 21140 2372 21146
rect 2320 21082 2372 21088
rect 2424 20777 2452 24550
rect 2516 24070 2544 25298
rect 2504 24064 2556 24070
rect 2504 24006 2556 24012
rect 2516 21026 2544 24006
rect 2608 21350 2636 27520
rect 2688 26104 2740 26110
rect 2688 26046 2740 26052
rect 2596 21344 2648 21350
rect 2596 21286 2648 21292
rect 2516 20998 2636 21026
rect 2410 20768 2466 20777
rect 2410 20703 2466 20712
rect 2412 20460 2464 20466
rect 2412 20402 2464 20408
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 2424 20369 2452 20402
rect 2410 20360 2466 20369
rect 2410 20295 2466 20304
rect 2320 20256 2372 20262
rect 2320 20198 2372 20204
rect 2332 20058 2360 20198
rect 2320 20052 2372 20058
rect 2320 19994 2372 20000
rect 2516 19242 2544 20402
rect 2504 19236 2556 19242
rect 2504 19178 2556 19184
rect 2608 18986 2636 20998
rect 2516 18958 2636 18986
rect 2516 18902 2544 18958
rect 2504 18896 2556 18902
rect 2504 18838 2556 18844
rect 2596 18896 2648 18902
rect 2596 18838 2648 18844
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2320 17536 2372 17542
rect 2320 17478 2372 17484
rect 2332 15026 2360 17478
rect 2424 16697 2452 18770
rect 2504 18692 2556 18698
rect 2504 18634 2556 18640
rect 2516 17610 2544 18634
rect 2608 17882 2636 18838
rect 2596 17876 2648 17882
rect 2596 17818 2648 17824
rect 2504 17604 2556 17610
rect 2504 17546 2556 17552
rect 2502 17504 2558 17513
rect 2502 17439 2558 17448
rect 2410 16688 2466 16697
rect 2410 16623 2466 16632
rect 2412 16448 2464 16454
rect 2410 16416 2412 16425
rect 2464 16416 2466 16425
rect 2410 16351 2466 16360
rect 2424 15570 2452 16351
rect 2516 16114 2544 17439
rect 2700 17218 2728 26046
rect 2778 25392 2834 25401
rect 2778 25327 2834 25336
rect 2792 23186 2820 25327
rect 3160 25242 3188 27520
rect 3160 25214 3280 25242
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 3148 25152 3200 25158
rect 3148 25094 3200 25100
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2792 22642 2820 23122
rect 2780 22636 2832 22642
rect 2780 22578 2832 22584
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 2792 21554 2820 21966
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2792 21010 2820 21490
rect 2884 21321 2912 25094
rect 3056 24608 3108 24614
rect 3056 24550 3108 24556
rect 2964 24200 3016 24206
rect 2964 24142 3016 24148
rect 2976 23594 3004 24142
rect 2964 23588 3016 23594
rect 2964 23530 3016 23536
rect 2976 22166 3004 23530
rect 3068 23322 3096 24550
rect 3160 23866 3188 25094
rect 3252 24721 3280 25214
rect 3424 25152 3476 25158
rect 3424 25094 3476 25100
rect 3700 25152 3752 25158
rect 3700 25094 3752 25100
rect 3436 24886 3464 25094
rect 3424 24880 3476 24886
rect 3424 24822 3476 24828
rect 3238 24712 3294 24721
rect 3238 24647 3294 24656
rect 3148 23860 3200 23866
rect 3148 23802 3200 23808
rect 3056 23316 3108 23322
rect 3056 23258 3108 23264
rect 3056 22704 3108 22710
rect 3056 22646 3108 22652
rect 2964 22160 3016 22166
rect 2964 22102 3016 22108
rect 2870 21312 2926 21321
rect 2870 21247 2926 21256
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 2792 20466 2820 20946
rect 2872 20868 2924 20874
rect 2872 20810 2924 20816
rect 2884 20534 2912 20810
rect 2872 20528 2924 20534
rect 2872 20470 2924 20476
rect 2780 20460 2832 20466
rect 2780 20402 2832 20408
rect 2870 20224 2926 20233
rect 2870 20159 2926 20168
rect 2884 19990 2912 20159
rect 2872 19984 2924 19990
rect 3068 19938 3096 22646
rect 3160 22642 3188 23802
rect 3240 23180 3292 23186
rect 3240 23122 3292 23128
rect 3148 22636 3200 22642
rect 3148 22578 3200 22584
rect 3148 22500 3200 22506
rect 3148 22442 3200 22448
rect 3160 21146 3188 22442
rect 3252 22098 3280 23122
rect 3332 22636 3384 22642
rect 3332 22578 3384 22584
rect 3344 22438 3372 22578
rect 3436 22574 3464 24822
rect 3516 23248 3568 23254
rect 3516 23190 3568 23196
rect 3528 23089 3556 23190
rect 3514 23080 3570 23089
rect 3514 23015 3516 23024
rect 3568 23015 3570 23024
rect 3516 22986 3568 22992
rect 3424 22568 3476 22574
rect 3424 22510 3476 22516
rect 3332 22432 3384 22438
rect 3330 22400 3332 22409
rect 3384 22400 3386 22409
rect 3330 22335 3386 22344
rect 3344 22309 3372 22335
rect 3240 22092 3292 22098
rect 3240 22034 3292 22040
rect 3608 22024 3660 22030
rect 3608 21966 3660 21972
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 3516 21888 3568 21894
rect 3516 21830 3568 21836
rect 3252 21593 3280 21830
rect 3422 21720 3478 21729
rect 3422 21655 3478 21664
rect 3436 21622 3464 21655
rect 3424 21616 3476 21622
rect 3238 21584 3294 21593
rect 3424 21558 3476 21564
rect 3528 21554 3556 21830
rect 3238 21519 3294 21528
rect 3516 21548 3568 21554
rect 3516 21490 3568 21496
rect 3422 21448 3478 21457
rect 3422 21383 3478 21392
rect 3148 21140 3200 21146
rect 3148 21082 3200 21088
rect 3160 20874 3188 21082
rect 3332 21072 3384 21078
rect 3238 21040 3294 21049
rect 3332 21014 3384 21020
rect 3238 20975 3294 20984
rect 3148 20868 3200 20874
rect 3148 20810 3200 20816
rect 3160 20602 3188 20810
rect 3148 20596 3200 20602
rect 3148 20538 3200 20544
rect 2872 19926 2924 19932
rect 2976 19910 3096 19938
rect 2778 19000 2834 19009
rect 2778 18935 2780 18944
rect 2832 18935 2834 18944
rect 2780 18906 2832 18912
rect 2792 18442 2820 18906
rect 2792 18426 2912 18442
rect 2792 18420 2924 18426
rect 2792 18414 2872 18420
rect 2872 18362 2924 18368
rect 2780 17808 2832 17814
rect 2780 17750 2832 17756
rect 2792 17338 2820 17750
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2608 17190 2728 17218
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2516 15706 2544 16050
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2424 15201 2452 15302
rect 2410 15192 2466 15201
rect 2410 15127 2466 15136
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2516 14822 2544 15438
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2410 14648 2466 14657
rect 2410 14583 2412 14592
rect 2464 14583 2466 14592
rect 2412 14554 2464 14560
rect 2228 13796 2280 13802
rect 2228 13738 2280 13744
rect 2424 13530 2452 14554
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2042 13152 2098 13161
rect 2042 13087 2098 13096
rect 2056 12986 2084 13087
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 2136 12912 2188 12918
rect 2136 12854 2188 12860
rect 2148 12442 2176 12854
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 1950 12064 2006 12073
rect 1950 11999 2006 12008
rect 1952 11688 2004 11694
rect 1858 11656 1914 11665
rect 1952 11630 2004 11636
rect 1858 11591 1914 11600
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1780 10146 1808 11494
rect 1964 11354 1992 11630
rect 2056 11354 2084 12310
rect 2240 11801 2268 13466
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2424 12481 2452 12582
rect 2410 12472 2466 12481
rect 2410 12407 2466 12416
rect 2608 12356 2636 17190
rect 2778 16960 2834 16969
rect 2778 16895 2834 16904
rect 2792 16794 2820 16895
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2780 16584 2832 16590
rect 2700 16544 2780 16572
rect 2700 15978 2728 16544
rect 2780 16526 2832 16532
rect 2780 16448 2832 16454
rect 2884 16436 2912 17614
rect 2976 17241 3004 19910
rect 3056 19848 3108 19854
rect 3056 19790 3108 19796
rect 3068 19378 3096 19790
rect 3252 19394 3280 20975
rect 3344 20398 3372 21014
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3056 19372 3108 19378
rect 3252 19366 3372 19394
rect 3056 19314 3108 19320
rect 3240 19236 3292 19242
rect 3240 19178 3292 19184
rect 3252 18630 3280 19178
rect 3344 18902 3372 19366
rect 3332 18896 3384 18902
rect 3332 18838 3384 18844
rect 3056 18624 3108 18630
rect 3056 18566 3108 18572
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3068 17746 3096 18566
rect 3056 17740 3108 17746
rect 3056 17682 3108 17688
rect 3252 17678 3280 18566
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 2962 17232 3018 17241
rect 2962 17167 3018 17176
rect 3252 16794 3280 17614
rect 3344 17066 3372 18022
rect 3436 17814 3464 21383
rect 3516 21344 3568 21350
rect 3516 21286 3568 21292
rect 3528 20806 3556 21286
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 3528 20505 3556 20742
rect 3514 20496 3570 20505
rect 3514 20431 3570 20440
rect 3516 20324 3568 20330
rect 3516 20266 3568 20272
rect 3528 19990 3556 20266
rect 3516 19984 3568 19990
rect 3516 19926 3568 19932
rect 3620 19174 3648 21966
rect 3712 21865 3740 25094
rect 3804 24857 3832 27520
rect 4356 25514 4384 27520
rect 4356 25486 4660 25514
rect 4068 25356 4120 25362
rect 4068 25298 4120 25304
rect 3790 24848 3846 24857
rect 3790 24783 3846 24792
rect 4080 24614 4108 25298
rect 4344 25220 4396 25226
rect 4344 25162 4396 25168
rect 3792 24608 3844 24614
rect 3792 24550 3844 24556
rect 4068 24608 4120 24614
rect 4068 24550 4120 24556
rect 3804 22438 3832 24550
rect 4356 24154 4384 25162
rect 3884 24132 3936 24138
rect 3884 24074 3936 24080
rect 4172 24126 4384 24154
rect 3896 23769 3924 24074
rect 4068 24064 4120 24070
rect 4068 24006 4120 24012
rect 3882 23760 3938 23769
rect 4080 23730 4108 24006
rect 3882 23695 3938 23704
rect 4068 23724 4120 23730
rect 3896 23662 3924 23695
rect 4068 23666 4120 23672
rect 3884 23656 3936 23662
rect 3884 23598 3936 23604
rect 3974 23624 4030 23633
rect 3974 23559 4030 23568
rect 3884 22772 3936 22778
rect 3884 22714 3936 22720
rect 3792 22432 3844 22438
rect 3792 22374 3844 22380
rect 3792 21888 3844 21894
rect 3698 21856 3754 21865
rect 3792 21830 3844 21836
rect 3698 21791 3754 21800
rect 3700 20528 3752 20534
rect 3700 20470 3752 20476
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3620 18154 3648 19110
rect 3608 18148 3660 18154
rect 3608 18090 3660 18096
rect 3620 17814 3648 18090
rect 3424 17808 3476 17814
rect 3424 17750 3476 17756
rect 3608 17808 3660 17814
rect 3608 17750 3660 17756
rect 3712 17762 3740 20470
rect 3804 19922 3832 21830
rect 3896 21622 3924 22714
rect 3884 21616 3936 21622
rect 3884 21558 3936 21564
rect 3792 19916 3844 19922
rect 3792 19858 3844 19864
rect 3988 18714 4016 23559
rect 4066 23488 4122 23497
rect 4066 23423 4122 23432
rect 4080 22545 4108 23423
rect 4172 23066 4200 24126
rect 4344 24064 4396 24070
rect 4344 24006 4396 24012
rect 4250 23896 4306 23905
rect 4250 23831 4306 23840
rect 4264 23633 4292 23831
rect 4250 23624 4306 23633
rect 4250 23559 4306 23568
rect 4172 23038 4292 23066
rect 4160 22976 4212 22982
rect 4160 22918 4212 22924
rect 4066 22536 4122 22545
rect 4066 22471 4122 22480
rect 4068 22228 4120 22234
rect 4068 22170 4120 22176
rect 4080 21146 4108 22170
rect 4172 22030 4200 22918
rect 4264 22794 4292 23038
rect 4356 22953 4384 24006
rect 4528 23724 4580 23730
rect 4528 23666 4580 23672
rect 4342 22944 4398 22953
rect 4342 22879 4398 22888
rect 4264 22766 4476 22794
rect 4342 22672 4398 22681
rect 4342 22607 4398 22616
rect 4356 22234 4384 22607
rect 4344 22228 4396 22234
rect 4344 22170 4396 22176
rect 4160 22024 4212 22030
rect 4160 21966 4212 21972
rect 4068 21140 4120 21146
rect 4068 21082 4120 21088
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 4172 19990 4200 20946
rect 4344 20256 4396 20262
rect 4344 20198 4396 20204
rect 4160 19984 4212 19990
rect 4160 19926 4212 19932
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 3896 18686 4016 18714
rect 3332 17060 3384 17066
rect 3332 17002 3384 17008
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 3054 16688 3110 16697
rect 3054 16623 3110 16632
rect 2884 16408 3004 16436
rect 2780 16390 2832 16396
rect 2792 16114 2820 16390
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 2700 15162 2728 15506
rect 2792 15434 2820 16050
rect 2780 15428 2832 15434
rect 2780 15370 2832 15376
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 2780 15088 2832 15094
rect 2780 15030 2832 15036
rect 2792 14618 2820 15030
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2700 14074 2728 14350
rect 2792 14074 2820 14418
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2700 13394 2728 13806
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2792 12986 2820 14010
rect 2884 13308 2912 14758
rect 2976 13462 3004 16408
rect 3068 14618 3096 16623
rect 3146 16552 3202 16561
rect 3146 16487 3202 16496
rect 3160 15881 3188 16487
rect 3436 16250 3464 16934
rect 3516 16516 3568 16522
rect 3516 16458 3568 16464
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3332 15904 3384 15910
rect 3146 15872 3202 15881
rect 3332 15846 3384 15852
rect 3146 15807 3202 15816
rect 3160 14958 3188 15807
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 3344 13852 3372 15846
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 3252 13824 3372 13852
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3160 13530 3188 13670
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 2964 13456 3016 13462
rect 2964 13398 3016 13404
rect 2884 13280 3004 13308
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2516 12328 2636 12356
rect 2700 12345 2728 12582
rect 2686 12336 2742 12345
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2410 12200 2466 12209
rect 2226 11792 2282 11801
rect 2226 11727 2282 11736
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 1860 11280 1912 11286
rect 2056 11257 2084 11290
rect 1860 11222 1912 11228
rect 2042 11248 2098 11257
rect 1872 10266 1900 11222
rect 2042 11183 2098 11192
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 2042 10568 2098 10577
rect 2042 10503 2044 10512
rect 2096 10503 2098 10512
rect 2044 10474 2096 10480
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1596 10118 1808 10146
rect 1398 10024 1454 10033
rect 1398 9959 1454 9968
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 1412 5846 1440 9551
rect 1596 9382 1624 10118
rect 1768 9648 1820 9654
rect 1766 9616 1768 9625
rect 1820 9616 1822 9625
rect 1766 9551 1822 9560
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 8786 1624 9318
rect 1504 8758 1624 8786
rect 1400 5840 1452 5846
rect 1400 5782 1452 5788
rect 662 3088 718 3097
rect 662 3023 718 3032
rect 202 1728 258 1737
rect 202 1663 258 1672
rect 216 480 244 1663
rect 676 480 704 3023
rect 1216 2848 1268 2854
rect 1216 2790 1268 2796
rect 1228 480 1256 2790
rect 1504 785 1532 8758
rect 1780 8498 1808 9551
rect 2148 9489 2176 11018
rect 2332 10305 2360 12174
rect 2410 12135 2412 12144
rect 2464 12135 2466 12144
rect 2412 12106 2464 12112
rect 2424 11694 2452 12106
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2318 10296 2374 10305
rect 2318 10231 2374 10240
rect 2134 9480 2190 9489
rect 2134 9415 2136 9424
rect 2188 9415 2190 9424
rect 2136 9386 2188 9392
rect 2148 9355 2176 9386
rect 2042 9344 2098 9353
rect 2042 9279 2098 9288
rect 1950 8800 2006 8809
rect 1950 8735 2006 8744
rect 1858 8528 1914 8537
rect 1768 8492 1820 8498
rect 1858 8463 1914 8472
rect 1768 8434 1820 8440
rect 1872 8430 1900 8463
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1964 7342 1992 8735
rect 2056 8634 2084 9279
rect 2410 9208 2466 9217
rect 2410 9143 2412 9152
rect 2464 9143 2466 9152
rect 2412 9114 2464 9120
rect 2134 9072 2190 9081
rect 2134 9007 2190 9016
rect 2228 9036 2280 9042
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2042 7440 2098 7449
rect 2042 7375 2044 7384
rect 2096 7375 2098 7384
rect 2044 7346 2096 7352
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 7041 1624 7142
rect 1582 7032 1638 7041
rect 1964 7002 1992 7278
rect 1582 6967 1638 6976
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1858 6216 1914 6225
rect 1858 6151 1914 6160
rect 1872 5574 1900 6151
rect 2148 5914 2176 9007
rect 2228 8978 2280 8984
rect 2240 8090 2268 8978
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2240 6322 2268 7346
rect 2332 6934 2360 8570
rect 2424 8090 2452 9114
rect 2516 8276 2544 12328
rect 2686 12271 2742 12280
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2608 11898 2636 12174
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2870 11520 2926 11529
rect 2870 11455 2926 11464
rect 2884 11354 2912 11455
rect 2872 11348 2924 11354
rect 2700 11308 2872 11336
rect 2700 10266 2728 11308
rect 2872 11290 2924 11296
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2608 8344 2636 9862
rect 2700 9518 2728 10066
rect 2792 9586 2820 10474
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2884 9722 2912 10202
rect 2976 9994 3004 13280
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3160 11898 3188 12242
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3160 11150 3188 11834
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3160 10198 3188 11086
rect 3252 10538 3280 13824
rect 3436 12322 3464 15642
rect 3344 12294 3464 12322
rect 3240 10532 3292 10538
rect 3240 10474 3292 10480
rect 3344 10266 3372 12294
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3436 11354 3464 12174
rect 3528 11898 3556 16458
rect 3620 15026 3648 17750
rect 3712 17734 3832 17762
rect 3698 17640 3754 17649
rect 3698 17575 3754 17584
rect 3712 16046 3740 17575
rect 3804 17338 3832 17734
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 3896 17270 3924 18686
rect 3976 18624 4028 18630
rect 3976 18566 4028 18572
rect 3884 17264 3936 17270
rect 3884 17206 3936 17212
rect 3792 17060 3844 17066
rect 3792 17002 3844 17008
rect 3804 16794 3832 17002
rect 3792 16788 3844 16794
rect 3792 16730 3844 16736
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 3804 16182 3832 16594
rect 3792 16176 3844 16182
rect 3790 16144 3792 16153
rect 3844 16144 3846 16153
rect 3790 16079 3846 16088
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 3700 16040 3752 16046
rect 3700 15982 3752 15988
rect 3896 15706 3924 16050
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 3988 15473 4016 18566
rect 4080 18329 4108 19858
rect 4160 19780 4212 19786
rect 4160 19722 4212 19728
rect 4172 19242 4200 19722
rect 4356 19718 4384 20198
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 4160 19236 4212 19242
rect 4160 19178 4212 19184
rect 4158 18864 4214 18873
rect 4158 18799 4160 18808
rect 4212 18799 4214 18808
rect 4160 18770 4212 18776
rect 4172 18426 4200 18770
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4066 18320 4122 18329
rect 4066 18255 4122 18264
rect 4172 17513 4200 18362
rect 4158 17504 4214 17513
rect 4158 17439 4214 17448
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4172 16794 4200 16934
rect 4264 16833 4292 19654
rect 4344 18352 4396 18358
rect 4342 18320 4344 18329
rect 4396 18320 4398 18329
rect 4342 18255 4398 18264
rect 4344 17264 4396 17270
rect 4344 17206 4396 17212
rect 4250 16824 4306 16833
rect 4160 16788 4212 16794
rect 4250 16759 4306 16768
rect 4160 16730 4212 16736
rect 4066 16688 4122 16697
rect 4356 16640 4384 17206
rect 4066 16623 4122 16632
rect 4080 16017 4108 16623
rect 4172 16612 4384 16640
rect 4066 16008 4122 16017
rect 4066 15943 4122 15952
rect 4172 15858 4200 16612
rect 4080 15830 4200 15858
rect 4080 15638 4108 15830
rect 4068 15632 4120 15638
rect 4068 15574 4120 15580
rect 3974 15464 4030 15473
rect 3974 15399 4030 15408
rect 3700 15360 3752 15366
rect 3700 15302 3752 15308
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 3620 14346 3648 14962
rect 3712 14822 3740 15302
rect 3790 15192 3846 15201
rect 3790 15127 3846 15136
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3608 14340 3660 14346
rect 3608 14282 3660 14288
rect 3620 14006 3648 14282
rect 3608 14000 3660 14006
rect 3608 13942 3660 13948
rect 3804 13734 3832 15127
rect 3988 15094 4016 15302
rect 3976 15088 4028 15094
rect 3976 15030 4028 15036
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3804 13569 3832 13670
rect 3790 13560 3846 13569
rect 3790 13495 3846 13504
rect 3790 13424 3846 13433
rect 3790 13359 3846 13368
rect 3804 12782 3832 13359
rect 4080 13326 4108 15574
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 4250 14920 4306 14929
rect 4356 14890 4384 15506
rect 4250 14855 4252 14864
rect 4304 14855 4306 14864
rect 4344 14884 4396 14890
rect 4252 14826 4304 14832
rect 4344 14826 4396 14832
rect 4264 14618 4292 14826
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 4172 13258 4200 14418
rect 4252 14408 4304 14414
rect 4356 14396 4384 14826
rect 4304 14368 4384 14396
rect 4252 14350 4304 14356
rect 4250 13696 4306 13705
rect 4250 13631 4306 13640
rect 4160 13252 4212 13258
rect 4160 13194 4212 13200
rect 4172 13138 4200 13194
rect 3896 13110 4200 13138
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3698 12608 3754 12617
rect 3620 12481 3648 12582
rect 3698 12543 3754 12552
rect 3606 12472 3662 12481
rect 3606 12407 3662 12416
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3606 11656 3662 11665
rect 3606 11591 3662 11600
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3514 10976 3570 10985
rect 3514 10911 3570 10920
rect 3528 10441 3556 10911
rect 3514 10432 3570 10441
rect 3514 10367 3570 10376
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3148 10192 3200 10198
rect 3148 10134 3200 10140
rect 3160 10062 3188 10134
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2872 8968 2924 8974
rect 2870 8936 2872 8945
rect 2924 8936 2926 8945
rect 2870 8871 2926 8880
rect 2884 8566 2912 8871
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2608 8316 2820 8344
rect 2516 8248 2728 8276
rect 2502 8120 2558 8129
rect 2412 8084 2464 8090
rect 2502 8055 2558 8064
rect 2412 8026 2464 8032
rect 2412 7744 2464 7750
rect 2410 7712 2412 7721
rect 2464 7712 2466 7721
rect 2410 7647 2466 7656
rect 2320 6928 2372 6934
rect 2320 6870 2372 6876
rect 2410 6760 2466 6769
rect 2410 6695 2412 6704
rect 2464 6695 2466 6704
rect 2412 6666 2464 6672
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2332 6322 2360 6598
rect 2516 6458 2544 8055
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2136 5908 2188 5914
rect 2056 5868 2136 5896
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1780 5234 1808 5510
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1872 4457 1900 5510
rect 2056 5166 2084 5868
rect 2136 5850 2188 5856
rect 2136 5296 2188 5302
rect 2136 5238 2188 5244
rect 2318 5264 2374 5273
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 1858 4448 1914 4457
rect 1858 4383 1914 4392
rect 2148 4078 2176 5238
rect 2318 5199 2374 5208
rect 2332 4826 2360 5199
rect 2516 5166 2544 6394
rect 2596 6248 2648 6254
rect 2594 6216 2596 6225
rect 2648 6216 2650 6225
rect 2594 6151 2650 6160
rect 2700 6089 2728 8248
rect 2792 7206 2820 8316
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 8022 3004 8230
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2976 7857 3004 7958
rect 3068 7886 3096 9658
rect 3160 9450 3188 9998
rect 3332 9988 3384 9994
rect 3332 9930 3384 9936
rect 3238 9752 3294 9761
rect 3238 9687 3294 9696
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 3160 8974 3188 9386
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3146 8528 3202 8537
rect 3146 8463 3202 8472
rect 3056 7880 3108 7886
rect 2962 7848 3018 7857
rect 3056 7822 3108 7828
rect 2962 7783 3018 7792
rect 3068 7478 3096 7822
rect 3160 7546 3188 8463
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3056 7472 3108 7478
rect 3056 7414 3108 7420
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 3148 6928 3200 6934
rect 3148 6870 3200 6876
rect 3056 6724 3108 6730
rect 2884 6684 3056 6712
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2686 6080 2742 6089
rect 2686 6015 2742 6024
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2700 5302 2728 5578
rect 2688 5296 2740 5302
rect 2688 5238 2740 5244
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 2792 4842 2820 6598
rect 2700 4826 2820 4842
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2688 4820 2820 4826
rect 2740 4814 2820 4820
rect 2688 4762 2740 4768
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2332 4214 2360 4626
rect 2320 4208 2372 4214
rect 2226 4176 2282 4185
rect 2320 4150 2372 4156
rect 2226 4111 2282 4120
rect 2136 4072 2188 4078
rect 2136 4014 2188 4020
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 2056 3194 2084 3538
rect 2240 3534 2268 4111
rect 2332 3670 2360 4150
rect 2700 4078 2728 4762
rect 2778 4720 2834 4729
rect 2778 4655 2834 4664
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 2320 3664 2372 3670
rect 2320 3606 2372 3612
rect 2228 3528 2280 3534
rect 2516 3482 2544 3946
rect 2688 3936 2740 3942
rect 2228 3470 2280 3476
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 1768 3120 1820 3126
rect 1768 3062 1820 3068
rect 1584 2304 1636 2310
rect 1582 2272 1584 2281
rect 1636 2272 1638 2281
rect 1582 2207 1638 2216
rect 1490 776 1546 785
rect 1490 711 1546 720
rect 1780 480 1808 3062
rect 2240 2650 2268 3470
rect 2332 3454 2544 3482
rect 2608 3896 2688 3924
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 1964 2310 1992 2450
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 1964 1873 1992 2246
rect 1950 1864 2006 1873
rect 1950 1799 2006 1808
rect 2332 480 2360 3454
rect 2608 3346 2636 3896
rect 2792 3924 2820 4655
rect 2740 3896 2820 3924
rect 2688 3878 2740 3884
rect 2884 3754 2912 6684
rect 3056 6666 3108 6672
rect 3160 6118 3188 6870
rect 3252 6798 3280 9687
rect 3344 8673 3372 9930
rect 3422 9208 3478 9217
rect 3422 9143 3478 9152
rect 3330 8664 3386 8673
rect 3330 8599 3386 8608
rect 3330 8528 3386 8537
rect 3330 8463 3386 8472
rect 3344 8430 3372 8463
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3252 6458 3280 6734
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2976 5370 3004 5850
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 3068 5273 3096 5714
rect 3054 5264 3110 5273
rect 3054 5199 3110 5208
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2976 4282 3004 4558
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2700 3738 2912 3754
rect 2688 3732 2912 3738
rect 2740 3726 2912 3732
rect 2688 3674 2740 3680
rect 2608 3318 2820 3346
rect 2688 3120 2740 3126
rect 2688 3062 2740 3068
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 2516 1329 2544 2926
rect 2700 2922 2728 3062
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 2792 2582 2820 3318
rect 2884 2650 2912 3726
rect 2976 3058 3004 4218
rect 3160 3233 3188 6054
rect 3252 5370 3280 6190
rect 3344 5914 3372 8366
rect 3436 7585 3464 9143
rect 3422 7576 3478 7585
rect 3422 7511 3478 7520
rect 3528 7290 3556 10367
rect 3620 7954 3648 11591
rect 3712 9625 3740 12543
rect 3790 12472 3846 12481
rect 3790 12407 3846 12416
rect 3804 12374 3832 12407
rect 3792 12368 3844 12374
rect 3792 12310 3844 12316
rect 3896 12238 3924 13110
rect 3974 13016 4030 13025
rect 3974 12951 4030 12960
rect 3884 12232 3936 12238
rect 3988 12209 4016 12951
rect 4066 12880 4122 12889
rect 4066 12815 4068 12824
rect 4120 12815 4122 12824
rect 4068 12786 4120 12792
rect 4066 12744 4122 12753
rect 4066 12679 4068 12688
rect 4120 12679 4122 12688
rect 4068 12650 4120 12656
rect 4264 12442 4292 13631
rect 4344 13456 4396 13462
rect 4344 13398 4396 13404
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4356 12322 4384 13398
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4264 12294 4384 12322
rect 3884 12174 3936 12180
rect 3974 12200 4030 12209
rect 3974 12135 4030 12144
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3896 11626 3924 12038
rect 3974 11928 4030 11937
rect 3974 11863 4030 11872
rect 3884 11620 3936 11626
rect 3884 11562 3936 11568
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10606 3832 10950
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3896 10470 3924 11562
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3698 9616 3754 9625
rect 3698 9551 3754 9560
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3790 8936 3846 8945
rect 3712 8498 3740 8910
rect 3790 8871 3846 8880
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3712 7886 3740 8298
rect 3700 7880 3752 7886
rect 3698 7848 3700 7857
rect 3752 7848 3754 7857
rect 3698 7783 3754 7792
rect 3528 7262 3648 7290
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3528 6905 3556 7142
rect 3514 6896 3570 6905
rect 3514 6831 3570 6840
rect 3422 5944 3478 5953
rect 3332 5908 3384 5914
rect 3422 5879 3478 5888
rect 3332 5850 3384 5856
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3252 5166 3280 5306
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 3252 4554 3280 5102
rect 3436 4690 3464 5879
rect 3620 5778 3648 7262
rect 3712 6934 3740 7783
rect 3804 7342 3832 8871
rect 3896 8294 3924 10406
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 7750 3924 8230
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3700 6928 3752 6934
rect 3700 6870 3752 6876
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3528 5166 3556 5646
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3240 4548 3292 4554
rect 3240 4490 3292 4496
rect 3436 4282 3464 4626
rect 3528 4622 3556 5102
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3146 3224 3202 3233
rect 3712 3194 3740 6598
rect 3988 5914 4016 11863
rect 4080 11354 4108 12242
rect 4264 11626 4292 12294
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4264 11218 4292 11562
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4264 10810 4292 11154
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 4080 8945 4108 9862
rect 4158 9616 4214 9625
rect 4158 9551 4214 9560
rect 4066 8936 4122 8945
rect 4066 8871 4122 8880
rect 4172 8090 4200 9551
rect 4264 9450 4292 10746
rect 4356 9994 4384 12174
rect 4344 9988 4396 9994
rect 4344 9930 4396 9936
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 4264 9042 4292 9386
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4066 7032 4122 7041
rect 4066 6967 4068 6976
rect 4120 6967 4122 6976
rect 4068 6938 4120 6944
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4080 5794 4108 6190
rect 3988 5766 4108 5794
rect 3988 5574 4016 5766
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3988 4486 4016 5510
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4080 4593 4108 4762
rect 4172 4729 4200 7142
rect 4264 6186 4292 8978
rect 4252 6180 4304 6186
rect 4252 6122 4304 6128
rect 4158 4720 4214 4729
rect 4158 4655 4214 4664
rect 4066 4584 4122 4593
rect 4066 4519 4122 4528
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3988 4146 4016 4422
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3882 4040 3938 4049
rect 3882 3975 3884 3984
rect 3936 3975 3938 3984
rect 3884 3946 3936 3952
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3804 3738 3832 3878
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3146 3159 3202 3168
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 2962 2952 3018 2961
rect 2962 2887 3018 2896
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 2502 1320 2558 1329
rect 2502 1255 2558 1264
rect 2976 1034 3004 2887
rect 3528 1034 3556 3062
rect 3804 2961 3832 3674
rect 3988 3534 4016 4082
rect 4080 3738 4108 4519
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 4172 3777 4200 3946
rect 4158 3768 4214 3777
rect 4068 3732 4120 3738
rect 4158 3703 4214 3712
rect 4068 3674 4120 3680
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3988 3058 4016 3470
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 3790 2952 3846 2961
rect 3790 2887 3846 2896
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3712 2582 3740 2790
rect 3700 2576 3752 2582
rect 3698 2544 3700 2553
rect 3752 2544 3754 2553
rect 3698 2479 3754 2488
rect 3712 2453 3740 2479
rect 4264 2446 4292 4422
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4066 2000 4122 2009
rect 4066 1935 4122 1944
rect 4080 1601 4108 1935
rect 4066 1592 4122 1601
rect 4066 1527 4122 1536
rect 4356 1465 4384 9522
rect 4448 7721 4476 22766
rect 4540 22574 4568 23666
rect 4528 22568 4580 22574
rect 4528 22510 4580 22516
rect 4540 22098 4568 22510
rect 4528 22092 4580 22098
rect 4528 22034 4580 22040
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4540 18970 4568 19246
rect 4528 18964 4580 18970
rect 4528 18906 4580 18912
rect 4528 17536 4580 17542
rect 4528 17478 4580 17484
rect 4540 11642 4568 17478
rect 4632 14958 4660 25486
rect 4712 25152 4764 25158
rect 4712 25094 4764 25100
rect 4724 24886 4752 25094
rect 4712 24880 4764 24886
rect 4712 24822 4764 24828
rect 4724 23730 4752 24822
rect 4802 24712 4858 24721
rect 4802 24647 4858 24656
rect 4712 23724 4764 23730
rect 4712 23666 4764 23672
rect 4712 22500 4764 22506
rect 4712 22442 4764 22448
rect 4724 22166 4752 22442
rect 4712 22160 4764 22166
rect 4712 22102 4764 22108
rect 4724 20398 4752 22102
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 4724 19922 4752 20334
rect 4712 19916 4764 19922
rect 4712 19858 4764 19864
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4632 12238 4660 14894
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4620 12096 4672 12102
rect 4618 12064 4620 12073
rect 4672 12064 4674 12073
rect 4618 11999 4674 12008
rect 4540 11614 4660 11642
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4540 11218 4568 11494
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4540 9761 4568 11154
rect 4632 10146 4660 11614
rect 4724 10606 4752 19654
rect 4816 17542 4844 24647
rect 4908 22137 4936 27520
rect 5172 26104 5224 26110
rect 5172 26046 5224 26052
rect 5080 25968 5132 25974
rect 5080 25910 5132 25916
rect 4988 25152 5040 25158
rect 4988 25094 5040 25100
rect 5000 24750 5028 25094
rect 4988 24744 5040 24750
rect 4988 24686 5040 24692
rect 5000 24410 5028 24686
rect 4988 24404 5040 24410
rect 4988 24346 5040 24352
rect 5092 24290 5120 25910
rect 5184 25226 5212 26046
rect 5552 25498 5580 27520
rect 5540 25492 5592 25498
rect 5540 25434 5592 25440
rect 5264 25424 5316 25430
rect 5264 25366 5316 25372
rect 5172 25220 5224 25226
rect 5172 25162 5224 25168
rect 5170 24848 5226 24857
rect 5170 24783 5226 24792
rect 5000 24262 5120 24290
rect 5000 22778 5028 24262
rect 5080 24200 5132 24206
rect 5080 24142 5132 24148
rect 5092 23254 5120 24142
rect 5080 23248 5132 23254
rect 5080 23190 5132 23196
rect 4988 22772 5040 22778
rect 4988 22714 5040 22720
rect 4894 22128 4950 22137
rect 4894 22063 4950 22072
rect 4896 22024 4948 22030
rect 4896 21966 4948 21972
rect 4988 22024 5040 22030
rect 4988 21966 5040 21972
rect 4908 21690 4936 21966
rect 4896 21684 4948 21690
rect 4896 21626 4948 21632
rect 5000 20806 5028 21966
rect 5080 21684 5132 21690
rect 5080 21626 5132 21632
rect 4988 20800 5040 20806
rect 4988 20742 5040 20748
rect 5000 20330 5028 20742
rect 4988 20324 5040 20330
rect 4988 20266 5040 20272
rect 5000 20058 5028 20266
rect 4988 20052 5040 20058
rect 4988 19994 5040 20000
rect 4988 19916 5040 19922
rect 4988 19858 5040 19864
rect 5000 19242 5028 19858
rect 4988 19236 5040 19242
rect 4988 19178 5040 19184
rect 5000 18834 5028 19178
rect 4988 18828 5040 18834
rect 4988 18770 5040 18776
rect 5092 17864 5120 21626
rect 5184 18170 5212 24783
rect 5276 24410 5304 25366
rect 5552 24868 5580 25434
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5460 24840 5580 24868
rect 5264 24404 5316 24410
rect 5264 24346 5316 24352
rect 5276 23322 5304 24346
rect 5460 23730 5488 24840
rect 6000 24608 6052 24614
rect 6000 24550 6052 24556
rect 5540 24268 5592 24274
rect 5540 24210 5592 24216
rect 5552 23866 5580 24210
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5448 23724 5500 23730
rect 5448 23666 5500 23672
rect 5632 23588 5684 23594
rect 5632 23530 5684 23536
rect 5264 23316 5316 23322
rect 5264 23258 5316 23264
rect 5644 23186 5672 23530
rect 6012 23186 6040 24550
rect 6104 24154 6132 27520
rect 6366 26072 6422 26081
rect 6366 26007 6422 26016
rect 6184 24336 6236 24342
rect 6182 24304 6184 24313
rect 6236 24304 6238 24313
rect 6182 24239 6238 24248
rect 6104 24126 6224 24154
rect 6380 24138 6408 26007
rect 6552 25356 6604 25362
rect 6552 25298 6604 25304
rect 6460 25152 6512 25158
rect 6460 25094 6512 25100
rect 6092 24064 6144 24070
rect 6092 24006 6144 24012
rect 6104 23730 6132 24006
rect 6092 23724 6144 23730
rect 6092 23666 6144 23672
rect 5448 23180 5500 23186
rect 5448 23122 5500 23128
rect 5632 23180 5684 23186
rect 5632 23122 5684 23128
rect 6000 23180 6052 23186
rect 6000 23122 6052 23128
rect 5356 22772 5408 22778
rect 5356 22714 5408 22720
rect 5264 22432 5316 22438
rect 5264 22374 5316 22380
rect 5276 20466 5304 22374
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5276 19310 5304 20198
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5276 18290 5304 18566
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5184 18142 5304 18170
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 17921 5212 18022
rect 4908 17836 5120 17864
rect 5170 17912 5226 17921
rect 5170 17847 5226 17856
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4816 15910 4844 16594
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4816 15570 4844 15846
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4802 14512 4858 14521
rect 4802 14447 4858 14456
rect 4816 13530 4844 14447
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4802 11656 4858 11665
rect 4802 11591 4804 11600
rect 4856 11591 4858 11600
rect 4804 11562 4856 11568
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4724 10266 4752 10542
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4632 10130 4752 10146
rect 4632 10124 4764 10130
rect 4632 10118 4712 10124
rect 4712 10066 4764 10072
rect 4526 9752 4582 9761
rect 4526 9687 4582 9696
rect 4724 9625 4752 10066
rect 4710 9616 4766 9625
rect 4710 9551 4766 9560
rect 4724 9178 4752 9551
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4816 9110 4844 10474
rect 4908 9178 4936 17836
rect 5078 17776 5134 17785
rect 4988 17740 5040 17746
rect 5078 17711 5134 17720
rect 4988 17682 5040 17688
rect 5000 17202 5028 17682
rect 5092 17678 5120 17711
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5092 17338 5120 17614
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 4988 17196 5040 17202
rect 5276 17184 5304 18142
rect 4988 17138 5040 17144
rect 5092 17156 5304 17184
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 5000 16833 5028 16934
rect 4986 16824 5042 16833
rect 4986 16759 5042 16768
rect 4988 14000 5040 14006
rect 4986 13968 4988 13977
rect 5040 13968 5042 13977
rect 4986 13903 5042 13912
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 5000 10810 5028 13262
rect 5092 13258 5120 17156
rect 5368 17082 5396 22714
rect 5460 22234 5488 23122
rect 6000 22976 6052 22982
rect 6000 22918 6052 22924
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5632 22432 5684 22438
rect 5630 22400 5632 22409
rect 5684 22400 5686 22409
rect 5630 22335 5686 22344
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 5644 22166 5672 22335
rect 5632 22160 5684 22166
rect 5632 22102 5684 22108
rect 6012 22001 6040 22918
rect 6196 22817 6224 24126
rect 6368 24132 6420 24138
rect 6368 24074 6420 24080
rect 6366 23896 6422 23905
rect 6366 23831 6422 23840
rect 6380 23662 6408 23831
rect 6368 23656 6420 23662
rect 6368 23598 6420 23604
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6366 22944 6422 22953
rect 6182 22808 6238 22817
rect 6182 22743 6238 22752
rect 6288 22574 6316 22918
rect 6366 22879 6422 22888
rect 6276 22568 6328 22574
rect 6276 22510 6328 22516
rect 6276 22432 6328 22438
rect 6276 22374 6328 22380
rect 6184 22228 6236 22234
rect 6184 22170 6236 22176
rect 5998 21992 6054 22001
rect 5998 21927 6054 21936
rect 6092 21888 6144 21894
rect 5998 21856 6054 21865
rect 5622 21788 5918 21808
rect 6092 21830 6144 21836
rect 5998 21791 6054 21800
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5460 21146 5488 21286
rect 5448 21140 5500 21146
rect 5448 21082 5500 21088
rect 5448 20936 5500 20942
rect 5552 20924 5580 21490
rect 6012 21457 6040 21791
rect 5998 21448 6054 21457
rect 5998 21383 6054 21392
rect 6104 21078 6132 21830
rect 6196 21418 6224 22170
rect 6184 21412 6236 21418
rect 6184 21354 6236 21360
rect 6092 21072 6144 21078
rect 6092 21014 6144 21020
rect 6000 21004 6052 21010
rect 6000 20946 6052 20952
rect 5500 20896 5580 20924
rect 5448 20878 5500 20884
rect 5552 19922 5580 20896
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6012 20602 6040 20946
rect 6092 20936 6144 20942
rect 6196 20924 6224 21354
rect 6144 20896 6224 20924
rect 6092 20878 6144 20884
rect 6000 20596 6052 20602
rect 6000 20538 6052 20544
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 5816 20392 5868 20398
rect 5814 20360 5816 20369
rect 5868 20360 5870 20369
rect 5814 20295 5870 20304
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5448 19780 5500 19786
rect 5448 19722 5500 19728
rect 5460 18970 5488 19722
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5644 18902 5672 19110
rect 5632 18896 5684 18902
rect 5552 18856 5632 18884
rect 5552 18426 5580 18856
rect 5632 18838 5684 18844
rect 6012 18737 6040 20402
rect 6104 20398 6132 20878
rect 6092 20392 6144 20398
rect 6092 20334 6144 20340
rect 6090 20224 6146 20233
rect 6090 20159 6146 20168
rect 5998 18728 6054 18737
rect 5998 18663 6054 18672
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5448 18148 5500 18154
rect 5448 18090 5500 18096
rect 5460 17882 5488 18090
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5644 17785 5672 18022
rect 5630 17776 5686 17785
rect 5460 17734 5630 17762
rect 5460 17338 5488 17734
rect 5630 17711 5686 17720
rect 5540 17604 5592 17610
rect 5540 17546 5592 17552
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5552 17202 5580 17546
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5276 17054 5396 17082
rect 5170 16008 5226 16017
rect 5170 15943 5226 15952
rect 5184 15910 5212 15943
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5184 14006 5212 14758
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 5092 10198 5120 13194
rect 5184 13161 5212 13466
rect 5170 13152 5226 13161
rect 5170 13087 5226 13096
rect 5184 12617 5212 13087
rect 5170 12608 5226 12617
rect 5170 12543 5226 12552
rect 5172 10736 5224 10742
rect 5170 10704 5172 10713
rect 5224 10704 5226 10713
rect 5170 10639 5226 10648
rect 5080 10192 5132 10198
rect 5080 10134 5132 10140
rect 5092 9722 5120 10134
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4710 8664 4766 8673
rect 4710 8599 4766 8608
rect 4724 8430 4752 8599
rect 4816 8498 4844 9046
rect 4908 8634 4936 9114
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5078 8528 5134 8537
rect 4804 8492 4856 8498
rect 5078 8463 5134 8472
rect 4804 8434 4856 8440
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4724 8090 4752 8366
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 5000 8090 5028 8230
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 4620 7744 4672 7750
rect 4434 7712 4490 7721
rect 4620 7686 4672 7692
rect 4434 7647 4490 7656
rect 4448 7002 4476 7647
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 4632 6798 4660 7686
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4724 6866 4752 7142
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4632 5914 4660 6734
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4986 6624 5042 6633
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4632 4758 4660 4966
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4620 4752 4672 4758
rect 4620 4694 4672 4700
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4526 3768 4582 3777
rect 4526 3703 4528 3712
rect 4580 3703 4582 3712
rect 4528 3674 4580 3680
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4448 3194 4476 3538
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4540 3126 4568 3674
rect 4632 3670 4660 3878
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 4436 2508 4488 2514
rect 4632 2496 4660 3606
rect 4816 3398 4844 4762
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4488 2468 4660 2496
rect 4436 2450 4488 2456
rect 4342 1456 4398 1465
rect 4342 1391 4398 1400
rect 2884 1006 3004 1034
rect 3436 1006 3556 1034
rect 2884 480 2912 1006
rect 3436 480 3464 1006
rect 4066 912 4122 921
rect 4066 847 4122 856
rect 3896 598 4016 626
rect 202 0 258 480
rect 662 0 718 480
rect 1214 0 1270 480
rect 1766 0 1822 480
rect 2318 0 2374 480
rect 2870 0 2926 480
rect 3422 0 3478 480
rect 3896 377 3924 598
rect 3988 480 4016 598
rect 3882 368 3938 377
rect 3882 303 3938 312
rect 3974 0 4030 480
rect 4080 241 4108 847
rect 4540 480 4568 2468
rect 4908 1465 4936 6598
rect 4986 6559 5042 6568
rect 5000 4146 5028 6559
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5092 3942 5120 8463
rect 5184 7449 5212 8774
rect 5276 8566 5304 17054
rect 5460 16833 5488 17138
rect 5446 16824 5502 16833
rect 5552 16794 5580 17138
rect 5446 16759 5502 16768
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5448 16448 5500 16454
rect 5354 16416 5410 16425
rect 5448 16390 5500 16396
rect 5354 16351 5410 16360
rect 5368 15484 5396 16351
rect 5460 15745 5488 16390
rect 5552 16250 5580 16730
rect 6104 16726 6132 20159
rect 6182 19680 6238 19689
rect 6182 19615 6238 19624
rect 6092 16720 6144 16726
rect 6092 16662 6144 16668
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5446 15736 5502 15745
rect 5644 15706 5672 15846
rect 5446 15671 5502 15680
rect 5632 15700 5684 15706
rect 5460 15638 5488 15671
rect 5632 15642 5684 15648
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5368 15456 5580 15484
rect 5552 15450 5580 15456
rect 5552 15422 6040 15450
rect 6104 15434 6132 16050
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5368 14482 5396 14758
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 5460 13938 5488 14758
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5354 13832 5410 13841
rect 5354 13767 5410 13776
rect 5368 13326 5396 13767
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5356 13320 5408 13326
rect 5460 13297 5488 13330
rect 5356 13262 5408 13268
rect 5446 13288 5502 13297
rect 5368 12986 5396 13262
rect 5446 13223 5502 13232
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5460 12918 5488 13223
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5368 12238 5396 12718
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5460 12442 5488 12582
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5552 12374 5580 14214
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6012 13705 6040 15422
rect 6092 15428 6144 15434
rect 6092 15370 6144 15376
rect 6196 14770 6224 19615
rect 6288 15609 6316 22374
rect 6380 22098 6408 22879
rect 6368 22092 6420 22098
rect 6368 22034 6420 22040
rect 6472 21962 6500 25094
rect 6564 24614 6592 25298
rect 6552 24608 6604 24614
rect 6552 24550 6604 24556
rect 6656 24313 6684 27520
rect 6828 25900 6880 25906
rect 6828 25842 6880 25848
rect 6736 24948 6788 24954
rect 6736 24890 6788 24896
rect 6642 24304 6698 24313
rect 6642 24239 6698 24248
rect 6644 24200 6696 24206
rect 6644 24142 6696 24148
rect 6552 24132 6604 24138
rect 6552 24074 6604 24080
rect 6564 22438 6592 24074
rect 6656 23594 6684 24142
rect 6644 23588 6696 23594
rect 6644 23530 6696 23536
rect 6552 22432 6604 22438
rect 6552 22374 6604 22380
rect 6748 22148 6776 24890
rect 6840 23882 6868 25842
rect 7104 24336 7156 24342
rect 7104 24278 7156 24284
rect 6840 23854 6960 23882
rect 6826 23760 6882 23769
rect 6826 23695 6882 23704
rect 6840 22778 6868 23695
rect 6932 23066 6960 23854
rect 7012 23520 7064 23526
rect 7010 23488 7012 23497
rect 7064 23488 7066 23497
rect 7010 23423 7066 23432
rect 6932 23038 7052 23066
rect 6920 22976 6972 22982
rect 6920 22918 6972 22924
rect 6828 22772 6880 22778
rect 6828 22714 6880 22720
rect 6932 22574 6960 22918
rect 6920 22568 6972 22574
rect 6920 22510 6972 22516
rect 7024 22506 7052 23038
rect 7012 22500 7064 22506
rect 7012 22442 7064 22448
rect 7116 22148 7144 24278
rect 7196 24268 7248 24274
rect 7196 24210 7248 24216
rect 7208 23322 7236 24210
rect 7300 23769 7328 27520
rect 7380 26172 7432 26178
rect 7380 26114 7432 26120
rect 7286 23760 7342 23769
rect 7286 23695 7342 23704
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 7392 22624 7420 26114
rect 7852 25158 7880 27520
rect 7932 25220 7984 25226
rect 7932 25162 7984 25168
rect 7656 25152 7708 25158
rect 7840 25152 7892 25158
rect 7656 25094 7708 25100
rect 7746 25120 7802 25129
rect 7472 24744 7524 24750
rect 7472 24686 7524 24692
rect 7484 23866 7512 24686
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7472 23860 7524 23866
rect 7472 23802 7524 23808
rect 7484 23662 7512 23802
rect 7472 23656 7524 23662
rect 7472 23598 7524 23604
rect 7470 23352 7526 23361
rect 7470 23287 7526 23296
rect 7300 22596 7420 22624
rect 7196 22568 7248 22574
rect 7196 22510 7248 22516
rect 6564 22120 6776 22148
rect 7024 22120 7144 22148
rect 6460 21956 6512 21962
rect 6460 21898 6512 21904
rect 6368 21888 6420 21894
rect 6368 21830 6420 21836
rect 6274 15600 6330 15609
rect 6274 15535 6330 15544
rect 6380 14822 6408 21830
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 6472 20602 6500 20878
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6472 18834 6500 19110
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 6472 18426 6500 18770
rect 6460 18420 6512 18426
rect 6460 18362 6512 18368
rect 6458 17640 6514 17649
rect 6458 17575 6514 17584
rect 6472 17542 6500 17575
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6564 17218 6592 22120
rect 6644 22024 6696 22030
rect 6644 21966 6696 21972
rect 6736 22024 6788 22030
rect 6736 21966 6788 21972
rect 6472 17190 6592 17218
rect 6368 14816 6420 14822
rect 6104 14742 6224 14770
rect 6366 14784 6368 14793
rect 6420 14784 6422 14793
rect 5998 13696 6054 13705
rect 5998 13631 6054 13640
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6012 12850 6040 13126
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5736 12481 5764 12582
rect 5722 12472 5778 12481
rect 6012 12442 6040 12786
rect 6104 12782 6132 14742
rect 6366 14719 6422 14728
rect 6182 14648 6238 14657
rect 6182 14583 6184 14592
rect 6236 14583 6238 14592
rect 6366 14648 6422 14657
rect 6366 14583 6422 14592
rect 6184 14554 6236 14560
rect 6380 14550 6408 14583
rect 6368 14544 6420 14550
rect 6368 14486 6420 14492
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 6288 13462 6316 13670
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6196 13190 6224 13330
rect 6288 13326 6316 13398
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 5722 12407 5778 12416
rect 6000 12436 6052 12442
rect 5540 12368 5592 12374
rect 5446 12336 5502 12345
rect 5540 12310 5592 12316
rect 5736 12322 5764 12407
rect 6000 12378 6052 12384
rect 5736 12294 5948 12322
rect 5446 12271 5502 12280
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5368 11830 5396 12174
rect 5460 12170 5488 12271
rect 5538 12200 5594 12209
rect 5448 12164 5500 12170
rect 5538 12135 5594 12144
rect 5920 12152 5948 12294
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 5448 12106 5500 12112
rect 5552 11898 5580 12135
rect 5920 12124 6040 12152
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5368 10742 5396 11290
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5460 10826 5488 11154
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5460 10810 5580 10826
rect 5460 10804 5592 10810
rect 5460 10798 5540 10804
rect 5540 10746 5592 10752
rect 5356 10736 5408 10742
rect 5356 10678 5408 10684
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5540 10192 5592 10198
rect 5538 10160 5540 10169
rect 5592 10160 5594 10169
rect 5538 10095 5594 10104
rect 5736 9994 5764 10406
rect 5828 10169 5856 10610
rect 5906 10432 5962 10441
rect 5906 10367 5962 10376
rect 5920 10266 5948 10367
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5814 10160 5870 10169
rect 5814 10095 5816 10104
rect 5868 10095 5870 10104
rect 5816 10066 5868 10072
rect 5828 10035 5856 10066
rect 5724 9988 5776 9994
rect 5724 9930 5776 9936
rect 5354 9888 5410 9897
rect 5410 9846 5580 9874
rect 5354 9823 5410 9832
rect 5552 9058 5580 9846
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 9217 5948 9318
rect 5906 9208 5962 9217
rect 5906 9143 5962 9152
rect 5816 9104 5868 9110
rect 5368 9030 5580 9058
rect 5814 9072 5816 9081
rect 5868 9072 5870 9081
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 5170 7440 5226 7449
rect 5170 7375 5172 7384
rect 5224 7375 5226 7384
rect 5172 7346 5224 7352
rect 5276 7274 5304 8502
rect 5368 7698 5396 9030
rect 5814 9007 5870 9016
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5460 8498 5488 8910
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5552 8265 5580 8774
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5630 8528 5686 8537
rect 5630 8463 5686 8472
rect 5644 8362 5672 8463
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5538 8256 5594 8265
rect 5538 8191 5594 8200
rect 5540 7744 5592 7750
rect 5368 7670 5488 7698
rect 5540 7686 5592 7692
rect 5354 7576 5410 7585
rect 5354 7511 5410 7520
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 5368 7177 5396 7511
rect 5354 7168 5410 7177
rect 5354 7103 5410 7112
rect 5262 6896 5318 6905
rect 5262 6831 5318 6840
rect 5276 6798 5304 6831
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5276 6304 5304 6734
rect 5184 6276 5304 6304
rect 5184 5817 5212 6276
rect 5460 6202 5488 7670
rect 5552 7342 5580 7686
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5276 6174 5488 6202
rect 5170 5808 5226 5817
rect 5170 5743 5226 5752
rect 5276 4010 5304 6174
rect 5448 6112 5500 6118
rect 5354 6080 5410 6089
rect 5448 6054 5500 6060
rect 5354 6015 5410 6024
rect 5368 5914 5396 6015
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5460 5710 5488 6054
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5368 5030 5396 5578
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5368 4282 5396 4966
rect 5460 4706 5488 5646
rect 5552 5642 5580 7278
rect 6012 6798 6040 12124
rect 6104 12073 6132 12242
rect 6196 12238 6224 13126
rect 6288 12646 6316 13262
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 6366 12608 6422 12617
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6090 12064 6146 12073
rect 6090 11999 6146 12008
rect 6090 11928 6146 11937
rect 6090 11863 6146 11872
rect 6104 11830 6132 11863
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 6196 11558 6224 12174
rect 6288 11830 6316 12582
rect 6366 12543 6422 12552
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6196 11234 6224 11494
rect 6288 11354 6316 11630
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6196 11206 6316 11234
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 6104 8022 6132 11018
rect 6196 9568 6224 11086
rect 6288 9994 6316 11206
rect 6380 10470 6408 12543
rect 6472 12209 6500 17190
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6564 16046 6592 16526
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6564 15910 6592 15982
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6564 15570 6592 15846
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6564 15094 6592 15506
rect 6552 15088 6604 15094
rect 6552 15030 6604 15036
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6564 13938 6592 14214
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6564 12889 6592 13874
rect 6550 12880 6606 12889
rect 6550 12815 6606 12824
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6458 12200 6514 12209
rect 6458 12135 6514 12144
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6472 11286 6500 12038
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6458 10296 6514 10305
rect 6458 10231 6460 10240
rect 6512 10231 6514 10240
rect 6460 10202 6512 10208
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 6288 9722 6316 9930
rect 6380 9897 6408 9998
rect 6366 9888 6422 9897
rect 6366 9823 6422 9832
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6196 9540 6316 9568
rect 6182 9480 6238 9489
rect 6182 9415 6238 9424
rect 6196 9217 6224 9415
rect 6182 9208 6238 9217
rect 6182 9143 6238 9152
rect 6182 8936 6238 8945
rect 6182 8871 6238 8880
rect 6196 8430 6224 8871
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 6104 7546 6132 7958
rect 6196 7954 6224 8230
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6104 6882 6132 7482
rect 6196 7342 6224 7890
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6288 7002 6316 9540
rect 6380 9382 6408 9823
rect 6472 9722 6500 10202
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6380 7750 6408 8978
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6276 6996 6328 7002
rect 6196 6934 6224 6965
rect 6276 6938 6328 6944
rect 6184 6928 6236 6934
rect 6104 6876 6184 6882
rect 6104 6870 6236 6876
rect 6104 6854 6224 6870
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6090 6760 6146 6769
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6012 6458 6040 6734
rect 6090 6695 6092 6704
rect 6144 6695 6146 6704
rect 6092 6666 6144 6672
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 6104 5914 6132 6666
rect 6196 6390 6224 6854
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6184 6384 6236 6390
rect 6184 6326 6236 6332
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6182 5808 6238 5817
rect 6092 5772 6144 5778
rect 6182 5743 6238 5752
rect 6092 5714 6144 5720
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5722 5264 5778 5273
rect 5722 5199 5724 5208
rect 5776 5199 5778 5208
rect 5724 5170 5776 5176
rect 6000 4752 6052 4758
rect 5460 4678 5580 4706
rect 6000 4694 6052 4700
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5448 4208 5500 4214
rect 5448 4150 5500 4156
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5276 3738 5304 3946
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5170 3632 5226 3641
rect 5170 3567 5226 3576
rect 5184 3534 5212 3567
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5184 3194 5212 3470
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 4894 1456 4950 1465
rect 4894 1391 4950 1400
rect 4066 232 4122 241
rect 4066 167 4122 176
rect 4526 0 4582 480
rect 5000 377 5028 3130
rect 5460 2938 5488 4150
rect 5552 3058 5580 4678
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5908 3596 5960 3602
rect 6012 3584 6040 4694
rect 6104 4214 6132 5714
rect 6092 4208 6144 4214
rect 6092 4150 6144 4156
rect 6196 4078 6224 5743
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 5960 3556 6040 3584
rect 5908 3538 5960 3544
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 6000 2984 6052 2990
rect 5460 2910 5580 2938
rect 6000 2926 6052 2932
rect 5552 2650 5580 2910
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 5092 480 5120 2450
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6012 2145 6040 2926
rect 5998 2136 6054 2145
rect 5998 2071 6054 2080
rect 5632 1692 5684 1698
rect 5632 1634 5684 1640
rect 5644 480 5672 1634
rect 6104 1329 6132 4014
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6196 3670 6224 3878
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6090 1320 6146 1329
rect 6090 1255 6146 1264
rect 6196 480 6224 3130
rect 6288 513 6316 6802
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6380 4185 6408 5510
rect 6366 4176 6422 4185
rect 6366 4111 6422 4120
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6380 2922 6408 4014
rect 6472 3641 6500 8774
rect 6564 6662 6592 12718
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6564 5846 6592 6598
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6564 5030 6592 5646
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6564 4622 6592 4966
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6564 3942 6592 4558
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6458 3632 6514 3641
rect 6458 3567 6514 3576
rect 6368 2916 6420 2922
rect 6368 2858 6420 2864
rect 6564 2650 6592 3878
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6656 1698 6684 21966
rect 6748 21350 6776 21966
rect 6828 21616 6880 21622
rect 6828 21558 6880 21564
rect 6736 21344 6788 21350
rect 6736 21286 6788 21292
rect 6748 21185 6776 21286
rect 6734 21176 6790 21185
rect 6734 21111 6790 21120
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6748 20097 6776 20742
rect 6840 20602 6868 21558
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6932 20233 6960 20742
rect 6918 20224 6974 20233
rect 6918 20159 6974 20168
rect 6734 20088 6790 20097
rect 6734 20023 6790 20032
rect 6736 19916 6788 19922
rect 6736 19858 6788 19864
rect 6748 19174 6776 19858
rect 6736 19168 6788 19174
rect 6736 19110 6788 19116
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6748 18630 6776 19110
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6748 16726 6776 18158
rect 6932 18057 6960 19110
rect 6918 18048 6974 18057
rect 6918 17983 6974 17992
rect 6828 17808 6880 17814
rect 6828 17750 6880 17756
rect 6840 17338 6868 17750
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6736 16720 6788 16726
rect 6736 16662 6788 16668
rect 6748 16250 6776 16662
rect 6840 16538 6868 17274
rect 6932 16969 6960 17614
rect 7024 17218 7052 22120
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7116 21486 7144 21966
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 7116 21146 7144 21422
rect 7104 21140 7156 21146
rect 7104 21082 7156 21088
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7116 18698 7144 20402
rect 7208 20369 7236 22510
rect 7300 21894 7328 22596
rect 7380 22500 7432 22506
rect 7380 22442 7432 22448
rect 7288 21888 7340 21894
rect 7288 21830 7340 21836
rect 7288 20868 7340 20874
rect 7288 20810 7340 20816
rect 7194 20360 7250 20369
rect 7194 20295 7250 20304
rect 7196 20256 7248 20262
rect 7300 20244 7328 20810
rect 7248 20216 7328 20244
rect 7196 20198 7248 20204
rect 7208 20058 7236 20198
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7392 18873 7420 22442
rect 7484 19718 7512 23287
rect 7576 22642 7604 24006
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 7564 21888 7616 21894
rect 7564 21830 7616 21836
rect 7576 21486 7604 21830
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7576 20330 7604 21422
rect 7564 20324 7616 20330
rect 7564 20266 7616 20272
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7576 19514 7604 20266
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 7378 18864 7434 18873
rect 7378 18799 7434 18808
rect 7104 18692 7156 18698
rect 7104 18634 7156 18640
rect 7116 18426 7144 18634
rect 7378 18592 7434 18601
rect 7378 18527 7434 18536
rect 7104 18420 7156 18426
rect 7104 18362 7156 18368
rect 7392 17320 7420 18527
rect 7484 18465 7512 19110
rect 7668 18902 7696 25094
rect 7840 25094 7892 25100
rect 7746 25055 7802 25064
rect 7656 18896 7708 18902
rect 7656 18838 7708 18844
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7470 18456 7526 18465
rect 7470 18391 7526 18400
rect 7472 18080 7524 18086
rect 7470 18048 7472 18057
rect 7576 18068 7604 18770
rect 7668 18222 7696 18838
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7524 18048 7604 18068
rect 7526 18040 7604 18048
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7470 17983 7526 17992
rect 7668 17882 7696 18022
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7392 17292 7512 17320
rect 7024 17190 7420 17218
rect 7012 16992 7064 16998
rect 6918 16960 6974 16969
rect 7012 16934 7064 16940
rect 7194 16960 7250 16969
rect 6918 16895 6974 16904
rect 7024 16697 7052 16934
rect 7194 16895 7250 16904
rect 7010 16688 7066 16697
rect 7010 16623 7066 16632
rect 6840 16510 7052 16538
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6748 15638 6776 16186
rect 7024 16130 7052 16510
rect 7024 16102 7144 16130
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 6734 15056 6790 15065
rect 6734 14991 6790 15000
rect 6748 14482 6776 14991
rect 6840 14600 6868 15846
rect 7010 15328 7066 15337
rect 7010 15263 7066 15272
rect 6920 14612 6972 14618
rect 6840 14572 6920 14600
rect 6920 14554 6972 14560
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6918 14376 6974 14385
rect 6918 14311 6920 14320
rect 6972 14311 6974 14320
rect 6920 14282 6972 14288
rect 6734 13424 6790 13433
rect 6734 13359 6790 13368
rect 6748 13161 6776 13359
rect 6734 13152 6790 13161
rect 6734 13087 6790 13096
rect 6748 12617 6776 13087
rect 7024 12918 7052 15263
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 6828 12640 6880 12646
rect 6734 12608 6790 12617
rect 6828 12582 6880 12588
rect 6734 12543 6790 12552
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6748 11898 6776 12378
rect 6840 12306 6868 12582
rect 7024 12442 7052 12854
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6734 11656 6790 11665
rect 6734 11591 6790 11600
rect 6748 9586 6776 11591
rect 6840 11529 6868 12242
rect 6826 11520 6882 11529
rect 6826 11455 6882 11464
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6840 10810 6868 11290
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6644 1692 6696 1698
rect 6644 1634 6696 1640
rect 6274 504 6330 513
rect 4986 368 5042 377
rect 4986 303 5042 312
rect 5078 0 5134 480
rect 5630 0 5686 480
rect 6182 0 6238 480
rect 6748 480 6776 9386
rect 6840 6984 6868 10746
rect 6932 7993 6960 12310
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7024 12102 7052 12242
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7024 11626 7052 11834
rect 7012 11620 7064 11626
rect 7012 11562 7064 11568
rect 7024 11354 7052 11562
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 7012 10736 7064 10742
rect 7012 10678 7064 10684
rect 7024 9586 7052 10678
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7012 9104 7064 9110
rect 7012 9046 7064 9052
rect 7024 8498 7052 9046
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 6918 7984 6974 7993
rect 6918 7919 6974 7928
rect 7024 7750 7052 8230
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7116 7562 7144 16102
rect 7208 15162 7236 16895
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7208 13394 7236 14894
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7300 12782 7328 13126
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 12306 7328 12582
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7024 7534 7144 7562
rect 6840 6956 6960 6984
rect 6826 6896 6882 6905
rect 6826 6831 6882 6840
rect 6840 6322 6868 6831
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6932 6202 6960 6956
rect 6840 6174 6960 6202
rect 6840 5778 6868 6174
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6828 5364 6880 5370
rect 6932 5352 6960 5782
rect 7024 5370 7052 7534
rect 7104 7472 7156 7478
rect 7102 7440 7104 7449
rect 7156 7440 7158 7449
rect 7102 7375 7158 7384
rect 7208 7313 7236 11494
rect 7300 10849 7328 12106
rect 7392 11218 7420 17190
rect 7484 15638 7512 17292
rect 7654 17232 7710 17241
rect 7760 17218 7788 25055
rect 7852 21049 7880 25094
rect 7944 24886 7972 25162
rect 7932 24880 7984 24886
rect 7932 24822 7984 24828
rect 8404 24834 8432 27520
rect 8760 25152 8812 25158
rect 8760 25094 8812 25100
rect 7944 24614 7972 24822
rect 8404 24806 8616 24834
rect 7932 24608 7984 24614
rect 7932 24550 7984 24556
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 8208 24608 8260 24614
rect 8208 24550 8260 24556
rect 7944 22506 7972 24550
rect 8022 23080 8078 23089
rect 8022 23015 8024 23024
rect 8076 23015 8078 23024
rect 8024 22986 8076 22992
rect 7932 22500 7984 22506
rect 7932 22442 7984 22448
rect 7838 21040 7894 21049
rect 7838 20975 7894 20984
rect 7932 21004 7984 21010
rect 7932 20946 7984 20952
rect 7840 20392 7892 20398
rect 7840 20334 7892 20340
rect 7852 20058 7880 20334
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 7944 19825 7972 20946
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 7930 19816 7986 19825
rect 7930 19751 7932 19760
rect 7984 19751 7986 19760
rect 7932 19722 7984 19728
rect 7932 19236 7984 19242
rect 7932 19178 7984 19184
rect 7944 18630 7972 19178
rect 8036 18970 8064 19858
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7932 18624 7984 18630
rect 7932 18566 7984 18572
rect 7852 18358 7880 18566
rect 7840 18352 7892 18358
rect 7840 18294 7892 18300
rect 7840 18148 7892 18154
rect 7840 18090 7892 18096
rect 7852 18057 7880 18090
rect 7838 18048 7894 18057
rect 7838 17983 7894 17992
rect 7944 17626 7972 18566
rect 8128 18290 8156 24550
rect 8220 24138 8248 24550
rect 8208 24132 8260 24138
rect 8208 24074 8260 24080
rect 8220 22234 8248 24074
rect 8484 23112 8536 23118
rect 8484 23054 8536 23060
rect 8496 22953 8524 23054
rect 8482 22944 8538 22953
rect 8482 22879 8538 22888
rect 8208 22228 8260 22234
rect 8208 22170 8260 22176
rect 8392 22160 8444 22166
rect 8392 22102 8444 22108
rect 8300 21956 8352 21962
rect 8300 21898 8352 21904
rect 8312 21418 8340 21898
rect 8300 21412 8352 21418
rect 8300 21354 8352 21360
rect 8312 21146 8340 21354
rect 8404 21350 8432 22102
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8404 21185 8432 21286
rect 8390 21176 8446 21185
rect 8300 21140 8352 21146
rect 8390 21111 8446 21120
rect 8300 21082 8352 21088
rect 8208 21072 8260 21078
rect 8260 21020 8432 21026
rect 8208 21014 8432 21020
rect 8220 20998 8432 21014
rect 8206 20768 8262 20777
rect 8206 20703 8262 20712
rect 8220 18290 8248 20703
rect 8298 20088 8354 20097
rect 8298 20023 8300 20032
rect 8352 20023 8354 20032
rect 8300 19994 8352 20000
rect 8312 19514 8340 19994
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8404 18426 8432 20998
rect 8496 20874 8524 21966
rect 8484 20868 8536 20874
rect 8484 20810 8536 20816
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 8220 17882 8248 18226
rect 8208 17876 8260 17882
rect 8588 17864 8616 24806
rect 8772 24614 8800 25094
rect 8760 24608 8812 24614
rect 8760 24550 8812 24556
rect 8850 24576 8906 24585
rect 8668 24064 8720 24070
rect 8666 24032 8668 24041
rect 8720 24032 8722 24041
rect 8666 23967 8722 23976
rect 8680 23662 8708 23967
rect 8668 23656 8720 23662
rect 8668 23598 8720 23604
rect 8772 21593 8800 24550
rect 8850 24511 8906 24520
rect 8758 21584 8814 21593
rect 8758 21519 8814 21528
rect 8760 20256 8812 20262
rect 8760 20198 8812 20204
rect 8772 19854 8800 20198
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 8680 18329 8708 18634
rect 8772 18358 8800 19790
rect 8864 18834 8892 24511
rect 9048 24177 9076 27520
rect 9496 25492 9548 25498
rect 9496 25434 9548 25440
rect 9218 25392 9274 25401
rect 9218 25327 9274 25336
rect 9126 24440 9182 24449
rect 9126 24375 9182 24384
rect 9034 24168 9090 24177
rect 9034 24103 9090 24112
rect 9036 23044 9088 23050
rect 9036 22986 9088 22992
rect 8944 22500 8996 22506
rect 8944 22442 8996 22448
rect 8956 21690 8984 22442
rect 8944 21684 8996 21690
rect 8944 21626 8996 21632
rect 9048 21146 9076 22986
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8760 18352 8812 18358
rect 8666 18320 8722 18329
rect 8760 18294 8812 18300
rect 8666 18255 8722 18264
rect 8864 18086 8892 18770
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8942 18456 8998 18465
rect 8942 18391 8998 18400
rect 8956 18222 8984 18391
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 8208 17818 8260 17824
rect 8404 17836 8616 17864
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 7944 17598 8156 17626
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 7760 17190 7972 17218
rect 7654 17167 7710 17176
rect 7562 15736 7618 15745
rect 7562 15671 7618 15680
rect 7472 15632 7524 15638
rect 7472 15574 7524 15580
rect 7484 14822 7512 15574
rect 7576 15026 7604 15671
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7286 10840 7342 10849
rect 7286 10775 7288 10784
rect 7340 10775 7342 10784
rect 7288 10746 7340 10752
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7300 9926 7328 10406
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7194 7304 7250 7313
rect 7194 7239 7250 7248
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 7116 6458 7144 6938
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7194 6352 7250 6361
rect 7194 6287 7250 6296
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 6880 5324 6960 5352
rect 6828 5306 6880 5312
rect 6932 3942 6960 5324
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6828 3120 6880 3126
rect 6826 3088 6828 3097
rect 6880 3088 6882 3097
rect 6826 3023 6882 3032
rect 7116 2922 7144 5850
rect 7208 5846 7236 6287
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7194 5536 7250 5545
rect 7194 5471 7250 5480
rect 7208 3194 7236 5471
rect 7300 4298 7328 9862
rect 7392 9382 7420 9998
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 8106 7420 9318
rect 7484 8242 7512 14758
rect 7576 14550 7604 14962
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7576 10010 7604 12310
rect 7668 10713 7696 17167
rect 7746 15464 7802 15473
rect 7746 15399 7748 15408
rect 7800 15399 7802 15408
rect 7748 15370 7800 15376
rect 7746 15192 7802 15201
rect 7746 15127 7802 15136
rect 7760 14958 7788 15127
rect 7748 14952 7800 14958
rect 7800 14900 7880 14906
rect 7748 14894 7880 14900
rect 7760 14878 7880 14894
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 7760 13530 7788 13806
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7760 11558 7788 12242
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7746 11248 7802 11257
rect 7746 11183 7802 11192
rect 7654 10704 7710 10713
rect 7654 10639 7710 10648
rect 7654 10024 7710 10033
rect 7576 9982 7654 10010
rect 7654 9959 7656 9968
rect 7708 9959 7710 9968
rect 7656 9930 7708 9936
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7576 9761 7604 9862
rect 7562 9752 7618 9761
rect 7562 9687 7618 9696
rect 7760 9450 7788 11183
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7668 9081 7696 9318
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7654 9072 7710 9081
rect 7654 9007 7710 9016
rect 7484 8214 7604 8242
rect 7392 8078 7512 8106
rect 7378 7304 7434 7313
rect 7378 7239 7380 7248
rect 7432 7239 7434 7248
rect 7380 7210 7432 7216
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7392 6186 7420 6598
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7484 5545 7512 8078
rect 7576 7698 7604 8214
rect 7576 7670 7696 7698
rect 7562 7576 7618 7585
rect 7562 7511 7618 7520
rect 7576 7342 7604 7511
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7470 5536 7526 5545
rect 7470 5471 7526 5480
rect 7576 4729 7604 7142
rect 7562 4720 7618 4729
rect 7562 4655 7618 4664
rect 7300 4270 7420 4298
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7300 3058 7328 3334
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7196 2984 7248 2990
rect 7392 2938 7420 4270
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7484 3058 7512 3946
rect 7562 3904 7618 3913
rect 7562 3839 7618 3848
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7196 2926 7248 2932
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 7208 921 7236 2926
rect 7300 2910 7420 2938
rect 7194 912 7250 921
rect 7194 847 7250 856
rect 7300 480 7328 2910
rect 7470 640 7526 649
rect 7576 626 7604 3839
rect 7668 2836 7696 7670
rect 7760 7206 7788 9114
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 7760 6254 7788 6802
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7760 5030 7788 6190
rect 7852 5370 7880 14878
rect 7944 12306 7972 17190
rect 8036 17105 8064 17478
rect 8022 17096 8078 17105
rect 8022 17031 8078 17040
rect 8128 16454 8156 17598
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8022 16144 8078 16153
rect 8022 16079 8078 16088
rect 8036 15473 8064 16079
rect 8116 15632 8168 15638
rect 8116 15574 8168 15580
rect 8022 15464 8078 15473
rect 8022 15399 8078 15408
rect 8128 15162 8156 15574
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8024 14612 8076 14618
rect 8220 14600 8248 17070
rect 8312 16998 8340 17682
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8312 16794 8340 16934
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8404 16266 8432 17836
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8496 16289 8524 17614
rect 8588 17377 8616 17614
rect 8760 17604 8812 17610
rect 8760 17546 8812 17552
rect 8574 17368 8630 17377
rect 8574 17303 8576 17312
rect 8628 17303 8630 17312
rect 8576 17274 8628 17280
rect 8588 17243 8616 17274
rect 8772 17202 8800 17546
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8312 16238 8432 16266
rect 8482 16280 8538 16289
rect 8312 15570 8340 16238
rect 8482 16215 8538 16224
rect 8390 16144 8446 16153
rect 8390 16079 8446 16088
rect 8404 15638 8432 16079
rect 8574 15736 8630 15745
rect 8758 15736 8814 15745
rect 8574 15671 8630 15680
rect 8680 15694 8758 15722
rect 8392 15632 8444 15638
rect 8392 15574 8444 15580
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8312 15162 8340 15506
rect 8588 15502 8616 15671
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8484 15428 8536 15434
rect 8484 15370 8536 15376
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8392 14884 8444 14890
rect 8392 14826 8444 14832
rect 8300 14612 8352 14618
rect 8220 14572 8300 14600
rect 8024 14554 8076 14560
rect 8300 14554 8352 14560
rect 8036 14385 8064 14554
rect 8022 14376 8078 14385
rect 8022 14311 8078 14320
rect 8206 14104 8262 14113
rect 8206 14039 8262 14048
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 8128 12186 8156 13466
rect 8220 12442 8248 14039
rect 8312 13530 8340 14554
rect 8404 14006 8432 14826
rect 8496 14074 8524 15370
rect 8680 15337 8708 15694
rect 8758 15671 8814 15680
rect 8864 15337 8892 18022
rect 8944 17808 8996 17814
rect 8944 17750 8996 17756
rect 8956 17649 8984 17750
rect 8942 17640 8998 17649
rect 8942 17575 8998 17584
rect 9048 17134 9076 18566
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 9140 16250 9168 24375
rect 9232 21622 9260 25327
rect 9402 24984 9458 24993
rect 9402 24919 9458 24928
rect 9416 24342 9444 24919
rect 9508 24857 9536 25434
rect 9494 24848 9550 24857
rect 9494 24783 9550 24792
rect 9496 24744 9548 24750
rect 9496 24686 9548 24692
rect 9508 24614 9536 24686
rect 9496 24608 9548 24614
rect 9496 24550 9548 24556
rect 9508 24449 9536 24550
rect 9494 24440 9550 24449
rect 9494 24375 9550 24384
rect 9404 24336 9456 24342
rect 9404 24278 9456 24284
rect 9496 23520 9548 23526
rect 9496 23462 9548 23468
rect 9508 23254 9536 23462
rect 9496 23248 9548 23254
rect 9496 23190 9548 23196
rect 9600 23066 9628 27520
rect 10046 26480 10102 26489
rect 10046 26415 10102 26424
rect 9956 25696 10008 25702
rect 9956 25638 10008 25644
rect 9968 25498 9996 25638
rect 9956 25492 10008 25498
rect 9956 25434 10008 25440
rect 9772 25356 9824 25362
rect 9772 25298 9824 25304
rect 9784 25158 9812 25298
rect 9772 25152 9824 25158
rect 9772 25094 9824 25100
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9692 23322 9720 24550
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 9680 23180 9732 23186
rect 9680 23122 9732 23128
rect 9324 23038 9628 23066
rect 9220 21616 9272 21622
rect 9220 21558 9272 21564
rect 9218 21176 9274 21185
rect 9218 21111 9274 21120
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9036 15360 9088 15366
rect 8666 15328 8722 15337
rect 8666 15263 8722 15272
rect 8850 15328 8906 15337
rect 9036 15302 9088 15308
rect 8850 15263 8906 15272
rect 9048 14890 9076 15302
rect 9036 14884 9088 14890
rect 9036 14826 9088 14832
rect 8574 14648 8630 14657
rect 8574 14583 8630 14592
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 8404 13841 8432 13942
rect 8390 13832 8446 13841
rect 8390 13767 8446 13776
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8496 13410 8524 14010
rect 8312 13382 8524 13410
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8312 12345 8340 13382
rect 8392 12912 8444 12918
rect 8390 12880 8392 12889
rect 8444 12880 8446 12889
rect 8390 12815 8446 12824
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8298 12336 8354 12345
rect 8298 12271 8354 12280
rect 7944 12158 8156 12186
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 7944 10826 7972 12158
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11801 8064 12038
rect 8220 11898 8248 12174
rect 8298 12064 8354 12073
rect 8298 11999 8354 12008
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8022 11792 8078 11801
rect 8206 11792 8262 11801
rect 8022 11727 8078 11736
rect 8128 11750 8206 11778
rect 8128 11082 8156 11750
rect 8206 11727 8262 11736
rect 8206 11656 8262 11665
rect 8206 11591 8262 11600
rect 8220 11354 8248 11591
rect 8312 11354 8340 11999
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8298 11248 8354 11257
rect 8208 11212 8260 11218
rect 8298 11183 8354 11192
rect 8208 11154 8260 11160
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 7944 10798 8156 10826
rect 7930 10704 7986 10713
rect 7930 10639 7986 10648
rect 8024 10668 8076 10674
rect 7944 10606 7972 10639
rect 8024 10610 8076 10616
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7944 9586 7972 10066
rect 8036 9994 8064 10610
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 8022 9616 8078 9625
rect 7932 9580 7984 9586
rect 8022 9551 8078 9560
rect 7932 9522 7984 9528
rect 7944 9178 7972 9522
rect 8036 9518 8064 9551
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 7944 8362 7972 8774
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7944 7886 7972 8298
rect 7932 7880 7984 7886
rect 7930 7848 7932 7857
rect 7984 7848 7986 7857
rect 7930 7783 7986 7792
rect 7944 7410 7972 7783
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 7930 7032 7986 7041
rect 7930 6967 7986 6976
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7944 5302 7972 6967
rect 7932 5296 7984 5302
rect 8036 5273 8064 7686
rect 8128 7018 8156 10798
rect 8220 10470 8248 11154
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8220 9586 8248 9862
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8220 7546 8248 7822
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8312 7426 8340 11183
rect 8404 9654 8432 12718
rect 8496 12238 8524 12786
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8588 11898 8616 14583
rect 9128 14544 9180 14550
rect 9128 14486 9180 14492
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8680 13530 8708 14350
rect 9034 13968 9090 13977
rect 9034 13903 9090 13912
rect 8942 13560 8998 13569
rect 8668 13524 8720 13530
rect 9048 13530 9076 13903
rect 9140 13870 9168 14486
rect 9128 13864 9180 13870
rect 9126 13832 9128 13841
rect 9180 13832 9182 13841
rect 9126 13767 9182 13776
rect 9126 13696 9182 13705
rect 9126 13631 9182 13640
rect 8942 13495 8998 13504
rect 9036 13524 9088 13530
rect 8668 13466 8720 13472
rect 8956 13410 8984 13495
rect 9036 13466 9088 13472
rect 8956 13382 9076 13410
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8666 12336 8722 12345
rect 8666 12271 8722 12280
rect 8760 12300 8812 12306
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8404 7546 8432 7890
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8312 7398 8432 7426
rect 8128 6990 8248 7018
rect 8220 6866 8248 6990
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8128 6497 8156 6802
rect 8114 6488 8170 6497
rect 8114 6423 8116 6432
rect 8168 6423 8170 6432
rect 8116 6394 8168 6400
rect 8128 6363 8156 6394
rect 8220 6118 8248 6802
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8220 5896 8248 6054
rect 8312 5914 8340 6122
rect 8128 5868 8248 5896
rect 8300 5908 8352 5914
rect 7932 5238 7984 5244
rect 8022 5264 8078 5273
rect 8022 5199 8078 5208
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 8036 3641 8064 5102
rect 8022 3632 8078 3641
rect 8022 3567 8078 3576
rect 7838 3496 7894 3505
rect 7838 3431 7840 3440
rect 7892 3431 7894 3440
rect 7840 3402 7892 3408
rect 8128 2990 8156 5868
rect 8300 5850 8352 5856
rect 8312 5817 8340 5850
rect 8298 5808 8354 5817
rect 8298 5743 8354 5752
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8312 3777 8340 4694
rect 8298 3768 8354 3777
rect 8298 3703 8354 3712
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 7944 2854 7972 2885
rect 8220 2854 8248 2926
rect 7932 2848 7984 2854
rect 7668 2808 7788 2836
rect 7760 2666 7788 2808
rect 7930 2816 7932 2825
rect 8208 2848 8260 2854
rect 7984 2816 7986 2825
rect 8208 2790 8260 2796
rect 7930 2751 7986 2760
rect 7760 2638 7880 2666
rect 7526 598 7604 626
rect 7470 575 7526 584
rect 7852 480 7880 2638
rect 7944 2582 7972 2751
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 8220 2514 8248 2790
rect 8312 2650 8340 3703
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8404 480 8432 7398
rect 8496 3913 8524 10406
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8588 9110 8616 9998
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8680 8090 8708 12271
rect 8760 12242 8812 12248
rect 8772 10554 8800 12242
rect 8864 11801 8892 12582
rect 8850 11792 8906 11801
rect 8850 11727 8906 11736
rect 8772 10526 8892 10554
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 8588 7585 8616 7958
rect 8574 7576 8630 7585
rect 8574 7511 8630 7520
rect 8588 7478 8616 7511
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8680 6882 8708 8026
rect 8588 6854 8708 6882
rect 8588 5250 8616 6854
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8680 5370 8708 6734
rect 8772 6225 8800 10406
rect 8864 7041 8892 10526
rect 8956 9518 8984 12922
rect 9048 12442 9076 13382
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 9140 11898 9168 13631
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 9048 10674 9076 10950
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9232 10130 9260 21111
rect 9324 20913 9352 23038
rect 9496 22976 9548 22982
rect 9494 22944 9496 22953
rect 9548 22944 9550 22953
rect 9692 22930 9720 23122
rect 9494 22879 9550 22888
rect 9600 22902 9720 22930
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 9416 22098 9444 22714
rect 9404 22092 9456 22098
rect 9404 22034 9456 22040
rect 9600 22030 9628 22902
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9692 21622 9720 22034
rect 9680 21616 9732 21622
rect 9680 21558 9732 21564
rect 9680 21480 9732 21486
rect 9680 21422 9732 21428
rect 9692 21010 9720 21422
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9310 20904 9366 20913
rect 9310 20839 9366 20848
rect 9588 20868 9640 20874
rect 9588 20810 9640 20816
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9310 20632 9366 20641
rect 9310 20567 9366 20576
rect 9324 15434 9352 20567
rect 9416 18154 9444 20742
rect 9600 20602 9628 20810
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 9692 20398 9720 20946
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9678 20224 9734 20233
rect 9678 20159 9734 20168
rect 9692 20058 9720 20159
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9588 19780 9640 19786
rect 9588 19722 9640 19728
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9508 19514 9536 19654
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9494 19408 9550 19417
rect 9494 19343 9550 19352
rect 9404 18148 9456 18154
rect 9404 18090 9456 18096
rect 9508 18034 9536 19343
rect 9600 18290 9628 19722
rect 9678 18864 9734 18873
rect 9678 18799 9680 18808
rect 9732 18799 9734 18808
rect 9680 18770 9732 18776
rect 9692 18426 9720 18770
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9508 18006 9628 18034
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9416 17241 9444 17478
rect 9402 17232 9458 17241
rect 9402 17167 9458 17176
rect 9496 17196 9548 17202
rect 9496 17138 9548 17144
rect 9508 17066 9536 17138
rect 9496 17060 9548 17066
rect 9496 17002 9548 17008
rect 9508 16794 9536 17002
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9600 16130 9628 18006
rect 9678 17912 9734 17921
rect 9678 17847 9680 17856
rect 9732 17847 9734 17856
rect 9680 17818 9732 17824
rect 9692 17270 9720 17818
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9692 16250 9720 17070
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9600 16102 9720 16130
rect 9692 15434 9720 16102
rect 9312 15428 9364 15434
rect 9312 15370 9364 15376
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9402 15192 9458 15201
rect 9312 15156 9364 15162
rect 9402 15127 9458 15136
rect 9312 15098 9364 15104
rect 9324 13977 9352 15098
rect 9310 13968 9366 13977
rect 9310 13903 9366 13912
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9324 12442 9352 13330
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9416 12306 9444 15127
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9600 14278 9628 14894
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9600 13870 9628 14214
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9678 13832 9734 13841
rect 9496 13796 9548 13802
rect 9678 13767 9734 13776
rect 9496 13738 9548 13744
rect 9508 13530 9536 13738
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9508 12986 9536 13262
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9692 12594 9720 13767
rect 9600 12566 9720 12594
rect 9600 12306 9628 12566
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8956 9178 8984 9454
rect 9048 9382 9076 9454
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 9048 8974 9076 9318
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9048 8430 9076 8910
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 8850 7032 8906 7041
rect 8850 6967 8906 6976
rect 9048 6798 9076 8366
rect 9218 7304 9274 7313
rect 9218 7239 9274 7248
rect 9232 7206 9260 7239
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8758 6216 8814 6225
rect 8758 6151 8814 6160
rect 8850 5944 8906 5953
rect 8850 5879 8852 5888
rect 8904 5879 8906 5888
rect 8852 5850 8904 5856
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8588 5222 8708 5250
rect 8574 4448 8630 4457
rect 8574 4383 8630 4392
rect 8482 3904 8538 3913
rect 8482 3839 8538 3848
rect 8588 3602 8616 4383
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8680 3516 8708 5222
rect 8956 5001 8984 6666
rect 9232 5710 9260 6734
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 8942 4992 8998 5001
rect 8942 4927 8998 4936
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8864 3942 8892 4422
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8864 3670 8892 3878
rect 8852 3664 8904 3670
rect 8852 3606 8904 3612
rect 8680 3488 8892 3516
rect 8668 3392 8720 3398
rect 8574 3360 8630 3369
rect 8668 3334 8720 3340
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8574 3295 8630 3304
rect 8588 2961 8616 3295
rect 8680 2990 8708 3334
rect 8668 2984 8720 2990
rect 8574 2952 8630 2961
rect 8772 2961 8800 3334
rect 8668 2926 8720 2932
rect 8758 2952 8814 2961
rect 8574 2887 8630 2896
rect 8680 2553 8708 2926
rect 8758 2887 8814 2896
rect 8864 2666 8892 3488
rect 8956 3097 8984 4762
rect 9140 4146 9168 5578
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9232 4593 9260 5510
rect 9218 4584 9274 4593
rect 9218 4519 9274 4528
rect 9218 4312 9274 4321
rect 9218 4247 9274 4256
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 8942 3088 8998 3097
rect 8942 3023 8998 3032
rect 9232 2689 9260 4247
rect 9324 4078 9352 12174
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9416 9450 9444 12106
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9508 11354 9536 11698
rect 9692 11642 9720 12378
rect 9600 11614 9720 11642
rect 9600 11393 9628 11614
rect 9678 11520 9734 11529
rect 9678 11455 9734 11464
rect 9586 11384 9642 11393
rect 9496 11348 9548 11354
rect 9586 11319 9642 11328
rect 9496 11290 9548 11296
rect 9508 10266 9536 11290
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9508 9994 9536 10202
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9508 9722 9536 9930
rect 9600 9926 9628 10406
rect 9692 10266 9720 11455
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9494 9616 9550 9625
rect 9494 9551 9550 9560
rect 9508 9518 9536 9551
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 9508 9178 9536 9454
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9402 8800 9458 8809
rect 9402 8735 9458 8744
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9324 3738 9352 4014
rect 9416 3942 9444 8735
rect 9508 8634 9536 9114
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9600 7834 9628 9862
rect 9678 9480 9734 9489
rect 9678 9415 9680 9424
rect 9732 9415 9734 9424
rect 9680 9386 9732 9392
rect 9784 9178 9812 25094
rect 9862 23216 9918 23225
rect 9862 23151 9918 23160
rect 9876 22234 9904 23151
rect 10060 22574 10088 26415
rect 10152 24721 10180 27520
rect 10796 26246 10824 27520
rect 11348 26625 11376 27520
rect 11334 26616 11390 26625
rect 11334 26551 11390 26560
rect 11610 26616 11666 26625
rect 11610 26551 11666 26560
rect 10784 26240 10836 26246
rect 10784 26182 10836 26188
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10232 24812 10284 24818
rect 10232 24754 10284 24760
rect 10138 24712 10194 24721
rect 10138 24647 10194 24656
rect 10244 24596 10272 24754
rect 10152 24568 10272 24596
rect 10152 24274 10180 24568
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10140 24268 10192 24274
rect 10140 24210 10192 24216
rect 10152 24070 10180 24210
rect 10416 24200 10468 24206
rect 10416 24142 10468 24148
rect 10690 24168 10746 24177
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 10324 24064 10376 24070
rect 10324 24006 10376 24012
rect 10152 23526 10180 24006
rect 10336 23730 10364 24006
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10428 23594 10456 24142
rect 10690 24103 10746 24112
rect 10416 23588 10468 23594
rect 10416 23530 10468 23536
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 10152 22710 10180 23462
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10324 23112 10376 23118
rect 10324 23054 10376 23060
rect 10336 22778 10364 23054
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10140 22704 10192 22710
rect 10704 22681 10732 24103
rect 10796 23905 10824 26182
rect 11520 26104 11572 26110
rect 11520 26046 11572 26052
rect 10876 26036 10928 26042
rect 10876 25978 10928 25984
rect 10782 23896 10838 23905
rect 10782 23831 10838 23840
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10796 23089 10824 23462
rect 10888 23202 10916 25978
rect 11336 25832 11388 25838
rect 11336 25774 11388 25780
rect 11348 25362 11376 25774
rect 11336 25356 11388 25362
rect 11336 25298 11388 25304
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 11072 24886 11100 25230
rect 11532 24886 11560 26046
rect 11060 24880 11112 24886
rect 11058 24848 11060 24857
rect 11520 24880 11572 24886
rect 11112 24848 11114 24857
rect 11058 24783 11114 24792
rect 11426 24848 11482 24857
rect 11520 24822 11572 24828
rect 11426 24783 11482 24792
rect 11440 24614 11468 24783
rect 11428 24608 11480 24614
rect 11428 24550 11480 24556
rect 11426 24304 11482 24313
rect 11426 24239 11482 24248
rect 11440 24206 11468 24239
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 10966 24032 11022 24041
rect 10966 23967 11022 23976
rect 10980 23798 11008 23967
rect 10968 23792 11020 23798
rect 10968 23734 11020 23740
rect 11334 23760 11390 23769
rect 10980 23322 11008 23734
rect 11334 23695 11390 23704
rect 11152 23520 11204 23526
rect 11152 23462 11204 23468
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 11058 23216 11114 23225
rect 10888 23174 11008 23202
rect 10782 23080 10838 23089
rect 10782 23015 10838 23024
rect 10140 22646 10192 22652
rect 10690 22672 10746 22681
rect 10690 22607 10746 22616
rect 10048 22568 10100 22574
rect 10048 22510 10100 22516
rect 9956 22500 10008 22506
rect 9956 22442 10008 22448
rect 9864 22228 9916 22234
rect 9864 22170 9916 22176
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 9876 21010 9904 21490
rect 9864 21004 9916 21010
rect 9864 20946 9916 20952
rect 9876 20466 9904 20946
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 9876 19718 9904 20402
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9968 18358 9996 22442
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 10060 22166 10088 22374
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10704 22234 10732 22607
rect 10784 22500 10836 22506
rect 10784 22442 10836 22448
rect 10692 22228 10744 22234
rect 10692 22170 10744 22176
rect 10048 22160 10100 22166
rect 10048 22102 10100 22108
rect 10060 20777 10088 22102
rect 10140 21888 10192 21894
rect 10140 21830 10192 21836
rect 10152 21350 10180 21830
rect 10704 21418 10732 22170
rect 10692 21412 10744 21418
rect 10692 21354 10744 21360
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 10152 20913 10180 21286
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10690 21040 10746 21049
rect 10690 20975 10746 20984
rect 10138 20904 10194 20913
rect 10138 20839 10194 20848
rect 10046 20768 10102 20777
rect 10046 20703 10102 20712
rect 10048 20256 10100 20262
rect 10046 20224 10048 20233
rect 10100 20224 10102 20233
rect 10046 20159 10102 20168
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 10060 18970 10088 19110
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 9956 18352 10008 18358
rect 9956 18294 10008 18300
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9968 16794 9996 17070
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9954 16416 10010 16425
rect 10060 16402 10088 18906
rect 10010 16374 10088 16402
rect 9954 16351 10010 16360
rect 9862 15872 9918 15881
rect 9862 15807 9918 15816
rect 9876 15638 9904 15807
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 9968 14498 9996 16351
rect 10152 15094 10180 19994
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10704 18873 10732 20975
rect 10796 20641 10824 22442
rect 10876 21344 10928 21350
rect 10876 21286 10928 21292
rect 10782 20632 10838 20641
rect 10782 20567 10838 20576
rect 10784 20324 10836 20330
rect 10784 20266 10836 20272
rect 10796 20058 10824 20266
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10784 19780 10836 19786
rect 10784 19722 10836 19728
rect 10796 19310 10824 19722
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10690 18864 10746 18873
rect 10796 18834 10824 19246
rect 10690 18799 10746 18808
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10796 18426 10824 18770
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10888 18034 10916 21286
rect 10704 18006 10916 18034
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10336 16250 10364 16594
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10704 15688 10732 18006
rect 10874 17912 10930 17921
rect 10874 17847 10876 17856
rect 10928 17847 10930 17856
rect 10876 17818 10928 17824
rect 10980 16402 11008 23174
rect 11058 23151 11060 23160
rect 11112 23151 11114 23160
rect 11060 23122 11112 23128
rect 11072 22778 11100 23122
rect 11164 22953 11192 23462
rect 11242 23080 11298 23089
rect 11242 23015 11298 23024
rect 11150 22944 11206 22953
rect 11150 22879 11206 22888
rect 11256 22817 11284 23015
rect 11242 22808 11298 22817
rect 11060 22772 11112 22778
rect 11242 22743 11298 22752
rect 11060 22714 11112 22720
rect 11060 22636 11112 22642
rect 11060 22578 11112 22584
rect 11072 22030 11100 22578
rect 11244 22568 11296 22574
rect 11244 22510 11296 22516
rect 11060 22024 11112 22030
rect 11112 21984 11192 22012
rect 11060 21966 11112 21972
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 11072 21049 11100 21626
rect 11164 21486 11192 21984
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 11058 21040 11114 21049
rect 11058 20975 11114 20984
rect 11072 20058 11100 20975
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11164 19786 11192 21422
rect 11256 20641 11284 22510
rect 11348 22386 11376 23695
rect 11426 23216 11482 23225
rect 11426 23151 11482 23160
rect 11440 22778 11468 23151
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11532 22556 11560 24822
rect 11624 24585 11652 26551
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 11716 25498 11744 25842
rect 11704 25492 11756 25498
rect 11704 25434 11756 25440
rect 11610 24576 11666 24585
rect 11610 24511 11666 24520
rect 11610 24304 11666 24313
rect 11610 24239 11666 24248
rect 11624 23633 11652 24239
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11704 23792 11756 23798
rect 11704 23734 11756 23740
rect 11610 23624 11666 23633
rect 11610 23559 11666 23568
rect 11532 22528 11652 22556
rect 11348 22358 11560 22386
rect 11336 22092 11388 22098
rect 11336 22034 11388 22040
rect 11348 21690 11376 22034
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 11428 21072 11480 21078
rect 11428 21014 11480 21020
rect 11242 20632 11298 20641
rect 11242 20567 11298 20576
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11152 19780 11204 19786
rect 11152 19722 11204 19728
rect 11256 19378 11284 19790
rect 11244 19372 11296 19378
rect 11244 19314 11296 19320
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 11072 18970 11100 19110
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 11256 18902 11284 19314
rect 11244 18896 11296 18902
rect 11244 18838 11296 18844
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 11072 18057 11100 18158
rect 11058 18048 11114 18057
rect 11058 17983 11114 17992
rect 11164 17882 11192 18362
rect 11256 18290 11284 18838
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11244 18284 11296 18290
rect 11244 18226 11296 18232
rect 11348 18086 11376 18770
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11256 17921 11284 18022
rect 11242 17912 11298 17921
rect 11152 17876 11204 17882
rect 11072 17836 11152 17864
rect 11072 17202 11100 17836
rect 11242 17847 11298 17856
rect 11152 17818 11204 17824
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11164 17338 11192 17614
rect 11242 17368 11298 17377
rect 11152 17332 11204 17338
rect 11348 17354 11376 18022
rect 11298 17326 11376 17354
rect 11242 17303 11298 17312
rect 11152 17274 11204 17280
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 11164 16726 11192 17274
rect 11256 17270 11284 17303
rect 11244 17264 11296 17270
rect 11244 17206 11296 17212
rect 11152 16720 11204 16726
rect 11152 16662 11204 16668
rect 10612 15660 10732 15688
rect 10796 16374 11008 16402
rect 10140 15088 10192 15094
rect 10140 15030 10192 15036
rect 10612 14958 10640 15660
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 9876 14470 9996 14498
rect 9876 13138 9904 14470
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9968 13433 9996 14350
rect 10060 13802 10088 14758
rect 10152 14618 10180 14894
rect 10704 14822 10732 15506
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 9954 13424 10010 13433
rect 9954 13359 10010 13368
rect 10060 13258 10088 13738
rect 10152 13530 10180 14554
rect 10598 14512 10654 14521
rect 10598 14447 10654 14456
rect 10612 14278 10640 14447
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10704 13734 10732 14758
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10230 13424 10286 13433
rect 10230 13359 10286 13368
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 9876 13110 10180 13138
rect 10046 12880 10102 12889
rect 10046 12815 10102 12824
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9692 8401 9720 8978
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9678 8392 9734 8401
rect 9678 8327 9734 8336
rect 9784 8294 9812 8910
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9508 7806 9628 7834
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9508 6730 9536 7806
rect 9588 7744 9640 7750
rect 9640 7704 9720 7732
rect 9588 7686 9640 7692
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9508 4865 9536 4966
rect 9494 4856 9550 4865
rect 9494 4791 9550 4800
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9508 4214 9536 4422
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9494 3632 9550 3641
rect 9494 3567 9550 3576
rect 9218 2680 9274 2689
rect 8864 2638 8984 2666
rect 8666 2544 8722 2553
rect 8666 2479 8722 2488
rect 8956 480 8984 2638
rect 9218 2615 9274 2624
rect 9508 480 9536 3567
rect 9600 3369 9628 7210
rect 9692 7206 9720 7704
rect 9784 7410 9812 7822
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 4826 9720 7142
rect 9784 7002 9812 7346
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9784 4457 9812 6598
rect 9770 4448 9826 4457
rect 9770 4383 9826 4392
rect 9678 4176 9734 4185
rect 9678 4111 9734 4120
rect 9692 3738 9720 4111
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9876 3602 9904 12242
rect 9968 12170 9996 12718
rect 10060 12646 10088 12815
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10060 12442 10088 12582
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 9954 12064 10010 12073
rect 9954 11999 10010 12008
rect 9968 6662 9996 11999
rect 10060 8634 10088 12242
rect 10152 11257 10180 13110
rect 10244 12986 10272 13359
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 10612 12850 10640 13262
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10138 11248 10194 11257
rect 10138 11183 10194 11192
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10428 10810 10456 11154
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10336 9926 10364 10066
rect 10324 9920 10376 9926
rect 10138 9888 10194 9897
rect 10612 9897 10640 10066
rect 10324 9862 10376 9868
rect 10598 9888 10654 9897
rect 10138 9823 10194 9832
rect 10152 9178 10180 9823
rect 10336 9450 10364 9862
rect 10598 9823 10654 9832
rect 10598 9752 10654 9761
rect 10598 9687 10654 9696
rect 10612 9489 10640 9687
rect 10598 9480 10654 9489
rect 10324 9444 10376 9450
rect 10598 9415 10654 9424
rect 10324 9386 10376 9392
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10600 8492 10652 8498
rect 10704 8480 10732 12922
rect 10796 12617 10824 16374
rect 11164 16250 11192 16662
rect 11242 16552 11298 16561
rect 11242 16487 11298 16496
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 10888 15570 10916 16186
rect 11256 16046 11284 16487
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 10968 15972 11020 15978
rect 11020 15932 11100 15960
rect 10968 15914 11020 15920
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10888 15162 10916 15506
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10874 15056 10930 15065
rect 11072 15026 11100 15932
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 10874 14991 10930 15000
rect 11060 15020 11112 15026
rect 10888 14618 10916 14991
rect 11060 14962 11112 14968
rect 11164 14822 11192 15574
rect 11334 15192 11390 15201
rect 11334 15127 11390 15136
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 10966 14648 11022 14657
rect 10876 14612 10928 14618
rect 11256 14634 11284 15030
rect 10966 14583 11022 14592
rect 11164 14606 11284 14634
rect 10876 14554 10928 14560
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10888 14074 10916 14350
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10980 13841 11008 14583
rect 10966 13832 11022 13841
rect 10966 13767 11022 13776
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 10874 13560 10930 13569
rect 10874 13495 10930 13504
rect 10888 13394 10916 13495
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10782 12608 10838 12617
rect 10782 12543 10838 12552
rect 10874 12336 10930 12345
rect 10980 12322 11008 13670
rect 11072 12442 11100 13670
rect 11164 13410 11192 14606
rect 11244 14408 11296 14414
rect 11242 14376 11244 14385
rect 11296 14376 11298 14385
rect 11242 14311 11298 14320
rect 11348 14249 11376 15127
rect 11334 14240 11390 14249
rect 11334 14175 11390 14184
rect 11440 14090 11468 21014
rect 11532 20058 11560 22358
rect 11624 20398 11652 22528
rect 11716 22137 11744 23734
rect 11808 23730 11836 24006
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 11900 23633 11928 27520
rect 12072 25356 12124 25362
rect 12072 25298 12124 25304
rect 11980 25152 12032 25158
rect 11980 25094 12032 25100
rect 11886 23624 11942 23633
rect 11886 23559 11942 23568
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 11808 22710 11836 23054
rect 11796 22704 11848 22710
rect 11796 22646 11848 22652
rect 11900 22438 11928 23122
rect 11992 22574 12020 25094
rect 12084 24070 12112 25298
rect 12440 25152 12492 25158
rect 12440 25094 12492 25100
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 12268 24614 12296 24754
rect 12348 24744 12400 24750
rect 12452 24698 12480 25094
rect 12400 24692 12480 24698
rect 12348 24686 12480 24692
rect 12360 24670 12480 24686
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 12164 24200 12216 24206
rect 12164 24142 12216 24148
rect 12072 24064 12124 24070
rect 12072 24006 12124 24012
rect 12084 22817 12112 24006
rect 12176 23866 12204 24142
rect 12164 23860 12216 23866
rect 12164 23802 12216 23808
rect 12268 23712 12296 24550
rect 12452 24041 12480 24670
rect 12544 24562 12572 27520
rect 13096 25514 13124 27520
rect 13544 26512 13596 26518
rect 13544 26454 13596 26460
rect 12808 25492 12860 25498
rect 12808 25434 12860 25440
rect 12900 25492 12952 25498
rect 13096 25486 13400 25514
rect 12900 25434 12952 25440
rect 12716 24608 12768 24614
rect 12544 24534 12664 24562
rect 12716 24550 12768 24556
rect 12530 24440 12586 24449
rect 12530 24375 12586 24384
rect 12438 24032 12494 24041
rect 12438 23967 12494 23976
rect 12544 23746 12572 24375
rect 12176 23684 12296 23712
rect 12452 23718 12572 23746
rect 12070 22808 12126 22817
rect 12070 22743 12126 22752
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11900 22137 11928 22374
rect 11702 22128 11758 22137
rect 11702 22063 11758 22072
rect 11886 22128 11942 22137
rect 11886 22063 11942 22072
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 11796 21412 11848 21418
rect 11796 21354 11848 21360
rect 11808 21146 11836 21354
rect 11796 21140 11848 21146
rect 11796 21082 11848 21088
rect 11612 20392 11664 20398
rect 11612 20334 11664 20340
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11532 19446 11560 19994
rect 11900 19922 11928 21626
rect 12084 20874 12112 22743
rect 12072 20868 12124 20874
rect 12072 20810 12124 20816
rect 12070 20360 12126 20369
rect 11980 20324 12032 20330
rect 12070 20295 12126 20304
rect 11980 20266 12032 20272
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11704 19848 11756 19854
rect 11702 19816 11704 19825
rect 11756 19816 11758 19825
rect 11702 19751 11758 19760
rect 11520 19440 11572 19446
rect 11520 19382 11572 19388
rect 11900 19378 11928 19858
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11520 18284 11572 18290
rect 11520 18226 11572 18232
rect 11532 17882 11560 18226
rect 11612 18216 11664 18222
rect 11612 18158 11664 18164
rect 11520 17876 11572 17882
rect 11520 17818 11572 17824
rect 11518 15464 11574 15473
rect 11518 15399 11574 15408
rect 11348 14062 11468 14090
rect 11242 13832 11298 13841
rect 11242 13767 11298 13776
rect 11256 13530 11284 13767
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11164 13382 11284 13410
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 13025 11192 13126
rect 11150 13016 11206 13025
rect 11256 12986 11284 13382
rect 11150 12951 11206 12960
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11244 12776 11296 12782
rect 11150 12744 11206 12753
rect 11244 12718 11296 12724
rect 11150 12679 11206 12688
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 10980 12294 11100 12322
rect 10874 12271 10876 12280
rect 10928 12271 10930 12280
rect 10876 12242 10928 12248
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10874 12200 10930 12209
rect 10796 11393 10824 12174
rect 10874 12135 10930 12144
rect 10888 11665 10916 12135
rect 10874 11656 10930 11665
rect 10874 11591 10930 11600
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10782 11384 10838 11393
rect 10782 11319 10838 11328
rect 10888 11286 10916 11494
rect 10876 11280 10928 11286
rect 10782 11248 10838 11257
rect 10876 11222 10928 11228
rect 10782 11183 10838 11192
rect 10652 8452 10732 8480
rect 10600 8434 10652 8440
rect 10060 6746 10088 8434
rect 10796 8362 10824 11183
rect 10888 10606 10916 11222
rect 10966 11112 11022 11121
rect 10966 11047 11022 11056
rect 10980 10674 11008 11047
rect 11072 10713 11100 12294
rect 11058 10704 11114 10713
rect 10968 10668 11020 10674
rect 11058 10639 11114 10648
rect 10968 10610 11020 10616
rect 10876 10600 10928 10606
rect 10928 10548 11008 10554
rect 10876 10542 11008 10548
rect 10888 10526 11008 10542
rect 10876 10464 10928 10470
rect 10874 10432 10876 10441
rect 10928 10432 10930 10441
rect 10874 10367 10930 10376
rect 10888 10266 10916 10367
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10980 10062 11008 10526
rect 11058 10296 11114 10305
rect 11164 10266 11192 12679
rect 11058 10231 11114 10240
rect 11152 10260 11204 10266
rect 11072 10198 11100 10231
rect 11152 10202 11204 10208
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10980 9897 11008 9998
rect 10966 9888 11022 9897
rect 10966 9823 11022 9832
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10690 8256 10746 8265
rect 10289 8188 10585 8208
rect 10690 8191 10746 8200
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 8090 10732 8191
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10784 8016 10836 8022
rect 10888 8004 10916 9658
rect 10980 9178 11008 9823
rect 11072 9722 11100 10134
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 11072 9217 11100 9386
rect 11058 9208 11114 9217
rect 10968 9172 11020 9178
rect 11058 9143 11114 9152
rect 10968 9114 11020 9120
rect 10980 8498 11008 9114
rect 11058 8528 11114 8537
rect 10968 8492 11020 8498
rect 11058 8463 11114 8472
rect 10968 8434 11020 8440
rect 10836 7976 10916 8004
rect 10968 8016 11020 8022
rect 10784 7958 10836 7964
rect 10968 7958 11020 7964
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10888 7546 10916 7822
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10416 6928 10468 6934
rect 10416 6870 10468 6876
rect 10428 6769 10456 6870
rect 10051 6718 10088 6746
rect 10414 6760 10470 6769
rect 9956 6656 10008 6662
rect 10051 6644 10079 6718
rect 10414 6695 10470 6704
rect 10598 6760 10654 6769
rect 10598 6695 10654 6704
rect 10140 6656 10192 6662
rect 10051 6616 10088 6644
rect 9956 6598 10008 6604
rect 9954 6488 10010 6497
rect 9954 6423 9956 6432
rect 10008 6423 10010 6432
rect 9956 6394 10008 6400
rect 9954 6216 10010 6225
rect 9954 6151 10010 6160
rect 9968 6118 9996 6151
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9968 5846 9996 6054
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 9968 4758 9996 5782
rect 9956 4752 10008 4758
rect 9956 4694 10008 4700
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9586 3360 9642 3369
rect 9586 3295 9642 3304
rect 9770 3360 9826 3369
rect 9770 3295 9826 3304
rect 9600 2281 9628 3295
rect 9784 2990 9812 3295
rect 9876 3194 9904 3538
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9784 2854 9812 2885
rect 9772 2848 9824 2854
rect 9770 2816 9772 2825
rect 9824 2816 9826 2825
rect 9770 2751 9826 2760
rect 9586 2272 9642 2281
rect 9586 2207 9642 2216
rect 9784 1057 9812 2751
rect 9770 1048 9826 1057
rect 9770 983 9826 992
rect 10060 480 10088 6616
rect 10140 6598 10192 6604
rect 10152 3738 10180 6598
rect 10506 6488 10562 6497
rect 10612 6458 10640 6695
rect 10506 6423 10562 6432
rect 10600 6452 10652 6458
rect 10520 6390 10548 6423
rect 10600 6394 10652 6400
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10322 5536 10378 5545
rect 10322 5471 10378 5480
rect 10506 5536 10562 5545
rect 10506 5471 10562 5480
rect 10336 5098 10364 5471
rect 10520 5370 10548 5471
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10888 5234 10916 7482
rect 10980 7274 11008 7958
rect 11072 7274 11100 8463
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11164 7342 11192 8026
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 10980 7177 11008 7210
rect 10966 7168 11022 7177
rect 10966 7103 11022 7112
rect 11256 6984 11284 12718
rect 11348 10146 11376 14062
rect 11532 13462 11560 15399
rect 11624 13530 11652 18158
rect 11704 17060 11756 17066
rect 11704 17002 11756 17008
rect 11716 16454 11744 17002
rect 11886 16552 11942 16561
rect 11886 16487 11942 16496
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11716 16114 11744 16390
rect 11900 16250 11928 16487
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11794 15600 11850 15609
rect 11794 15535 11850 15544
rect 11808 15337 11836 15535
rect 11794 15328 11850 15337
rect 11794 15263 11850 15272
rect 11992 15178 12020 20266
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11808 15150 12020 15178
rect 11716 14482 11744 15098
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11716 14006 11744 14418
rect 11704 14000 11756 14006
rect 11704 13942 11756 13948
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11440 12442 11468 13262
rect 11624 12986 11652 13466
rect 11702 13288 11758 13297
rect 11702 13223 11758 13232
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11624 12753 11652 12922
rect 11610 12744 11666 12753
rect 11610 12679 11666 12688
rect 11518 12472 11574 12481
rect 11428 12436 11480 12442
rect 11716 12442 11744 13223
rect 11518 12407 11574 12416
rect 11704 12436 11756 12442
rect 11428 12378 11480 12384
rect 11426 11928 11482 11937
rect 11426 11863 11482 11872
rect 11440 11257 11468 11863
rect 11426 11248 11482 11257
rect 11426 11183 11482 11192
rect 11348 10118 11468 10146
rect 11334 10024 11390 10033
rect 11334 9959 11336 9968
rect 11388 9959 11390 9968
rect 11336 9930 11388 9936
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11348 7206 11376 9590
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11072 6956 11284 6984
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10874 5128 10930 5137
rect 10324 5092 10376 5098
rect 10874 5063 10930 5072
rect 10324 5034 10376 5040
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10888 4826 10916 5063
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10324 4480 10376 4486
rect 10322 4448 10324 4457
rect 10376 4448 10378 4457
rect 10322 4383 10378 4392
rect 10796 3942 10824 4626
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10152 3126 10180 3674
rect 10796 3233 10824 3878
rect 10888 3738 10916 4762
rect 11072 4321 11100 6956
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11164 6322 11192 6802
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11164 5914 11192 6258
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11164 5234 11192 5850
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11164 4622 11192 5170
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11152 4616 11204 4622
rect 11204 4576 11284 4604
rect 11152 4558 11204 4564
rect 11058 4312 11114 4321
rect 11058 4247 11114 4256
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10782 3224 10838 3233
rect 10782 3159 10838 3168
rect 10876 3188 10928 3194
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10690 2680 10746 2689
rect 10612 2624 10690 2632
rect 10612 2615 10746 2624
rect 10612 2604 10732 2615
rect 10612 2417 10640 2604
rect 10796 2417 10824 3159
rect 10876 3130 10928 3136
rect 10888 2582 10916 3130
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 10598 2408 10654 2417
rect 10598 2343 10654 2352
rect 10782 2408 10838 2417
rect 10782 2343 10838 2352
rect 10980 2009 11008 3878
rect 10966 2000 11022 2009
rect 10966 1935 11022 1944
rect 11072 1737 11100 4014
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11164 3194 11192 3674
rect 11256 3602 11284 4576
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11242 3088 11298 3097
rect 11152 3052 11204 3058
rect 11242 3023 11298 3032
rect 11152 2994 11204 3000
rect 11058 1728 11114 1737
rect 11058 1663 11114 1672
rect 10598 1184 10654 1193
rect 10598 1119 10654 1128
rect 10612 480 10640 1119
rect 11164 480 11192 2994
rect 11256 2990 11284 3023
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11242 2544 11298 2553
rect 11242 2479 11298 2488
rect 11256 2310 11284 2479
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 11256 1737 11284 2246
rect 11348 2106 11376 4966
rect 11440 3058 11468 10118
rect 11532 9654 11560 12407
rect 11704 12378 11756 12384
rect 11702 12336 11758 12345
rect 11702 12271 11758 12280
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11624 10810 11652 11290
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11610 10296 11666 10305
rect 11610 10231 11666 10240
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11532 7750 11560 8230
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11624 6934 11652 10231
rect 11612 6928 11664 6934
rect 11612 6870 11664 6876
rect 11518 5264 11574 5273
rect 11518 5199 11574 5208
rect 11532 5098 11560 5199
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11532 4826 11560 5034
rect 11610 4856 11666 4865
rect 11520 4820 11572 4826
rect 11610 4791 11666 4800
rect 11520 4762 11572 4768
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11532 4049 11560 4082
rect 11518 4040 11574 4049
rect 11518 3975 11574 3984
rect 11624 3670 11652 4791
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 11624 2854 11652 3470
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11336 2100 11388 2106
rect 11336 2042 11388 2048
rect 11242 1728 11298 1737
rect 11242 1663 11298 1672
rect 11440 1193 11468 2790
rect 11426 1184 11482 1193
rect 11426 1119 11482 1128
rect 11716 480 11744 12271
rect 11808 9194 11836 15150
rect 11978 14240 12034 14249
rect 11978 14175 12034 14184
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11900 12714 11928 13330
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11900 12345 11928 12650
rect 11886 12336 11942 12345
rect 11886 12271 11942 12280
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11900 11558 11928 12174
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11900 11218 11928 11494
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11886 10840 11942 10849
rect 11886 10775 11888 10784
rect 11940 10775 11942 10784
rect 11888 10746 11940 10752
rect 11992 10266 12020 14175
rect 12084 13161 12112 20295
rect 12176 18057 12204 23684
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12360 22760 12388 23598
rect 12452 23497 12480 23718
rect 12532 23588 12584 23594
rect 12532 23530 12584 23536
rect 12438 23488 12494 23497
rect 12438 23423 12494 23432
rect 12544 23322 12572 23530
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12440 22772 12492 22778
rect 12360 22732 12440 22760
rect 12440 22714 12492 22720
rect 12544 21962 12572 23258
rect 12532 21956 12584 21962
rect 12532 21898 12584 21904
rect 12636 21690 12664 24534
rect 12728 22574 12756 24550
rect 12820 23254 12848 25434
rect 12912 25294 12940 25434
rect 12900 25288 12952 25294
rect 12900 25230 12952 25236
rect 13084 25288 13136 25294
rect 13084 25230 13136 25236
rect 12992 25152 13044 25158
rect 12992 25094 13044 25100
rect 13004 24886 13032 25094
rect 13096 24954 13124 25230
rect 13176 25152 13228 25158
rect 13176 25094 13228 25100
rect 13084 24948 13136 24954
rect 13084 24890 13136 24896
rect 12992 24880 13044 24886
rect 12992 24822 13044 24828
rect 12990 24712 13046 24721
rect 12990 24647 13046 24656
rect 13004 24274 13032 24647
rect 12992 24268 13044 24274
rect 12992 24210 13044 24216
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12808 23248 12860 23254
rect 12808 23190 12860 23196
rect 12912 23186 12940 24006
rect 12900 23180 12952 23186
rect 12900 23122 12952 23128
rect 12808 22976 12860 22982
rect 12806 22944 12808 22953
rect 12860 22944 12862 22953
rect 12806 22879 12862 22888
rect 12912 22642 12940 23122
rect 13004 23050 13032 24210
rect 13096 23322 13124 24890
rect 13084 23316 13136 23322
rect 13084 23258 13136 23264
rect 13096 23050 13124 23258
rect 12992 23044 13044 23050
rect 12992 22986 13044 22992
rect 13084 23044 13136 23050
rect 13084 22986 13136 22992
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12728 22166 12756 22510
rect 13004 22273 13032 22986
rect 13188 22658 13216 25094
rect 13372 24313 13400 25486
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13464 24614 13492 24754
rect 13452 24608 13504 24614
rect 13452 24550 13504 24556
rect 13358 24304 13414 24313
rect 13358 24239 13414 24248
rect 13464 24206 13492 24550
rect 13360 24200 13412 24206
rect 13360 24142 13412 24148
rect 13452 24200 13504 24206
rect 13452 24142 13504 24148
rect 13372 23769 13400 24142
rect 13358 23760 13414 23769
rect 13358 23695 13414 23704
rect 13464 23594 13492 24142
rect 13452 23588 13504 23594
rect 13452 23530 13504 23536
rect 13360 23112 13412 23118
rect 13360 23054 13412 23060
rect 13372 22710 13400 23054
rect 13452 23044 13504 23050
rect 13452 22986 13504 22992
rect 13096 22630 13216 22658
rect 13360 22704 13412 22710
rect 13360 22646 13412 22652
rect 12990 22264 13046 22273
rect 12990 22199 13046 22208
rect 12716 22160 12768 22166
rect 12716 22102 12768 22108
rect 12808 21956 12860 21962
rect 12808 21898 12860 21904
rect 12820 21690 12848 21898
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 12254 21584 12310 21593
rect 12254 21519 12310 21528
rect 12268 21146 12296 21519
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12714 21040 12770 21049
rect 12624 21004 12676 21010
rect 12714 20975 12716 20984
rect 12624 20946 12676 20952
rect 12768 20975 12770 20984
rect 12990 21040 13046 21049
rect 12990 20975 13046 20984
rect 12716 20946 12768 20952
rect 12256 20868 12308 20874
rect 12256 20810 12308 20816
rect 12268 19242 12296 20810
rect 12636 20602 12664 20946
rect 12900 20936 12952 20942
rect 12806 20904 12862 20913
rect 12900 20878 12952 20884
rect 12806 20839 12862 20848
rect 12624 20596 12676 20602
rect 12624 20538 12676 20544
rect 12820 19922 12848 20839
rect 12912 20602 12940 20878
rect 12900 20596 12952 20602
rect 12900 20538 12952 20544
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 12912 20097 12940 20198
rect 12898 20088 12954 20097
rect 12898 20023 12900 20032
rect 12952 20023 12954 20032
rect 12900 19994 12952 20000
rect 12912 19963 12940 19994
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12728 19514 12756 19790
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 12728 19310 12756 19450
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12256 19236 12308 19242
rect 12256 19178 12308 19184
rect 12624 19236 12676 19242
rect 12624 19178 12676 19184
rect 12636 18442 12664 19178
rect 12820 18970 12848 19858
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12544 18414 12664 18442
rect 12162 18048 12218 18057
rect 12162 17983 12218 17992
rect 12438 18048 12494 18057
rect 12438 17983 12494 17992
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12360 16436 12388 17478
rect 12452 17241 12480 17983
rect 12438 17232 12494 17241
rect 12544 17218 12572 18414
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12636 17490 12664 18226
rect 13004 17882 13032 20975
rect 13096 18222 13124 22630
rect 13360 22568 13412 22574
rect 13360 22510 13412 22516
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 13280 21554 13308 21830
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 13280 18970 13308 19314
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 13372 18902 13400 22510
rect 13464 22438 13492 22986
rect 13556 22574 13584 26454
rect 13648 23730 13676 27520
rect 13910 25528 13966 25537
rect 13910 25463 13966 25472
rect 14188 25492 14240 25498
rect 13924 24313 13952 25463
rect 14188 25434 14240 25440
rect 14096 25424 14148 25430
rect 14096 25366 14148 25372
rect 14004 25288 14056 25294
rect 14004 25230 14056 25236
rect 14016 24818 14044 25230
rect 14108 24954 14136 25366
rect 14096 24948 14148 24954
rect 14096 24890 14148 24896
rect 14004 24812 14056 24818
rect 14004 24754 14056 24760
rect 13910 24304 13966 24313
rect 13910 24239 13966 24248
rect 14016 24138 14044 24754
rect 14200 24342 14228 25434
rect 14292 24857 14320 27520
rect 14844 26353 14872 27520
rect 14830 26344 14886 26353
rect 14830 26279 14886 26288
rect 14462 26072 14518 26081
rect 14462 26007 14518 26016
rect 14646 26072 14702 26081
rect 14646 26007 14702 26016
rect 14476 25537 14504 26007
rect 14462 25528 14518 25537
rect 14462 25463 14518 25472
rect 14372 25356 14424 25362
rect 14372 25298 14424 25304
rect 14278 24848 14334 24857
rect 14278 24783 14334 24792
rect 14384 24750 14412 25298
rect 14660 25129 14688 26007
rect 14832 25152 14884 25158
rect 14646 25120 14702 25129
rect 14832 25094 14884 25100
rect 15292 25152 15344 25158
rect 15292 25094 15344 25100
rect 14646 25055 14702 25064
rect 14844 24818 14872 25094
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15106 24848 15162 24857
rect 14832 24812 14884 24818
rect 15106 24783 15162 24792
rect 14832 24754 14884 24760
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14464 24744 14516 24750
rect 14464 24686 14516 24692
rect 14188 24336 14240 24342
rect 14188 24278 14240 24284
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14004 24132 14056 24138
rect 14004 24074 14056 24080
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13544 22568 13596 22574
rect 13544 22510 13596 22516
rect 13452 22432 13504 22438
rect 13452 22374 13504 22380
rect 13544 22432 13596 22438
rect 13544 22374 13596 22380
rect 13464 21078 13492 22374
rect 13556 22234 13584 22374
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13648 21865 13676 23666
rect 13740 23322 13768 24006
rect 13912 23588 13964 23594
rect 13912 23530 13964 23536
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 13728 23316 13780 23322
rect 13728 23258 13780 23264
rect 13740 22438 13768 23258
rect 13832 23118 13860 23462
rect 13924 23322 13952 23530
rect 14004 23520 14056 23526
rect 14004 23462 14056 23468
rect 13912 23316 13964 23322
rect 13912 23258 13964 23264
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13728 22432 13780 22438
rect 13728 22374 13780 22380
rect 14016 22250 14044 23462
rect 13832 22222 14044 22250
rect 13634 21856 13690 21865
rect 13634 21791 13690 21800
rect 13634 21176 13690 21185
rect 13634 21111 13636 21120
rect 13688 21111 13690 21120
rect 13636 21082 13688 21088
rect 13452 21072 13504 21078
rect 13452 21014 13504 21020
rect 13832 20398 13860 22222
rect 13912 22160 13964 22166
rect 13912 22102 13964 22108
rect 13924 21185 13952 22102
rect 14004 22024 14056 22030
rect 14002 21992 14004 22001
rect 14056 21992 14058 22001
rect 14002 21927 14058 21936
rect 14016 21690 14044 21927
rect 14004 21684 14056 21690
rect 14004 21626 14056 21632
rect 14004 21412 14056 21418
rect 14004 21354 14056 21360
rect 13910 21176 13966 21185
rect 13910 21111 13966 21120
rect 14016 20806 14044 21354
rect 14004 20800 14056 20806
rect 14004 20742 14056 20748
rect 13910 20632 13966 20641
rect 13910 20567 13966 20576
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 13450 20088 13506 20097
rect 13450 20023 13506 20032
rect 13360 18896 13412 18902
rect 13360 18838 13412 18844
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12636 17462 12848 17490
rect 12544 17190 12756 17218
rect 12438 17167 12494 17176
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12544 16658 12572 17002
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12360 16408 12480 16436
rect 12346 16280 12402 16289
rect 12346 16215 12348 16224
rect 12400 16215 12402 16224
rect 12348 16186 12400 16192
rect 12452 15978 12480 16408
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12162 15736 12218 15745
rect 12162 15671 12164 15680
rect 12216 15671 12218 15680
rect 12164 15642 12216 15648
rect 12176 14550 12204 15642
rect 12544 15314 12572 16594
rect 12452 15286 12572 15314
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 12176 13938 12204 14486
rect 12268 14074 12296 14758
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12268 13326 12296 14010
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12070 13152 12126 13161
rect 12070 13087 12126 13096
rect 12084 12617 12112 13087
rect 12070 12608 12126 12617
rect 12070 12543 12126 12552
rect 12070 12472 12126 12481
rect 12070 12407 12126 12416
rect 12256 12436 12308 12442
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11808 9166 11928 9194
rect 11796 9104 11848 9110
rect 11796 9046 11848 9052
rect 11808 8294 11836 9046
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11808 7410 11836 8230
rect 11900 7546 11928 9166
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11808 7002 11836 7346
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11808 6730 11836 6938
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11808 5710 11836 6054
rect 11888 5840 11940 5846
rect 11886 5808 11888 5817
rect 11940 5808 11942 5817
rect 11992 5778 12020 8978
rect 12084 8634 12112 12407
rect 12256 12378 12308 12384
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12176 11354 12204 12242
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12176 10169 12204 10950
rect 12162 10160 12218 10169
rect 12162 10095 12218 10104
rect 12268 9926 12296 12378
rect 12360 10538 12388 14214
rect 12452 11014 12480 15286
rect 12636 14929 12664 16730
rect 12622 14920 12678 14929
rect 12622 14855 12678 14864
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12544 14074 12572 14418
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12440 11008 12492 11014
rect 12544 10985 12572 12922
rect 12440 10950 12492 10956
rect 12530 10976 12586 10985
rect 12452 10826 12480 10950
rect 12530 10911 12586 10920
rect 12530 10840 12586 10849
rect 12452 10798 12530 10826
rect 12530 10775 12586 10784
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 12360 10062 12388 10474
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12452 9466 12480 10406
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12544 9722 12572 9998
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12360 9438 12480 9466
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12070 8528 12126 8537
rect 12070 8463 12126 8472
rect 11886 5743 11942 5752
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11794 3904 11850 3913
rect 11794 3839 11850 3848
rect 11808 3505 11836 3839
rect 11794 3496 11850 3505
rect 11794 3431 11850 3440
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11808 2514 11836 2790
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11900 785 11928 5102
rect 12084 5001 12112 8463
rect 12176 7954 12204 8774
rect 12360 8090 12388 9438
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12452 9217 12480 9318
rect 12438 9208 12494 9217
rect 12438 9143 12494 9152
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12452 7970 12480 8230
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12268 7942 12480 7970
rect 12176 7585 12204 7890
rect 12162 7576 12218 7585
rect 12162 7511 12218 7520
rect 12070 4992 12126 5001
rect 12126 4950 12204 4978
rect 12070 4927 12126 4936
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 12084 4185 12112 4422
rect 12070 4176 12126 4185
rect 12070 4111 12126 4120
rect 11980 3936 12032 3942
rect 12176 3890 12204 4950
rect 11980 3878 12032 3884
rect 11992 2145 12020 3878
rect 12084 3862 12204 3890
rect 12084 3369 12112 3862
rect 12268 3720 12296 7942
rect 12440 7472 12492 7478
rect 12438 7440 12440 7449
rect 12492 7440 12494 7449
rect 12438 7375 12494 7384
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12544 7002 12572 7142
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12544 6662 12572 6938
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 6497 12572 6598
rect 12530 6488 12586 6497
rect 12530 6423 12586 6432
rect 12636 5370 12664 14758
rect 12728 12832 12756 17190
rect 12820 16794 12848 17462
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12912 16726 12940 17682
rect 13096 17377 13124 18022
rect 13082 17368 13138 17377
rect 13004 17326 13082 17354
rect 12900 16720 12952 16726
rect 12900 16662 12952 16668
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12820 16046 12848 16390
rect 12898 16144 12954 16153
rect 12898 16079 12954 16088
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12912 15178 12940 16079
rect 12820 15150 12940 15178
rect 12820 13190 12848 15150
rect 12898 14512 12954 14521
rect 13004 14482 13032 17326
rect 13082 17303 13138 17312
rect 13188 16810 13216 18770
rect 13372 18426 13400 18838
rect 13464 18834 13492 20023
rect 13740 19378 13768 20266
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13832 19242 13860 19722
rect 13820 19236 13872 19242
rect 13820 19178 13872 19184
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13556 18714 13584 19110
rect 13648 18970 13676 19110
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13452 18692 13504 18698
rect 13556 18686 13676 18714
rect 13452 18634 13504 18640
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13096 16782 13216 16810
rect 13096 15858 13124 16782
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 13188 16561 13216 16594
rect 13268 16584 13320 16590
rect 13174 16552 13230 16561
rect 13268 16526 13320 16532
rect 13174 16487 13230 16496
rect 13188 16114 13216 16487
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13096 15830 13216 15858
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13096 14958 13124 15642
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 12898 14447 12954 14456
rect 12992 14476 13044 14482
rect 12912 13870 12940 14447
rect 12992 14418 13044 14424
rect 12990 14376 13046 14385
rect 13096 14362 13124 14894
rect 13188 14822 13216 15830
rect 13280 15638 13308 16526
rect 13372 15706 13400 18362
rect 13464 17882 13492 18634
rect 13648 18630 13676 18686
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13648 18306 13676 18566
rect 13740 18426 13768 18770
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13648 18278 13860 18306
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13464 17338 13492 17614
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13464 16998 13492 17274
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 16590 13492 16934
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13464 16250 13492 16526
rect 13542 16416 13598 16425
rect 13542 16351 13598 16360
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13464 15881 13492 16050
rect 13450 15872 13506 15881
rect 13450 15807 13506 15816
rect 13556 15706 13584 16351
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13450 15600 13506 15609
rect 13450 15535 13506 15544
rect 13464 14958 13492 15535
rect 13544 15496 13596 15502
rect 13542 15464 13544 15473
rect 13596 15464 13598 15473
rect 13542 15399 13598 15408
rect 13556 15042 13584 15399
rect 13648 15201 13676 17682
rect 13740 16810 13768 18158
rect 13832 17882 13860 18278
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13924 17610 13952 20567
rect 14016 19718 14044 20742
rect 14108 20602 14136 24142
rect 14476 24070 14504 24686
rect 14556 24608 14608 24614
rect 14556 24550 14608 24556
rect 14464 24064 14516 24070
rect 14370 24032 14426 24041
rect 14464 24006 14516 24012
rect 14370 23967 14426 23976
rect 14278 23352 14334 23361
rect 14278 23287 14334 23296
rect 14188 22432 14240 22438
rect 14188 22374 14240 22380
rect 14200 21894 14228 22374
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 14186 21720 14242 21729
rect 14186 21655 14242 21664
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 14108 18426 14136 19246
rect 14096 18420 14148 18426
rect 14096 18362 14148 18368
rect 14004 18148 14056 18154
rect 14004 18090 14056 18096
rect 13912 17604 13964 17610
rect 13912 17546 13964 17552
rect 13740 16782 13860 16810
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13740 15978 13768 16594
rect 13832 16250 13860 16782
rect 13910 16688 13966 16697
rect 13910 16623 13966 16632
rect 13924 16590 13952 16623
rect 13912 16584 13964 16590
rect 13912 16526 13964 16532
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13728 15972 13780 15978
rect 13728 15914 13780 15920
rect 13832 15910 13860 16050
rect 13912 15972 13964 15978
rect 13912 15914 13964 15920
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13832 15745 13860 15846
rect 13818 15736 13874 15745
rect 13728 15700 13780 15706
rect 13818 15671 13874 15680
rect 13728 15642 13780 15648
rect 13740 15473 13768 15642
rect 13924 15586 13952 15914
rect 13832 15558 13952 15586
rect 13726 15464 13782 15473
rect 13726 15399 13782 15408
rect 13634 15192 13690 15201
rect 13634 15127 13690 15136
rect 13728 15156 13780 15162
rect 13832 15144 13860 15558
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13780 15116 13860 15144
rect 13728 15098 13780 15104
rect 13556 15014 13860 15042
rect 13452 14952 13504 14958
rect 13358 14920 13414 14929
rect 13452 14894 13504 14900
rect 13358 14855 13414 14864
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13372 14618 13400 14855
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13046 14334 13124 14362
rect 13174 14376 13230 14385
rect 12990 14311 13046 14320
rect 13174 14311 13230 14320
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12808 12844 12860 12850
rect 12728 12804 12808 12832
rect 12808 12786 12860 12792
rect 12714 11792 12770 11801
rect 12714 11727 12770 11736
rect 12728 11354 12756 11727
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12714 10704 12770 10713
rect 12714 10639 12770 10648
rect 12728 9722 12756 10639
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12728 5914 12756 6666
rect 12820 5914 12848 12786
rect 12912 10198 12940 13670
rect 13188 13530 13216 14311
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13174 13152 13230 13161
rect 13174 13087 13230 13096
rect 13188 12753 13216 13087
rect 13280 12986 13308 13262
rect 13358 13152 13414 13161
rect 13358 13087 13414 13096
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13268 12776 13320 12782
rect 13174 12744 13230 12753
rect 13372 12730 13400 13087
rect 13320 12724 13400 12730
rect 13268 12718 13400 12724
rect 13280 12702 13400 12718
rect 13464 12714 13492 14894
rect 13832 14822 13860 15014
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13832 14657 13860 14758
rect 13818 14648 13874 14657
rect 13924 14618 13952 15438
rect 14016 14958 14044 18090
rect 14200 17898 14228 21655
rect 14292 21146 14320 23287
rect 14280 21140 14332 21146
rect 14280 21082 14332 21088
rect 14280 21004 14332 21010
rect 14280 20946 14332 20952
rect 14292 20369 14320 20946
rect 14278 20360 14334 20369
rect 14278 20295 14334 20304
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14292 19786 14320 20198
rect 14280 19780 14332 19786
rect 14280 19722 14332 19728
rect 14384 18714 14412 23967
rect 14476 21418 14504 24006
rect 14464 21412 14516 21418
rect 14464 21354 14516 21360
rect 14568 21146 14596 24550
rect 14844 24410 14872 24754
rect 14922 24712 14978 24721
rect 14922 24647 14924 24656
rect 14976 24647 14978 24656
rect 14924 24618 14976 24624
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 15120 24206 15148 24783
rect 15304 24721 15332 25094
rect 15290 24712 15346 24721
rect 15290 24647 15346 24656
rect 15396 24614 15424 27520
rect 15568 25832 15620 25838
rect 15568 25774 15620 25780
rect 15476 25492 15528 25498
rect 15476 25434 15528 25440
rect 15384 24608 15436 24614
rect 15384 24550 15436 24556
rect 15396 24449 15424 24550
rect 15382 24440 15438 24449
rect 15382 24375 15438 24384
rect 15384 24336 15436 24342
rect 15384 24278 15436 24284
rect 15108 24200 15160 24206
rect 14738 24168 14794 24177
rect 15108 24142 15160 24148
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 14738 24103 14794 24112
rect 14832 24132 14884 24138
rect 14752 23866 14780 24103
rect 14832 24074 14884 24080
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 14844 23322 14872 24074
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15200 23792 15252 23798
rect 15304 23780 15332 24142
rect 15252 23752 15332 23780
rect 15200 23734 15252 23740
rect 15200 23656 15252 23662
rect 15200 23598 15252 23604
rect 14832 23316 14884 23322
rect 14832 23258 14884 23264
rect 14740 23180 14792 23186
rect 14740 23122 14792 23128
rect 14752 22817 14780 23122
rect 14738 22808 14794 22817
rect 14738 22743 14794 22752
rect 14648 22500 14700 22506
rect 14648 22442 14700 22448
rect 14660 21894 14688 22442
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14556 21140 14608 21146
rect 14556 21082 14608 21088
rect 14464 20868 14516 20874
rect 14464 20810 14516 20816
rect 14476 20466 14504 20810
rect 14660 20466 14688 21830
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14752 20330 14780 21286
rect 14844 20913 14872 23258
rect 15212 23118 15240 23598
rect 15396 23594 15424 24278
rect 15384 23588 15436 23594
rect 15384 23530 15436 23536
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15396 22778 15424 23530
rect 15384 22772 15436 22778
rect 15384 22714 15436 22720
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 15304 22098 15332 22374
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15304 21690 15332 22034
rect 15292 21684 15344 21690
rect 15292 21626 15344 21632
rect 15106 21312 15162 21321
rect 15106 21247 15162 21256
rect 15120 21078 15148 21247
rect 15108 21072 15160 21078
rect 15108 21014 15160 21020
rect 15292 21004 15344 21010
rect 15292 20946 15344 20952
rect 14830 20904 14886 20913
rect 14830 20839 14886 20848
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14740 20324 14792 20330
rect 14740 20266 14792 20272
rect 14830 20224 14886 20233
rect 14830 20159 14886 20168
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14568 19378 14596 19654
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14568 19174 14596 19314
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14738 19136 14794 19145
rect 14568 18766 14596 19110
rect 14738 19071 14794 19080
rect 14556 18760 14608 18766
rect 14384 18686 14504 18714
rect 14556 18702 14608 18708
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14384 18193 14412 18566
rect 14370 18184 14426 18193
rect 14370 18119 14426 18128
rect 14200 17870 14320 17898
rect 14188 17808 14240 17814
rect 14186 17776 14188 17785
rect 14240 17776 14242 17785
rect 14186 17711 14242 17720
rect 14292 16250 14320 17870
rect 14372 17128 14424 17134
rect 14370 17096 14372 17105
rect 14424 17096 14426 17105
rect 14370 17031 14426 17040
rect 14280 16244 14332 16250
rect 14280 16186 14332 16192
rect 14370 16144 14426 16153
rect 14370 16079 14426 16088
rect 14278 16008 14334 16017
rect 14278 15943 14334 15952
rect 14292 15706 14320 15943
rect 14384 15910 14412 16079
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 14186 15328 14242 15337
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 13818 14583 13874 14592
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13740 13326 13768 13806
rect 13818 13560 13874 13569
rect 13924 13530 13952 14554
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 14016 13569 14044 13942
rect 14108 13802 14136 15302
rect 14186 15263 14242 15272
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 14002 13560 14058 13569
rect 13818 13495 13874 13504
rect 13912 13524 13964 13530
rect 13832 13462 13860 13495
rect 14200 13530 14228 15263
rect 14278 15192 14334 15201
rect 14476 15162 14504 18686
rect 14554 17504 14610 17513
rect 14554 17439 14610 17448
rect 14568 16794 14596 17439
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14278 15127 14334 15136
rect 14464 15156 14516 15162
rect 14292 14618 14320 15127
rect 14464 15098 14516 15104
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14384 14249 14412 14554
rect 14568 14550 14596 16186
rect 14660 15706 14688 16526
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 14646 15464 14702 15473
rect 14646 15399 14702 15408
rect 14660 15094 14688 15399
rect 14648 15088 14700 15094
rect 14648 15030 14700 15036
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 14370 14240 14426 14249
rect 14370 14175 14426 14184
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14476 13841 14504 13874
rect 14462 13832 14518 13841
rect 14462 13767 14518 13776
rect 14370 13696 14426 13705
rect 14370 13631 14426 13640
rect 14002 13495 14058 13504
rect 14188 13524 14240 13530
rect 13912 13466 13964 13472
rect 14188 13466 14240 13472
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13924 13190 13952 13466
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13542 13016 13598 13025
rect 13542 12951 13598 12960
rect 13174 12679 13230 12688
rect 13372 12646 13400 12702
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13188 11626 13216 12038
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 13082 11520 13138 11529
rect 13082 11455 13138 11464
rect 12990 11248 13046 11257
rect 12990 11183 13046 11192
rect 13004 11150 13032 11183
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13004 10810 13032 11086
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 13004 10010 13032 10066
rect 12912 9982 13032 10010
rect 12912 9897 12940 9982
rect 12898 9888 12954 9897
rect 12898 9823 12954 9832
rect 12912 9654 12940 9823
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12898 8528 12954 8537
rect 13004 8498 13032 9318
rect 12898 8463 12954 8472
rect 12992 8492 13044 8498
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12806 5672 12862 5681
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12728 5030 12756 5646
rect 12912 5658 12940 8463
rect 12992 8434 13044 8440
rect 13004 7750 13032 8434
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 13004 7206 13032 7686
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 13004 6254 13032 7142
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 13004 5681 13032 5714
rect 12862 5630 12940 5658
rect 12990 5672 13046 5681
rect 12806 5607 12862 5616
rect 12990 5607 13046 5616
rect 13096 5216 13124 11455
rect 13188 10062 13216 11562
rect 13450 11384 13506 11393
rect 13268 11348 13320 11354
rect 13320 11308 13400 11336
rect 13556 11354 13584 12951
rect 13924 12850 13952 13126
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13910 12200 13966 12209
rect 13910 12135 13966 12144
rect 13924 11898 13952 12135
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13450 11319 13506 11328
rect 13544 11348 13596 11354
rect 13268 11290 13320 11296
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13188 9081 13216 9114
rect 13372 9110 13400 11308
rect 13464 10266 13492 11319
rect 13544 11290 13596 11296
rect 13556 10810 13584 11290
rect 13634 11248 13690 11257
rect 13634 11183 13690 11192
rect 13648 10985 13676 11183
rect 13634 10976 13690 10985
rect 13634 10911 13690 10920
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13542 10704 13598 10713
rect 13832 10674 13860 11494
rect 13542 10639 13598 10648
rect 13820 10668 13872 10674
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13360 9104 13412 9110
rect 13174 9072 13230 9081
rect 13360 9046 13412 9052
rect 13174 9007 13230 9016
rect 13464 8838 13492 9318
rect 13556 8906 13584 10639
rect 13820 10610 13872 10616
rect 13818 10432 13874 10441
rect 13818 10367 13874 10376
rect 13832 10266 13860 10367
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13740 9178 13768 10134
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13726 9072 13782 9081
rect 13726 9007 13782 9016
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13464 7750 13492 8774
rect 13740 8537 13768 9007
rect 13726 8528 13782 8537
rect 13726 8463 13782 8472
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13174 7168 13230 7177
rect 13174 7103 13230 7112
rect 12912 5188 13124 5216
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12452 4146 12480 4626
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12348 4140 12400 4146
rect 12440 4140 12492 4146
rect 12400 4100 12440 4128
rect 12348 4082 12400 4088
rect 12440 4082 12492 4088
rect 12544 4049 12572 4558
rect 12530 4040 12586 4049
rect 12530 3975 12586 3984
rect 12544 3942 12572 3975
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12176 3692 12296 3720
rect 12070 3360 12126 3369
rect 12070 3295 12126 3304
rect 12176 3126 12204 3692
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12268 3369 12296 3538
rect 12254 3360 12310 3369
rect 12254 3295 12310 3304
rect 12268 3194 12296 3295
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 11978 2136 12034 2145
rect 11978 2071 12034 2080
rect 11886 776 11942 785
rect 11886 711 11942 720
rect 12268 480 12296 2994
rect 12912 2666 12940 5188
rect 13082 5128 13138 5137
rect 13082 5063 13138 5072
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 12820 2638 12940 2666
rect 12820 480 12848 2638
rect 13004 2514 13032 4966
rect 13096 3738 13124 5063
rect 13188 4758 13216 7103
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13280 6458 13308 6870
rect 13360 6792 13412 6798
rect 13358 6760 13360 6769
rect 13412 6760 13414 6769
rect 13358 6695 13414 6704
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13280 5545 13308 6394
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13266 5536 13322 5545
rect 13266 5471 13322 5480
rect 13176 4752 13228 4758
rect 13176 4694 13228 4700
rect 13188 4146 13216 4694
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 13280 1873 13308 2790
rect 13266 1864 13322 1873
rect 13266 1799 13322 1808
rect 13372 480 13400 5850
rect 13464 5234 13492 7686
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13556 7206 13584 7346
rect 13648 7313 13676 8298
rect 13832 8265 13860 10066
rect 14002 9480 14058 9489
rect 14002 9415 14058 9424
rect 14016 9178 14044 9415
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14108 8945 14136 13330
rect 14384 12986 14412 13631
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14384 12782 14412 12922
rect 14372 12776 14424 12782
rect 14568 12730 14596 14486
rect 14752 13394 14780 19071
rect 14844 17082 14872 20159
rect 15304 20074 15332 20946
rect 15382 20632 15438 20641
rect 15382 20567 15438 20576
rect 15396 20233 15424 20567
rect 15382 20224 15438 20233
rect 15382 20159 15438 20168
rect 15120 20058 15332 20074
rect 15108 20052 15332 20058
rect 15160 20046 15332 20052
rect 15108 19994 15160 20000
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15108 19440 15160 19446
rect 15304 19394 15332 20046
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15160 19388 15332 19394
rect 15108 19382 15332 19388
rect 15120 19366 15332 19382
rect 15396 18986 15424 19654
rect 15120 18970 15424 18986
rect 15488 18970 15516 25434
rect 15580 23322 15608 25774
rect 15936 25356 15988 25362
rect 15936 25298 15988 25304
rect 15660 24880 15712 24886
rect 15660 24822 15712 24828
rect 15752 24880 15804 24886
rect 15752 24822 15804 24828
rect 15568 23316 15620 23322
rect 15568 23258 15620 23264
rect 15566 22536 15622 22545
rect 15566 22471 15622 22480
rect 15580 19310 15608 22471
rect 15672 20058 15700 24822
rect 15764 24410 15792 24822
rect 15948 24614 15976 25298
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 15752 24404 15804 24410
rect 15752 24346 15804 24352
rect 15764 23848 15792 24346
rect 15844 23860 15896 23866
rect 15764 23820 15844 23848
rect 15844 23802 15896 23808
rect 15948 22098 15976 24550
rect 16040 22114 16068 27520
rect 16304 24676 16356 24682
rect 16304 24618 16356 24624
rect 16118 23624 16174 23633
rect 16118 23559 16174 23568
rect 16132 22234 16160 23559
rect 16212 23180 16264 23186
rect 16212 23122 16264 23128
rect 16224 22778 16252 23122
rect 16212 22772 16264 22778
rect 16212 22714 16264 22720
rect 16316 22574 16344 24618
rect 16396 24608 16448 24614
rect 16396 24550 16448 24556
rect 16488 24608 16540 24614
rect 16488 24550 16540 24556
rect 16304 22568 16356 22574
rect 16304 22510 16356 22516
rect 16120 22228 16172 22234
rect 16120 22170 16172 22176
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 15844 22092 15896 22098
rect 15844 22034 15896 22040
rect 15936 22092 15988 22098
rect 16040 22086 16160 22114
rect 15936 22034 15988 22040
rect 15856 21350 15884 22034
rect 15934 21992 15990 22001
rect 15934 21927 15990 21936
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15764 20602 15792 21082
rect 15856 20942 15884 21286
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 15752 20596 15804 20602
rect 15752 20538 15804 20544
rect 15842 20088 15898 20097
rect 15660 20052 15712 20058
rect 15842 20023 15898 20032
rect 15660 19994 15712 20000
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15672 18970 15700 19994
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 15764 19378 15792 19790
rect 15856 19689 15884 20023
rect 15842 19680 15898 19689
rect 15842 19615 15898 19624
rect 15842 19408 15898 19417
rect 15752 19372 15804 19378
rect 15842 19343 15898 19352
rect 15752 19314 15804 19320
rect 15856 19242 15884 19343
rect 15844 19236 15896 19242
rect 15844 19178 15896 19184
rect 15108 18964 15424 18970
rect 15160 18958 15424 18964
rect 15476 18964 15528 18970
rect 15108 18906 15160 18912
rect 15476 18906 15528 18912
rect 15660 18964 15712 18970
rect 15660 18906 15712 18912
rect 15856 18902 15884 19178
rect 15844 18896 15896 18902
rect 15844 18838 15896 18844
rect 15384 18828 15436 18834
rect 15384 18770 15436 18776
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 15028 17678 15056 18226
rect 15106 18184 15162 18193
rect 15106 18119 15162 18128
rect 15120 17882 15148 18119
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15304 17338 15332 17750
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 14844 17054 15056 17082
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 14936 16833 14964 16934
rect 14922 16824 14978 16833
rect 14922 16759 14978 16768
rect 14832 16720 14884 16726
rect 14830 16688 14832 16697
rect 14884 16688 14886 16697
rect 14830 16623 14886 16632
rect 15028 16436 15056 17054
rect 15106 16688 15162 16697
rect 15106 16623 15108 16632
rect 15160 16623 15162 16632
rect 15108 16594 15160 16600
rect 14844 16408 15056 16436
rect 14844 15688 14872 16408
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14922 16008 14978 16017
rect 14922 15943 14924 15952
rect 14976 15943 14978 15952
rect 14924 15914 14976 15920
rect 14844 15660 14964 15688
rect 14936 15473 14964 15660
rect 15108 15496 15160 15502
rect 14922 15464 14978 15473
rect 14922 15399 14978 15408
rect 15106 15464 15108 15473
rect 15160 15464 15162 15473
rect 15106 15399 15162 15408
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14922 15056 14978 15065
rect 14922 14991 14978 15000
rect 14936 14958 14964 14991
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 15108 14612 15160 14618
rect 15396 14600 15424 18770
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15658 18592 15714 18601
rect 15658 18527 15714 18536
rect 15672 18222 15700 18527
rect 15856 18426 15884 18702
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15672 17338 15700 17478
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15580 15910 15608 16526
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15580 15570 15608 15846
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15568 15360 15620 15366
rect 15672 15337 15700 16390
rect 15568 15302 15620 15308
rect 15658 15328 15714 15337
rect 15488 15026 15516 15302
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15160 14572 15424 14600
rect 15108 14554 15160 14560
rect 15488 14482 15516 14962
rect 15476 14476 15528 14482
rect 15396 14436 15476 14464
rect 15292 14408 15344 14414
rect 15290 14376 15292 14385
rect 15344 14376 15346 14385
rect 15290 14311 15346 14320
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 15304 13326 15332 13942
rect 14924 13320 14976 13326
rect 14922 13288 14924 13297
rect 15292 13320 15344 13326
rect 14976 13288 14978 13297
rect 15292 13262 15344 13268
rect 14922 13223 14978 13232
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14660 12850 14688 13126
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14372 12718 14424 12724
rect 14476 12702 14596 12730
rect 14476 12628 14504 12702
rect 14384 12600 14504 12628
rect 14556 12640 14608 12646
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11665 14228 12038
rect 14186 11656 14242 11665
rect 14186 11591 14242 11600
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14200 11014 14228 11494
rect 14278 11384 14334 11393
rect 14278 11319 14280 11328
rect 14332 11319 14334 11328
rect 14280 11290 14332 11296
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14200 10538 14228 10950
rect 14188 10532 14240 10538
rect 14188 10474 14240 10480
rect 14200 10169 14228 10474
rect 14186 10160 14242 10169
rect 14186 10095 14242 10104
rect 14200 9994 14228 10095
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 14188 9716 14240 9722
rect 14240 9676 14320 9704
rect 14188 9658 14240 9664
rect 14292 9568 14320 9676
rect 14200 9540 14320 9568
rect 14200 9058 14228 9540
rect 14384 9500 14412 12600
rect 14556 12582 14608 12588
rect 14568 12481 14596 12582
rect 14554 12472 14610 12481
rect 14554 12407 14610 12416
rect 14554 12336 14610 12345
rect 14554 12271 14610 12280
rect 14462 10840 14518 10849
rect 14462 10775 14518 10784
rect 14476 10441 14504 10775
rect 14462 10432 14518 10441
rect 14462 10367 14518 10376
rect 14292 9472 14412 9500
rect 14292 9353 14320 9472
rect 14278 9344 14334 9353
rect 14278 9279 14334 9288
rect 14200 9030 14412 9058
rect 14188 8968 14240 8974
rect 14094 8936 14150 8945
rect 14188 8910 14240 8916
rect 14094 8871 14150 8880
rect 13818 8256 13874 8265
rect 13818 8191 13874 8200
rect 14002 7576 14058 7585
rect 14002 7511 14058 7520
rect 14016 7410 14044 7511
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 13820 7336 13872 7342
rect 13634 7304 13690 7313
rect 13634 7239 13690 7248
rect 13740 7296 13820 7324
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13556 6798 13584 7142
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13740 6662 13768 7296
rect 13820 7278 13872 7284
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13726 5808 13782 5817
rect 13924 5760 13952 7142
rect 14016 7002 14044 7346
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 14108 6440 14136 8871
rect 14200 8090 14228 8910
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14280 7200 14332 7206
rect 14186 7168 14242 7177
rect 14280 7142 14332 7148
rect 14186 7103 14242 7112
rect 13782 5752 13952 5760
rect 13726 5743 13952 5752
rect 13740 5732 13952 5743
rect 14016 6412 14136 6440
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13740 5166 13768 5732
rect 13910 5672 13966 5681
rect 13820 5636 13872 5642
rect 13910 5607 13966 5616
rect 13820 5578 13872 5584
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13832 4826 13860 5578
rect 13924 5370 13952 5607
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 14016 5250 14044 6412
rect 14094 6352 14150 6361
rect 14094 6287 14150 6296
rect 14108 6254 14136 6287
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14108 5914 14136 6190
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 13924 5222 14044 5250
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13740 4298 13768 4626
rect 13464 4270 13768 4298
rect 13464 4146 13492 4270
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13556 2689 13584 4150
rect 13740 3738 13768 4270
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13636 2848 13688 2854
rect 13634 2816 13636 2825
rect 13688 2816 13690 2825
rect 13634 2751 13690 2760
rect 13542 2680 13598 2689
rect 13542 2615 13598 2624
rect 13740 2582 13768 2994
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 13740 1873 13768 2518
rect 13726 1864 13782 1873
rect 13726 1799 13782 1808
rect 13924 480 13952 5222
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14016 2961 14044 4966
rect 14096 4616 14148 4622
rect 14094 4584 14096 4593
rect 14148 4584 14150 4593
rect 14094 4519 14150 4528
rect 14108 4214 14136 4519
rect 14096 4208 14148 4214
rect 14096 4150 14148 4156
rect 14200 3738 14228 7103
rect 14292 7041 14320 7142
rect 14278 7032 14334 7041
rect 14278 6967 14334 6976
rect 14292 5914 14320 6967
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14292 4457 14320 5102
rect 14384 4826 14412 9030
rect 14476 8634 14504 10367
rect 14568 9654 14596 12271
rect 14660 11694 14688 12786
rect 14924 12708 14976 12714
rect 14924 12650 14976 12656
rect 14936 12442 14964 12650
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 15200 12436 15252 12442
rect 15304 12424 15332 13262
rect 15252 12396 15332 12424
rect 15200 12378 15252 12384
rect 15396 12356 15424 14436
rect 15476 14418 15528 14424
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15304 12328 15424 12356
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15304 11898 15332 12328
rect 15382 12200 15438 12209
rect 15382 12135 15438 12144
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14830 11384 14886 11393
rect 14830 11319 14886 11328
rect 15290 11384 15346 11393
rect 15290 11319 15346 11328
rect 14740 11144 14792 11150
rect 14738 11112 14740 11121
rect 14792 11112 14794 11121
rect 14738 11047 14794 11056
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14660 8022 14688 9318
rect 14752 8974 14780 10406
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14648 8016 14700 8022
rect 14648 7958 14700 7964
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14476 7342 14504 7686
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14554 7304 14610 7313
rect 14554 7239 14610 7248
rect 14568 6390 14596 7239
rect 14660 6866 14688 7958
rect 14752 7041 14780 8774
rect 14738 7032 14794 7041
rect 14738 6967 14794 6976
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14740 6724 14792 6730
rect 14740 6666 14792 6672
rect 14752 6497 14780 6666
rect 14738 6488 14794 6497
rect 14738 6423 14794 6432
rect 14556 6384 14608 6390
rect 14556 6326 14608 6332
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14278 4448 14334 4457
rect 14278 4383 14334 4392
rect 14384 4078 14412 4762
rect 14568 4593 14596 4966
rect 14554 4584 14610 4593
rect 14554 4519 14610 4528
rect 14740 4480 14792 4486
rect 14554 4448 14610 4457
rect 14740 4422 14792 4428
rect 14554 4383 14610 4392
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14292 3641 14320 3878
rect 14278 3632 14334 3641
rect 14568 3618 14596 4383
rect 14646 4176 14702 4185
rect 14646 4111 14702 4120
rect 14660 4078 14688 4111
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14660 3738 14688 4014
rect 14752 4010 14780 4422
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14568 3590 14688 3618
rect 14278 3567 14334 3576
rect 14370 3496 14426 3505
rect 14370 3431 14426 3440
rect 14464 3460 14516 3466
rect 14002 2952 14058 2961
rect 14002 2887 14004 2896
rect 14056 2887 14058 2896
rect 14004 2858 14056 2864
rect 14384 480 14412 3431
rect 14464 3402 14516 3408
rect 14476 3233 14504 3402
rect 14554 3360 14610 3369
rect 14554 3295 14610 3304
rect 14462 3224 14518 3233
rect 14462 3159 14518 3168
rect 14568 3097 14596 3295
rect 14554 3088 14610 3097
rect 14554 3023 14610 3032
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14476 2514 14504 2790
rect 14568 2650 14596 3023
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14554 2408 14610 2417
rect 14554 2343 14610 2352
rect 14568 2310 14596 2343
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 14660 1902 14688 3590
rect 14648 1896 14700 1902
rect 14648 1838 14700 1844
rect 14844 1034 14872 11319
rect 15304 11218 15332 11319
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10305 15332 11154
rect 15290 10296 15346 10305
rect 15396 10266 15424 12135
rect 15488 12073 15516 13806
rect 15580 12714 15608 15302
rect 15658 15263 15714 15272
rect 15764 15178 15792 17818
rect 15842 17368 15898 17377
rect 15842 17303 15898 17312
rect 15672 15150 15792 15178
rect 15568 12708 15620 12714
rect 15568 12650 15620 12656
rect 15568 12096 15620 12102
rect 15474 12064 15530 12073
rect 15568 12038 15620 12044
rect 15474 11999 15530 12008
rect 15488 11529 15516 11999
rect 15580 11626 15608 12038
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15474 11520 15530 11529
rect 15474 11455 15530 11464
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15290 10231 15346 10240
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 14922 9344 14978 9353
rect 14922 9279 14978 9288
rect 14936 9178 14964 9279
rect 15120 9178 15148 9522
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15292 9104 15344 9110
rect 15292 9046 15344 9052
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15304 8616 15332 9046
rect 15120 8588 15332 8616
rect 15120 8090 15148 8588
rect 15488 8362 15516 11154
rect 15580 10674 15608 11562
rect 15672 11354 15700 15150
rect 15752 14884 15804 14890
rect 15752 14826 15804 14832
rect 15764 14618 15792 14826
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15764 13190 15792 14554
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15764 12442 15792 13126
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15658 10976 15714 10985
rect 15658 10911 15714 10920
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15580 10470 15608 10610
rect 15568 10464 15620 10470
rect 15672 10441 15700 10911
rect 15750 10704 15806 10713
rect 15750 10639 15806 10648
rect 15568 10406 15620 10412
rect 15658 10432 15714 10441
rect 15658 10367 15714 10376
rect 15658 10296 15714 10305
rect 15764 10266 15792 10639
rect 15658 10231 15714 10240
rect 15752 10260 15804 10266
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15476 8356 15528 8362
rect 15476 8298 15528 8304
rect 15580 8294 15608 8774
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15304 7886 15332 8230
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15304 6798 15332 7822
rect 15672 7342 15700 10231
rect 15752 10202 15804 10208
rect 15752 9444 15804 9450
rect 15752 9386 15804 9392
rect 15764 9081 15792 9386
rect 15856 9110 15884 17303
rect 15948 15348 15976 21927
rect 16026 21720 16082 21729
rect 16026 21655 16082 21664
rect 16040 21185 16068 21655
rect 16026 21176 16082 21185
rect 16026 21111 16082 21120
rect 16040 16776 16068 21111
rect 16132 17921 16160 22086
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 16224 19553 16252 20198
rect 16210 19544 16266 19553
rect 16210 19479 16266 19488
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 16224 18737 16252 19110
rect 16210 18728 16266 18737
rect 16210 18663 16266 18672
rect 16118 17912 16174 17921
rect 16118 17847 16174 17856
rect 16040 16748 16252 16776
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 16040 15473 16068 16594
rect 16026 15464 16082 15473
rect 16026 15399 16082 15408
rect 15948 15320 16068 15348
rect 15936 14544 15988 14550
rect 15936 14486 15988 14492
rect 15948 13734 15976 14486
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15936 13184 15988 13190
rect 15934 13152 15936 13161
rect 15988 13152 15990 13161
rect 15934 13087 15990 13096
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 15948 10062 15976 11222
rect 16040 10849 16068 15320
rect 16224 13512 16252 16748
rect 16316 16182 16344 22170
rect 16408 21486 16436 24550
rect 16500 24410 16528 24550
rect 16488 24404 16540 24410
rect 16488 24346 16540 24352
rect 16500 23526 16528 24346
rect 16488 23520 16540 23526
rect 16488 23462 16540 23468
rect 16592 23225 16620 27520
rect 17038 26344 17094 26353
rect 17038 26279 17094 26288
rect 16948 25968 17000 25974
rect 16684 25916 16948 25922
rect 16684 25910 17000 25916
rect 16684 25894 16988 25910
rect 16684 25702 16712 25894
rect 16672 25696 16724 25702
rect 16672 25638 16724 25644
rect 17052 25514 17080 26279
rect 16868 25486 17080 25514
rect 16868 25362 16896 25486
rect 16856 25356 16908 25362
rect 16856 25298 16908 25304
rect 16948 25356 17000 25362
rect 16948 25298 17000 25304
rect 16672 25152 16724 25158
rect 16672 25094 16724 25100
rect 16684 24274 16712 25094
rect 16672 24268 16724 24274
rect 16672 24210 16724 24216
rect 16960 24206 16988 25298
rect 16948 24200 17000 24206
rect 16946 24168 16948 24177
rect 17000 24168 17002 24177
rect 16672 24132 16724 24138
rect 16946 24103 17002 24112
rect 16672 24074 16724 24080
rect 16578 23216 16634 23225
rect 16578 23151 16634 23160
rect 16488 23112 16540 23118
rect 16488 23054 16540 23060
rect 16500 22506 16528 23054
rect 16488 22500 16540 22506
rect 16488 22442 16540 22448
rect 16500 22166 16528 22442
rect 16488 22160 16540 22166
rect 16488 22102 16540 22108
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16396 21480 16448 21486
rect 16396 21422 16448 21428
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 16408 21185 16436 21286
rect 16394 21176 16450 21185
rect 16394 21111 16450 21120
rect 16500 20641 16528 21898
rect 16684 21418 16712 24074
rect 17052 24018 17080 25486
rect 17144 24585 17172 27520
rect 17222 25664 17278 25673
rect 17222 25599 17278 25608
rect 17236 25265 17264 25599
rect 17500 25356 17552 25362
rect 17500 25298 17552 25304
rect 17316 25288 17368 25294
rect 17222 25256 17278 25265
rect 17316 25230 17368 25236
rect 17222 25191 17278 25200
rect 17328 25158 17356 25230
rect 17316 25152 17368 25158
rect 17316 25094 17368 25100
rect 17328 24818 17356 25094
rect 17316 24812 17368 24818
rect 17316 24754 17368 24760
rect 17408 24812 17460 24818
rect 17408 24754 17460 24760
rect 17130 24576 17186 24585
rect 17130 24511 17186 24520
rect 17052 23990 17172 24018
rect 17038 23896 17094 23905
rect 16764 23860 16816 23866
rect 17038 23831 17094 23840
rect 16764 23802 16816 23808
rect 16776 23254 16804 23802
rect 16764 23248 16816 23254
rect 16764 23190 16816 23196
rect 16776 22234 16804 23190
rect 17052 22710 17080 23831
rect 17040 22704 17092 22710
rect 17040 22646 17092 22652
rect 17144 22386 17172 23990
rect 17328 23866 17356 24754
rect 17420 24206 17448 24754
rect 17512 24614 17540 25298
rect 17592 24676 17644 24682
rect 17592 24618 17644 24624
rect 17500 24608 17552 24614
rect 17500 24550 17552 24556
rect 17408 24200 17460 24206
rect 17408 24142 17460 24148
rect 17316 23860 17368 23866
rect 17316 23802 17368 23808
rect 17222 23080 17278 23089
rect 17222 23015 17278 23024
rect 17236 22409 17264 23015
rect 16868 22358 17172 22386
rect 17222 22400 17278 22409
rect 16764 22228 16816 22234
rect 16764 22170 16816 22176
rect 16764 21684 16816 21690
rect 16764 21626 16816 21632
rect 16672 21412 16724 21418
rect 16672 21354 16724 21360
rect 16486 20632 16542 20641
rect 16486 20567 16542 20576
rect 16396 20528 16448 20534
rect 16394 20496 16396 20505
rect 16448 20496 16450 20505
rect 16394 20431 16450 20440
rect 16394 20360 16450 20369
rect 16394 20295 16450 20304
rect 16488 20324 16540 20330
rect 16408 17882 16436 20295
rect 16488 20266 16540 20272
rect 16500 20058 16528 20266
rect 16488 20052 16540 20058
rect 16488 19994 16540 20000
rect 16488 19916 16540 19922
rect 16488 19858 16540 19864
rect 16500 19174 16528 19858
rect 16578 19544 16634 19553
rect 16578 19479 16580 19488
rect 16632 19479 16634 19488
rect 16580 19450 16632 19456
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16488 18080 16540 18086
rect 16486 18048 16488 18057
rect 16540 18048 16542 18057
rect 16486 17983 16542 17992
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 16500 17814 16528 17983
rect 16488 17808 16540 17814
rect 16488 17750 16540 17756
rect 16776 17762 16804 21626
rect 16868 20058 16896 22358
rect 17222 22335 17278 22344
rect 16948 22228 17000 22234
rect 16948 22170 17000 22176
rect 16960 22098 16988 22170
rect 17038 22128 17094 22137
rect 16948 22092 17000 22098
rect 17038 22063 17094 22072
rect 16948 22034 17000 22040
rect 16960 21078 16988 22034
rect 17052 21690 17080 22063
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 17040 21344 17092 21350
rect 17038 21312 17040 21321
rect 17092 21312 17094 21321
rect 17038 21247 17094 21256
rect 16948 21072 17000 21078
rect 16948 21014 17000 21020
rect 16960 20466 16988 21014
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16960 19938 16988 20402
rect 17038 20088 17094 20097
rect 17038 20023 17094 20032
rect 16868 19922 16988 19938
rect 16868 19916 17000 19922
rect 16868 19910 16948 19916
rect 16868 19514 16896 19910
rect 16948 19858 17000 19864
rect 16960 19827 16988 19858
rect 17052 19786 17080 20023
rect 17144 19990 17172 21966
rect 17132 19984 17184 19990
rect 17132 19926 17184 19932
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 16948 19712 17000 19718
rect 16948 19654 17000 19660
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16960 19310 16988 19654
rect 16948 19304 17000 19310
rect 16946 19272 16948 19281
rect 17000 19272 17002 19281
rect 16946 19207 17002 19216
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17144 18737 17172 19110
rect 17130 18728 17186 18737
rect 17130 18663 17186 18672
rect 16776 17734 16988 17762
rect 16764 17604 16816 17610
rect 16764 17546 16816 17552
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16684 17377 16712 17478
rect 16670 17368 16726 17377
rect 16670 17303 16726 17312
rect 16486 17232 16542 17241
rect 16486 17167 16488 17176
rect 16540 17167 16542 17176
rect 16488 17138 16540 17144
rect 16776 17134 16804 17546
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16580 17060 16632 17066
rect 16580 17002 16632 17008
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16408 16794 16436 16934
rect 16396 16788 16448 16794
rect 16396 16730 16448 16736
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16408 16250 16436 16526
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 16316 15978 16344 16118
rect 16304 15972 16356 15978
rect 16304 15914 16356 15920
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16408 14550 16436 15506
rect 16592 14618 16620 17002
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16868 16658 16896 16934
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16776 16114 16804 16390
rect 16764 16108 16816 16114
rect 16764 16050 16816 16056
rect 16672 15972 16724 15978
rect 16672 15914 16724 15920
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16500 14074 16528 14418
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16580 13524 16632 13530
rect 16224 13484 16436 13512
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16118 13016 16174 13025
rect 16118 12951 16120 12960
rect 16172 12951 16174 12960
rect 16120 12922 16172 12928
rect 16316 12918 16344 13330
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16210 12744 16266 12753
rect 16210 12679 16266 12688
rect 16224 12646 16252 12679
rect 16316 12646 16344 12854
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16118 12336 16174 12345
rect 16118 12271 16174 12280
rect 16026 10840 16082 10849
rect 16026 10775 16082 10784
rect 16040 10305 16068 10775
rect 16026 10296 16082 10305
rect 16026 10231 16082 10240
rect 16026 10160 16082 10169
rect 16026 10095 16082 10104
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15948 9586 15976 9998
rect 16040 9654 16068 10095
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15844 9104 15896 9110
rect 15750 9072 15806 9081
rect 15844 9046 15896 9052
rect 15750 9007 15806 9016
rect 15750 8664 15806 8673
rect 15750 8599 15752 8608
rect 15804 8599 15806 8608
rect 15752 8570 15804 8576
rect 16040 8566 16068 9590
rect 16132 9382 16160 12271
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16224 11801 16252 12038
rect 16408 11937 16436 13484
rect 16580 13466 16632 13472
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16394 11928 16450 11937
rect 16394 11863 16450 11872
rect 16210 11792 16266 11801
rect 16408 11744 16436 11863
rect 16210 11727 16266 11736
rect 16316 11716 16436 11744
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16224 11150 16252 11630
rect 16316 11218 16344 11716
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16212 10600 16264 10606
rect 16210 10568 16212 10577
rect 16264 10568 16266 10577
rect 16210 10503 16266 10512
rect 16304 10464 16356 10470
rect 16210 10432 16266 10441
rect 16304 10406 16356 10412
rect 16210 10367 16266 10376
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16224 8616 16252 10367
rect 16316 9382 16344 10406
rect 16408 10266 16436 11086
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16394 10024 16450 10033
rect 16394 9959 16450 9968
rect 16408 9518 16436 9959
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 9081 16344 9318
rect 16302 9072 16358 9081
rect 16302 9007 16358 9016
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16132 8588 16252 8616
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15752 7268 15804 7274
rect 15752 7210 15804 7216
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15488 6118 15516 6802
rect 15580 6458 15608 7142
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15476 6112 15528 6118
rect 15474 6080 15476 6089
rect 15528 6080 15530 6089
rect 15474 6015 15530 6024
rect 15290 5944 15346 5953
rect 15580 5914 15608 6394
rect 15290 5879 15292 5888
rect 15344 5879 15346 5888
rect 15568 5908 15620 5914
rect 15292 5850 15344 5856
rect 15568 5850 15620 5856
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15304 5370 15332 5646
rect 15384 5636 15436 5642
rect 15384 5578 15436 5584
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15396 5166 15424 5578
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15108 5092 15160 5098
rect 15108 5034 15160 5040
rect 15120 4826 15148 5034
rect 15384 5024 15436 5030
rect 15488 4978 15516 5714
rect 15436 4972 15516 4978
rect 15384 4966 15516 4972
rect 15396 4950 15516 4966
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 15290 4720 15346 4729
rect 15290 4655 15346 4664
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15016 4208 15068 4214
rect 15014 4176 15016 4185
rect 15068 4176 15070 4185
rect 14924 4140 14976 4146
rect 15304 4146 15332 4655
rect 15396 4214 15424 4950
rect 15672 4729 15700 6598
rect 15658 4720 15714 4729
rect 15658 4655 15714 4664
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15384 4208 15436 4214
rect 15384 4150 15436 4156
rect 15014 4111 15070 4120
rect 15292 4140 15344 4146
rect 14924 4082 14976 4088
rect 15292 4082 15344 4088
rect 14936 3534 14964 4082
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 14936 2650 14964 2926
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 15304 2514 15332 3878
rect 15396 3777 15424 4150
rect 15672 3942 15700 4558
rect 15764 4049 15792 7210
rect 15750 4040 15806 4049
rect 15750 3975 15806 3984
rect 15660 3936 15712 3942
rect 15856 3924 15884 8366
rect 16132 8106 16160 8588
rect 16210 8528 16266 8537
rect 16210 8463 16212 8472
rect 16264 8463 16266 8472
rect 16212 8434 16264 8440
rect 15948 8078 16160 8106
rect 15948 6458 15976 8078
rect 16120 8016 16172 8022
rect 16120 7958 16172 7964
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 16040 5710 16068 7686
rect 16132 7410 16160 7958
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16132 6662 16160 6734
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16132 5778 16160 6598
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 16132 5302 16160 5714
rect 16120 5296 16172 5302
rect 16120 5238 16172 5244
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16040 4486 16068 5170
rect 16132 4622 16160 5238
rect 16120 4616 16172 4622
rect 16120 4558 16172 4564
rect 16028 4480 16080 4486
rect 16028 4422 16080 4428
rect 16316 4298 16344 8910
rect 16500 6984 16528 12922
rect 16592 12782 16620 13466
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16578 12336 16634 12345
rect 16684 12322 16712 15914
rect 16960 15858 16988 17734
rect 17236 16810 17264 22335
rect 17314 22128 17370 22137
rect 17314 22063 17370 22072
rect 17328 20262 17356 22063
rect 17420 21146 17448 24142
rect 17512 23769 17540 24550
rect 17498 23760 17554 23769
rect 17498 23695 17554 23704
rect 17604 23066 17632 24618
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 17696 23225 17724 24210
rect 17788 23361 17816 27520
rect 18340 25974 18368 27520
rect 18512 26716 18564 26722
rect 18512 26658 18564 26664
rect 18420 26036 18472 26042
rect 18420 25978 18472 25984
rect 18236 25968 18288 25974
rect 18236 25910 18288 25916
rect 18328 25968 18380 25974
rect 18328 25910 18380 25916
rect 18248 25242 18276 25910
rect 18248 25214 18368 25242
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 18236 25152 18288 25158
rect 18236 25094 18288 25100
rect 18156 24750 18184 25094
rect 18248 24818 18276 25094
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 18144 24744 18196 24750
rect 18144 24686 18196 24692
rect 17960 24608 18012 24614
rect 17960 24550 18012 24556
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 17880 23526 17908 24142
rect 17868 23520 17920 23526
rect 17868 23462 17920 23468
rect 17774 23352 17830 23361
rect 17774 23287 17830 23296
rect 17682 23216 17738 23225
rect 17682 23151 17738 23160
rect 17604 23038 17724 23066
rect 17880 23050 17908 23462
rect 17498 22944 17554 22953
rect 17498 22879 17554 22888
rect 17512 22098 17540 22879
rect 17592 22704 17644 22710
rect 17592 22646 17644 22652
rect 17500 22092 17552 22098
rect 17500 22034 17552 22040
rect 17500 21956 17552 21962
rect 17500 21898 17552 21904
rect 17408 21140 17460 21146
rect 17408 21082 17460 21088
rect 17316 20256 17368 20262
rect 17316 20198 17368 20204
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17420 19514 17448 19994
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17512 18850 17540 21898
rect 17604 21554 17632 22646
rect 17696 21962 17724 23038
rect 17868 23044 17920 23050
rect 17868 22986 17920 22992
rect 17880 22710 17908 22986
rect 17868 22704 17920 22710
rect 17868 22646 17920 22652
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 17776 22228 17828 22234
rect 17776 22170 17828 22176
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 17682 21856 17738 21865
rect 17682 21791 17738 21800
rect 17592 21548 17644 21554
rect 17592 21490 17644 21496
rect 17696 20913 17724 21791
rect 17682 20904 17738 20913
rect 17788 20874 17816 22170
rect 17880 22098 17908 22510
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17972 21434 18000 24550
rect 18052 24064 18104 24070
rect 18052 24006 18104 24012
rect 18064 22642 18092 24006
rect 18144 23656 18196 23662
rect 18144 23598 18196 23604
rect 18052 22636 18104 22642
rect 18052 22578 18104 22584
rect 18156 22506 18184 23598
rect 18234 23488 18290 23497
rect 18234 23423 18290 23432
rect 18144 22500 18196 22506
rect 18144 22442 18196 22448
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 18064 21690 18092 22374
rect 18052 21684 18104 21690
rect 18052 21626 18104 21632
rect 18156 21554 18184 22442
rect 18248 22438 18276 23423
rect 18236 22432 18288 22438
rect 18236 22374 18288 22380
rect 18234 22264 18290 22273
rect 18234 22199 18290 22208
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 18248 21434 18276 22199
rect 17880 21406 18000 21434
rect 18064 21406 18276 21434
rect 17880 21350 17908 21406
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 17682 20839 17738 20848
rect 17776 20868 17828 20874
rect 17696 18970 17724 20839
rect 17776 20810 17828 20816
rect 17880 20602 17908 20878
rect 17868 20596 17920 20602
rect 17868 20538 17920 20544
rect 17776 19984 17828 19990
rect 17776 19926 17828 19932
rect 17788 19174 17816 19926
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 17776 19168 17828 19174
rect 17774 19136 17776 19145
rect 17828 19136 17830 19145
rect 17774 19071 17830 19080
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17408 18828 17460 18834
rect 17512 18822 17724 18850
rect 17408 18770 17460 18776
rect 17420 18426 17448 18770
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17316 18148 17368 18154
rect 17316 18090 17368 18096
rect 17052 16782 17264 16810
rect 17052 16046 17080 16782
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 17144 15910 17172 16594
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17132 15904 17184 15910
rect 16960 15830 17080 15858
rect 17132 15846 17184 15852
rect 17052 14958 17080 15830
rect 17040 14952 17092 14958
rect 16854 14920 16910 14929
rect 17040 14894 17092 14900
rect 16854 14855 16910 14864
rect 16868 14822 16896 14855
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16868 14550 16896 14758
rect 16856 14544 16908 14550
rect 16856 14486 16908 14492
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16776 13938 16804 14418
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16776 12850 16804 13194
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16684 12294 16804 12322
rect 16578 12271 16580 12280
rect 16632 12271 16634 12280
rect 16580 12242 16632 12248
rect 16672 12232 16724 12238
rect 16670 12200 16672 12209
rect 16724 12200 16726 12209
rect 16670 12135 16726 12144
rect 16776 11393 16804 12294
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16762 11384 16818 11393
rect 16762 11319 16818 11328
rect 16868 11286 16896 11494
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16762 10568 16818 10577
rect 16762 10503 16764 10512
rect 16816 10503 16818 10512
rect 16764 10474 16816 10480
rect 16960 10452 16988 12582
rect 17052 10554 17080 14894
rect 17144 11121 17172 15846
rect 17236 15162 17264 16390
rect 17328 15366 17356 18090
rect 17420 15706 17448 18362
rect 17500 17740 17552 17746
rect 17500 17682 17552 17688
rect 17512 17338 17540 17682
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17604 16810 17632 17478
rect 17512 16782 17632 16810
rect 17512 16726 17540 16782
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17512 16114 17540 16662
rect 17696 16590 17724 18822
rect 17972 18630 18000 19246
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 17649 18000 18566
rect 17958 17640 18014 17649
rect 17958 17575 18014 17584
rect 18064 17082 18092 21406
rect 18234 21312 18290 21321
rect 18234 21247 18290 21256
rect 18142 21176 18198 21185
rect 18142 21111 18198 21120
rect 18156 21078 18184 21111
rect 18144 21072 18196 21078
rect 18144 21014 18196 21020
rect 18156 20058 18184 21014
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18156 17649 18184 18158
rect 18248 18034 18276 21247
rect 18340 20262 18368 25214
rect 18432 24138 18460 25978
rect 18524 24682 18552 26658
rect 18892 25770 18920 27520
rect 19248 25968 19300 25974
rect 19248 25910 19300 25916
rect 18880 25764 18932 25770
rect 18880 25706 18932 25712
rect 18604 25356 18656 25362
rect 18604 25298 18656 25304
rect 18696 25356 18748 25362
rect 18696 25298 18748 25304
rect 19064 25356 19116 25362
rect 19064 25298 19116 25304
rect 18616 24818 18644 25298
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18512 24676 18564 24682
rect 18512 24618 18564 24624
rect 18616 24206 18644 24754
rect 18708 24682 18736 25298
rect 18972 25288 19024 25294
rect 18972 25230 19024 25236
rect 18788 25152 18840 25158
rect 18788 25094 18840 25100
rect 18696 24676 18748 24682
rect 18696 24618 18748 24624
rect 18604 24200 18656 24206
rect 18604 24142 18656 24148
rect 18420 24132 18472 24138
rect 18420 24074 18472 24080
rect 18708 23497 18736 24618
rect 18800 24410 18828 25094
rect 18880 24880 18932 24886
rect 18880 24822 18932 24828
rect 18788 24404 18840 24410
rect 18788 24346 18840 24352
rect 18694 23488 18750 23497
rect 18694 23423 18750 23432
rect 18418 23080 18474 23089
rect 18418 23015 18474 23024
rect 18328 20256 18380 20262
rect 18328 20198 18380 20204
rect 18328 18352 18380 18358
rect 18326 18320 18328 18329
rect 18380 18320 18382 18329
rect 18326 18255 18382 18264
rect 18248 18006 18368 18034
rect 18234 17912 18290 17921
rect 18234 17847 18236 17856
rect 18288 17847 18290 17856
rect 18236 17818 18288 17824
rect 18142 17640 18198 17649
rect 18142 17575 18198 17584
rect 18248 17338 18276 17818
rect 18236 17332 18288 17338
rect 18236 17274 18288 17280
rect 18064 17054 18184 17082
rect 18052 16992 18104 16998
rect 17774 16960 17830 16969
rect 18052 16934 18104 16940
rect 17774 16895 17830 16904
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 17420 15026 17448 15642
rect 17512 15366 17540 16050
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 17406 14240 17462 14249
rect 17512 14226 17540 15302
rect 17462 14198 17540 14226
rect 17406 14175 17462 14184
rect 17420 14074 17448 14175
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17316 13456 17368 13462
rect 17314 13424 17316 13433
rect 17368 13424 17370 13433
rect 17314 13359 17370 13368
rect 17592 13320 17644 13326
rect 17498 13288 17554 13297
rect 17592 13262 17644 13268
rect 17498 13223 17500 13232
rect 17552 13223 17554 13232
rect 17500 13194 17552 13200
rect 17604 13138 17632 13262
rect 17512 13110 17632 13138
rect 17512 12918 17540 13110
rect 17500 12912 17552 12918
rect 17498 12880 17500 12889
rect 17592 12912 17644 12918
rect 17552 12880 17554 12889
rect 17592 12854 17644 12860
rect 17498 12815 17554 12824
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17420 11558 17448 12174
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17420 11354 17448 11494
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 17130 11112 17186 11121
rect 17130 11047 17186 11056
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17052 10526 17264 10554
rect 16960 10424 17080 10452
rect 16946 10296 17002 10305
rect 16580 10260 16632 10266
rect 16946 10231 17002 10240
rect 16580 10202 16632 10208
rect 16592 9024 16620 10202
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16868 9926 16896 10066
rect 16856 9920 16908 9926
rect 16854 9888 16856 9897
rect 16908 9888 16910 9897
rect 16854 9823 16910 9832
rect 16592 8996 16712 9024
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 15660 3878 15712 3884
rect 15764 3896 15884 3924
rect 16040 4270 16344 4298
rect 16408 6956 16528 6984
rect 15382 3768 15438 3777
rect 15382 3703 15438 3712
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15396 2990 15424 3470
rect 15488 3194 15516 3674
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15580 3194 15608 3334
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15764 3074 15792 3896
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 15856 3097 15884 3334
rect 15488 3046 15792 3074
rect 15842 3088 15898 3097
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15108 1624 15160 1630
rect 15106 1592 15108 1601
rect 15160 1592 15162 1601
rect 15106 1527 15162 1536
rect 15198 1320 15254 1329
rect 15198 1255 15254 1264
rect 14844 1006 14964 1034
rect 14936 480 14964 1006
rect 6274 439 6330 448
rect 6734 0 6790 480
rect 7286 0 7342 480
rect 7838 0 7894 480
rect 8390 0 8446 480
rect 8942 0 8998 480
rect 9494 0 9550 480
rect 10046 0 10102 480
rect 10598 0 10654 480
rect 11150 0 11206 480
rect 11702 0 11758 480
rect 12254 0 12310 480
rect 12806 0 12862 480
rect 13358 0 13414 480
rect 13910 0 13966 480
rect 14370 0 14426 480
rect 14832 264 14884 270
rect 14830 232 14832 241
rect 14884 232 14886 241
rect 14830 167 14886 176
rect 14922 0 14978 480
rect 15212 377 15240 1255
rect 15488 480 15516 3046
rect 15842 3023 15898 3032
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15580 2582 15608 2926
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 16040 480 16068 4270
rect 16408 4146 16436 6956
rect 16488 6860 16540 6866
rect 16592 6848 16620 8842
rect 16684 8430 16712 8996
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16854 7032 16910 7041
rect 16854 6967 16910 6976
rect 16540 6820 16620 6848
rect 16488 6802 16540 6808
rect 16592 6361 16620 6820
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16578 6352 16634 6361
rect 16578 6287 16634 6296
rect 16684 5914 16712 6802
rect 16762 6624 16818 6633
rect 16762 6559 16818 6568
rect 16776 6186 16804 6559
rect 16868 6458 16896 6967
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16868 6254 16896 6394
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16764 6180 16816 6186
rect 16764 6122 16816 6128
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16212 3936 16264 3942
rect 16212 3878 16264 3884
rect 16224 3233 16252 3878
rect 16302 3768 16358 3777
rect 16500 3738 16528 4966
rect 16960 4842 16988 10231
rect 16592 4814 16988 4842
rect 16302 3703 16304 3712
rect 16356 3703 16358 3712
rect 16488 3732 16540 3738
rect 16304 3674 16356 3680
rect 16488 3674 16540 3680
rect 16210 3224 16266 3233
rect 16210 3159 16266 3168
rect 16592 480 16620 4814
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16868 4146 16896 4422
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16762 3904 16818 3913
rect 16762 3839 16818 3848
rect 16776 3670 16804 3839
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16868 3534 16896 4082
rect 17052 3602 17080 10424
rect 17236 10130 17264 10526
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17236 9382 17264 10066
rect 17420 10062 17448 10610
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17236 8974 17264 9318
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17144 5846 17172 6258
rect 17132 5840 17184 5846
rect 17132 5782 17184 5788
rect 17144 5370 17172 5782
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17130 4720 17186 4729
rect 17236 4690 17264 8774
rect 17328 8673 17356 9998
rect 17420 9178 17448 9998
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17408 8832 17460 8838
rect 17408 8774 17460 8780
rect 17498 8800 17554 8809
rect 17314 8664 17370 8673
rect 17314 8599 17370 8608
rect 17328 8401 17356 8599
rect 17314 8392 17370 8401
rect 17314 8327 17370 8336
rect 17420 8294 17448 8774
rect 17498 8735 17554 8744
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 7750 17448 8230
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17420 5778 17448 6054
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17130 4655 17186 4664
rect 17224 4684 17276 4690
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16868 3126 16896 3470
rect 16856 3120 16908 3126
rect 16856 3062 16908 3068
rect 17052 2990 17080 3538
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16868 1873 16896 2246
rect 16854 1864 16910 1873
rect 16854 1799 16910 1808
rect 17038 640 17094 649
rect 17038 575 17094 584
rect 15198 368 15254 377
rect 15198 303 15254 312
rect 15474 0 15530 480
rect 16026 0 16082 480
rect 16578 0 16634 480
rect 17052 241 17080 575
rect 17144 480 17172 4655
rect 17224 4626 17276 4632
rect 17236 4078 17264 4626
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17236 3534 17264 4014
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17420 2961 17448 3334
rect 17406 2952 17462 2961
rect 17406 2887 17462 2896
rect 17512 2553 17540 8735
rect 17604 7478 17632 12854
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 17696 5370 17724 15982
rect 17788 14074 17816 16895
rect 17868 16516 17920 16522
rect 17868 16458 17920 16464
rect 17880 16182 17908 16458
rect 17868 16176 17920 16182
rect 17866 16144 17868 16153
rect 17920 16144 17922 16153
rect 17866 16079 17922 16088
rect 18064 15706 18092 16934
rect 18156 16425 18184 17054
rect 18142 16416 18198 16425
rect 18142 16351 18198 16360
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 18052 15700 18104 15706
rect 18052 15642 18104 15648
rect 17960 15564 18012 15570
rect 17880 15524 17960 15552
rect 17880 15162 17908 15524
rect 17960 15506 18012 15512
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 17880 14618 17908 14826
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17958 14104 18014 14113
rect 17776 14068 17828 14074
rect 17958 14039 18014 14048
rect 17776 14010 17828 14016
rect 17972 13802 18000 14039
rect 18064 13938 18092 14758
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 18156 13682 18184 15846
rect 18234 15464 18290 15473
rect 18234 15399 18236 15408
rect 18288 15399 18290 15408
rect 18236 15370 18288 15376
rect 17880 13654 18184 13682
rect 17880 13530 17908 13654
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17880 12442 17908 13330
rect 18340 12918 18368 18006
rect 18432 17202 18460 23015
rect 18800 22982 18828 24346
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18510 22808 18566 22817
rect 18510 22743 18566 22752
rect 18524 22642 18552 22743
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18616 22273 18644 22918
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18602 22264 18658 22273
rect 18602 22199 18658 22208
rect 18708 22166 18736 22578
rect 18696 22160 18748 22166
rect 18696 22102 18748 22108
rect 18892 22098 18920 24822
rect 18984 24818 19012 25230
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 18972 22976 19024 22982
rect 18972 22918 19024 22924
rect 18984 22574 19012 22918
rect 18972 22568 19024 22574
rect 18972 22510 19024 22516
rect 18970 22264 19026 22273
rect 18970 22199 19026 22208
rect 18512 22092 18564 22098
rect 18512 22034 18564 22040
rect 18880 22092 18932 22098
rect 18880 22034 18932 22040
rect 18524 21418 18552 22034
rect 18604 22024 18656 22030
rect 18604 21966 18656 21972
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18616 21690 18644 21966
rect 18604 21684 18656 21690
rect 18604 21626 18656 21632
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18512 21412 18564 21418
rect 18512 21354 18564 21360
rect 18524 21010 18552 21354
rect 18616 21350 18644 21490
rect 18708 21486 18736 21966
rect 18696 21480 18748 21486
rect 18696 21422 18748 21428
rect 18708 21350 18736 21422
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18512 21004 18564 21010
rect 18512 20946 18564 20952
rect 18512 20868 18564 20874
rect 18512 20810 18564 20816
rect 18524 20602 18552 20810
rect 18512 20596 18564 20602
rect 18512 20538 18564 20544
rect 18616 20466 18644 21286
rect 18708 21078 18736 21286
rect 18696 21072 18748 21078
rect 18696 21014 18748 21020
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18786 20088 18842 20097
rect 18984 20058 19012 22199
rect 18786 20023 18842 20032
rect 18972 20052 19024 20058
rect 18512 19916 18564 19922
rect 18512 19858 18564 19864
rect 18524 19174 18552 19858
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18616 19242 18644 19654
rect 18604 19236 18656 19242
rect 18604 19178 18656 19184
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18524 18873 18552 19110
rect 18510 18864 18566 18873
rect 18510 18799 18566 18808
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 18432 16794 18460 17138
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18524 16182 18552 18226
rect 18616 18193 18644 19178
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18602 18184 18658 18193
rect 18602 18119 18658 18128
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18616 17202 18644 17614
rect 18708 17513 18736 19110
rect 18800 17882 18828 20023
rect 18972 19994 19024 20000
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 18880 18624 18932 18630
rect 18880 18566 18932 18572
rect 18788 17876 18840 17882
rect 18788 17818 18840 17824
rect 18892 17785 18920 18566
rect 18984 18426 19012 19314
rect 19076 19310 19104 25298
rect 19260 25294 19288 25910
rect 19536 25498 19564 27520
rect 19984 25832 20036 25838
rect 19984 25774 20036 25780
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19996 25498 20024 25774
rect 19524 25492 19576 25498
rect 19524 25434 19576 25440
rect 19984 25492 20036 25498
rect 19984 25434 20036 25440
rect 19329 25392 19385 25401
rect 19329 25327 19385 25336
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 19154 24304 19210 24313
rect 19154 24239 19210 24248
rect 19168 22030 19196 24239
rect 19248 24064 19300 24070
rect 19248 24006 19300 24012
rect 19260 23338 19288 24006
rect 19352 23798 19380 25327
rect 19996 24750 20024 25434
rect 19984 24744 20036 24750
rect 19984 24686 20036 24692
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20088 23905 20116 27520
rect 20352 26580 20404 26586
rect 20352 26522 20404 26528
rect 20258 25800 20314 25809
rect 20258 25735 20314 25744
rect 20272 25537 20300 25735
rect 20258 25528 20314 25537
rect 20258 25463 20314 25472
rect 20364 25401 20392 26522
rect 20444 26308 20496 26314
rect 20444 26250 20496 26256
rect 20350 25392 20406 25401
rect 20350 25327 20406 25336
rect 20352 24812 20404 24818
rect 20352 24754 20404 24760
rect 20364 24070 20392 24754
rect 20456 24274 20484 26250
rect 20534 25800 20590 25809
rect 20534 25735 20590 25744
rect 20548 24857 20576 25735
rect 20640 25498 20668 27520
rect 20720 26852 20772 26858
rect 20720 26794 20772 26800
rect 20732 25838 20760 26794
rect 20904 25968 20956 25974
rect 20904 25910 20956 25916
rect 20996 25968 21048 25974
rect 20996 25910 21048 25916
rect 20720 25832 20772 25838
rect 20720 25774 20772 25780
rect 20732 25514 20760 25774
rect 20628 25492 20680 25498
rect 20732 25486 20852 25514
rect 20628 25434 20680 25440
rect 20720 25356 20772 25362
rect 20720 25298 20772 25304
rect 20628 24880 20680 24886
rect 20534 24848 20590 24857
rect 20628 24822 20680 24828
rect 20534 24783 20590 24792
rect 20536 24676 20588 24682
rect 20536 24618 20588 24624
rect 20444 24268 20496 24274
rect 20444 24210 20496 24216
rect 20352 24064 20404 24070
rect 20352 24006 20404 24012
rect 20074 23896 20130 23905
rect 20074 23831 20130 23840
rect 19340 23792 19392 23798
rect 19340 23734 19392 23740
rect 19524 23656 19576 23662
rect 19524 23598 19576 23604
rect 19982 23624 20038 23633
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 19260 23310 19380 23338
rect 19352 23186 19380 23310
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19248 22568 19300 22574
rect 19248 22510 19300 22516
rect 19260 22409 19288 22510
rect 19246 22400 19302 22409
rect 19246 22335 19302 22344
rect 19352 22080 19380 23122
rect 19444 22642 19472 23462
rect 19536 22778 19564 23598
rect 19982 23559 20038 23568
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19892 23248 19944 23254
rect 19892 23190 19944 23196
rect 19524 22772 19576 22778
rect 19524 22714 19576 22720
rect 19904 22710 19932 23190
rect 19616 22704 19668 22710
rect 19616 22646 19668 22652
rect 19892 22704 19944 22710
rect 19892 22646 19944 22652
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19430 22536 19486 22545
rect 19628 22522 19656 22646
rect 19800 22568 19852 22574
rect 19486 22494 19656 22522
rect 19798 22536 19800 22545
rect 19852 22536 19854 22545
rect 19430 22471 19486 22480
rect 19798 22471 19854 22480
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19996 22216 20024 23559
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 20180 23322 20208 23462
rect 20168 23316 20220 23322
rect 20168 23258 20220 23264
rect 20260 23248 20312 23254
rect 20260 23190 20312 23196
rect 20168 23112 20220 23118
rect 20168 23054 20220 23060
rect 20076 22772 20128 22778
rect 20076 22714 20128 22720
rect 20088 22574 20116 22714
rect 20076 22568 20128 22574
rect 20076 22510 20128 22516
rect 19628 22188 20024 22216
rect 20076 22228 20128 22234
rect 19352 22052 19472 22080
rect 19156 22024 19208 22030
rect 19156 21966 19208 21972
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19156 20936 19208 20942
rect 19156 20878 19208 20884
rect 19168 20097 19196 20878
rect 19260 20874 19288 21830
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19248 20868 19300 20874
rect 19248 20810 19300 20816
rect 19352 20398 19380 21286
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19154 20088 19210 20097
rect 19154 20023 19210 20032
rect 19248 19984 19300 19990
rect 19248 19926 19300 19932
rect 19352 19938 19380 20198
rect 19444 20058 19472 22052
rect 19628 21434 19656 22188
rect 20180 22216 20208 23054
rect 20272 22982 20300 23190
rect 20260 22976 20312 22982
rect 20260 22918 20312 22924
rect 20272 22234 20300 22918
rect 20128 22188 20208 22216
rect 20260 22228 20312 22234
rect 20076 22170 20128 22176
rect 20260 22170 20312 22176
rect 20364 22166 20392 24006
rect 20456 23594 20484 24210
rect 20548 23610 20576 24618
rect 20640 24410 20668 24822
rect 20732 24818 20760 25298
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20628 24404 20680 24410
rect 20628 24346 20680 24352
rect 20640 23730 20668 24346
rect 20720 24200 20772 24206
rect 20720 24142 20772 24148
rect 20732 23730 20760 24142
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20444 23588 20496 23594
rect 20548 23582 20668 23610
rect 20444 23530 20496 23536
rect 20456 23322 20484 23530
rect 20444 23316 20496 23322
rect 20444 23258 20496 23264
rect 20442 23080 20498 23089
rect 20442 23015 20498 23024
rect 20456 22982 20484 23015
rect 20444 22976 20496 22982
rect 20444 22918 20496 22924
rect 20444 22636 20496 22642
rect 20444 22578 20496 22584
rect 20352 22160 20404 22166
rect 20352 22102 20404 22108
rect 19708 22092 19760 22098
rect 19708 22034 19760 22040
rect 20168 22092 20220 22098
rect 20168 22034 20220 22040
rect 19720 21729 19748 22034
rect 19800 21956 19852 21962
rect 19800 21898 19852 21904
rect 20076 21956 20128 21962
rect 20076 21898 20128 21904
rect 19812 21865 19840 21898
rect 19892 21888 19944 21894
rect 19798 21856 19854 21865
rect 19892 21830 19944 21836
rect 19798 21791 19854 21800
rect 19706 21720 19762 21729
rect 19706 21655 19708 21664
rect 19760 21655 19762 21664
rect 19708 21626 19760 21632
rect 19720 21595 19748 21626
rect 19812 21554 19840 21791
rect 19904 21729 19932 21830
rect 19890 21720 19946 21729
rect 19890 21655 19946 21664
rect 19800 21548 19852 21554
rect 19800 21490 19852 21496
rect 19536 21406 19656 21434
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19064 19304 19116 19310
rect 19260 19258 19288 19926
rect 19352 19910 19472 19938
rect 19329 19816 19385 19825
rect 19385 19780 19392 19786
rect 19329 19751 19340 19760
rect 19340 19722 19392 19728
rect 19064 19246 19116 19252
rect 19168 19242 19380 19258
rect 19168 19236 19392 19242
rect 19168 19230 19340 19236
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 19076 18465 19104 18770
rect 19062 18456 19118 18465
rect 18972 18420 19024 18426
rect 19062 18391 19118 18400
rect 18972 18362 19024 18368
rect 18878 17776 18934 17785
rect 18878 17711 18934 17720
rect 18694 17504 18750 17513
rect 18694 17439 18750 17448
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18616 16726 18644 17138
rect 18604 16720 18656 16726
rect 18604 16662 18656 16668
rect 18984 16658 19012 18362
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 18970 16416 19026 16425
rect 18970 16351 19026 16360
rect 18512 16176 18564 16182
rect 18512 16118 18564 16124
rect 18696 16176 18748 16182
rect 18696 16118 18748 16124
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18432 14618 18460 15642
rect 18604 15360 18656 15366
rect 18510 15328 18566 15337
rect 18604 15302 18656 15308
rect 18510 15263 18566 15272
rect 18524 15026 18552 15263
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18524 14074 18552 14962
rect 18616 14822 18644 15302
rect 18708 14822 18736 16118
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18800 15094 18828 15438
rect 18788 15088 18840 15094
rect 18788 15030 18840 15036
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18696 14816 18748 14822
rect 18748 14776 18920 14804
rect 18696 14758 18748 14764
rect 18616 14521 18644 14758
rect 18694 14648 18750 14657
rect 18694 14583 18750 14592
rect 18602 14512 18658 14521
rect 18602 14447 18658 14456
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18512 14068 18564 14074
rect 18512 14010 18564 14016
rect 18512 13796 18564 13802
rect 18512 13738 18564 13744
rect 18524 13705 18552 13738
rect 18510 13696 18566 13705
rect 18510 13631 18566 13640
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18432 12986 18460 13330
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18510 12880 18566 12889
rect 18510 12815 18566 12824
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18234 12472 18290 12481
rect 17868 12436 17920 12442
rect 18234 12407 18290 12416
rect 17868 12378 17920 12384
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 18064 11665 18092 12174
rect 18050 11656 18106 11665
rect 18050 11591 18106 11600
rect 17958 11248 18014 11257
rect 17958 11183 18014 11192
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17788 9722 17816 10542
rect 17880 10441 17908 10678
rect 17866 10432 17922 10441
rect 17866 10367 17922 10376
rect 17972 10198 18000 11183
rect 18248 10606 18276 12407
rect 18432 12238 18460 12582
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18326 11248 18382 11257
rect 18326 11183 18382 11192
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 18064 10033 18092 10406
rect 18050 10024 18106 10033
rect 18050 9959 18106 9968
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17788 9518 17816 9658
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17972 9450 18000 9862
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 18052 9036 18104 9042
rect 18052 8978 18104 8984
rect 17972 7426 18000 8978
rect 18064 7546 18092 8978
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 17972 7398 18092 7426
rect 17958 6896 18014 6905
rect 17868 6860 17920 6866
rect 17958 6831 17960 6840
rect 17868 6802 17920 6808
rect 18012 6831 18014 6840
rect 17960 6802 18012 6808
rect 17880 6390 17908 6802
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17868 6384 17920 6390
rect 17868 6326 17920 6332
rect 17972 6322 18000 6598
rect 18064 6497 18092 7398
rect 18050 6488 18106 6497
rect 18050 6423 18106 6432
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 18052 6180 18104 6186
rect 18052 6122 18104 6128
rect 18064 5574 18092 6122
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17868 4752 17920 4758
rect 17868 4694 17920 4700
rect 17880 4593 17908 4694
rect 17682 4584 17738 4593
rect 17682 4519 17738 4528
rect 17866 4584 17922 4593
rect 17866 4519 17922 4528
rect 17592 3664 17644 3670
rect 17592 3606 17644 3612
rect 17604 2990 17632 3606
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17314 2544 17370 2553
rect 17314 2479 17370 2488
rect 17498 2544 17554 2553
rect 17498 2479 17554 2488
rect 17328 2281 17356 2479
rect 17314 2272 17370 2281
rect 17314 2207 17370 2216
rect 17408 2100 17460 2106
rect 17408 2042 17460 2048
rect 17314 1184 17370 1193
rect 17314 1119 17370 1128
rect 17328 785 17356 1119
rect 17420 921 17448 2042
rect 17500 1896 17552 1902
rect 17498 1864 17500 1873
rect 17552 1864 17554 1873
rect 17498 1799 17554 1808
rect 17406 912 17462 921
rect 17406 847 17462 856
rect 17314 776 17370 785
rect 17314 711 17370 720
rect 17696 480 17724 4519
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18064 3777 18092 3878
rect 18050 3768 18106 3777
rect 18050 3703 18106 3712
rect 17776 3664 17828 3670
rect 17774 3632 17776 3641
rect 17828 3632 17830 3641
rect 17774 3567 17830 3576
rect 17960 3528 18012 3534
rect 18156 3505 18184 10474
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 18248 9926 18276 10406
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18340 9466 18368 11183
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 18432 10674 18460 10950
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18420 10464 18472 10470
rect 18524 10452 18552 12815
rect 18472 10424 18552 10452
rect 18420 10406 18472 10412
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18432 9761 18460 9862
rect 18418 9752 18474 9761
rect 18616 9704 18644 14350
rect 18418 9687 18474 9696
rect 18524 9676 18644 9704
rect 18340 9438 18460 9466
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18248 8090 18276 8910
rect 18340 8673 18368 9318
rect 18326 8664 18382 8673
rect 18326 8599 18382 8608
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18248 7750 18276 7822
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18248 6798 18276 7686
rect 18432 7290 18460 9438
rect 18524 8022 18552 9676
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18616 8974 18644 9522
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18512 8016 18564 8022
rect 18512 7958 18564 7964
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18524 7478 18552 7754
rect 18512 7472 18564 7478
rect 18512 7414 18564 7420
rect 18340 7262 18460 7290
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18234 6352 18290 6361
rect 18234 6287 18236 6296
rect 18288 6287 18290 6296
rect 18236 6258 18288 6264
rect 18234 5672 18290 5681
rect 18234 5607 18236 5616
rect 18288 5607 18290 5616
rect 18236 5578 18288 5584
rect 18340 5302 18368 7262
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18432 7041 18460 7142
rect 18418 7032 18474 7041
rect 18418 6967 18474 6976
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18432 5953 18460 6190
rect 18418 5944 18474 5953
rect 18418 5879 18474 5888
rect 18328 5296 18380 5302
rect 18328 5238 18380 5244
rect 18340 5030 18368 5238
rect 18420 5160 18472 5166
rect 18420 5102 18472 5108
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 18432 4690 18460 5102
rect 18420 4684 18472 4690
rect 18420 4626 18472 4632
rect 18432 4214 18460 4626
rect 18524 4321 18552 7414
rect 18616 7410 18644 7822
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18708 7002 18736 14583
rect 18892 14006 18920 14776
rect 18984 14414 19012 16351
rect 19076 16250 19104 18391
rect 19168 17338 19196 19230
rect 19340 19178 19392 19184
rect 19248 19168 19300 19174
rect 19444 19156 19472 19910
rect 19536 19310 19564 21406
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 19996 20505 20024 20946
rect 19982 20496 20038 20505
rect 19982 20431 20038 20440
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19524 19304 19576 19310
rect 19524 19246 19576 19252
rect 19444 19128 19564 19156
rect 19300 19116 19380 19122
rect 19248 19110 19380 19116
rect 19260 19094 19380 19110
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19260 17882 19288 18158
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19248 17740 19300 17746
rect 19248 17682 19300 17688
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 19168 17066 19196 17274
rect 19156 17060 19208 17066
rect 19156 17002 19208 17008
rect 19260 16833 19288 17682
rect 19246 16824 19302 16833
rect 19246 16759 19248 16768
rect 19300 16759 19302 16768
rect 19248 16730 19300 16736
rect 19352 16674 19380 19094
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19444 18426 19472 18702
rect 19432 18420 19484 18426
rect 19432 18362 19484 18368
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 19444 16969 19472 17546
rect 19430 16960 19486 16969
rect 19430 16895 19486 16904
rect 19444 16794 19472 16895
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19156 16652 19208 16658
rect 19352 16646 19472 16674
rect 19156 16594 19208 16600
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 19168 15978 19196 16594
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19156 15972 19208 15978
rect 19156 15914 19208 15920
rect 19062 15328 19118 15337
rect 19062 15263 19118 15272
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 18880 14000 18932 14006
rect 18880 13942 18932 13948
rect 18788 13728 18840 13734
rect 18788 13670 18840 13676
rect 18800 13025 18828 13670
rect 18892 13462 18920 13942
rect 19076 13530 19104 15263
rect 19168 14346 19196 15914
rect 19352 15706 19380 16458
rect 19444 15978 19472 16646
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19430 15872 19486 15881
rect 19430 15807 19486 15816
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19248 15632 19300 15638
rect 19248 15574 19300 15580
rect 19260 14618 19288 15574
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19156 14340 19208 14346
rect 19156 14282 19208 14288
rect 19260 14074 19288 14350
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19156 13728 19208 13734
rect 19156 13670 19208 13676
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 18880 13456 18932 13462
rect 18932 13416 19012 13444
rect 18880 13398 18932 13404
rect 18786 13016 18842 13025
rect 18786 12951 18842 12960
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 18892 12617 18920 12922
rect 18984 12782 19012 13416
rect 19168 13410 19196 13670
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19076 13382 19196 13410
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18878 12608 18934 12617
rect 18878 12543 18934 12552
rect 18984 12442 19012 12718
rect 19076 12481 19104 13382
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 19168 12714 19196 13194
rect 19260 12986 19288 13466
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19156 12708 19208 12714
rect 19156 12650 19208 12656
rect 19062 12472 19118 12481
rect 18972 12436 19024 12442
rect 19062 12407 19118 12416
rect 18972 12378 19024 12384
rect 18984 11898 19012 12378
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 18786 11520 18842 11529
rect 18786 11455 18842 11464
rect 18800 10538 18828 11455
rect 18972 11212 19024 11218
rect 18972 11154 19024 11160
rect 18880 11076 18932 11082
rect 18880 11018 18932 11024
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18892 10169 18920 11018
rect 18984 10849 19012 11154
rect 18970 10840 19026 10849
rect 18970 10775 18972 10784
rect 19024 10775 19026 10784
rect 18972 10746 19024 10752
rect 19076 10169 19104 12242
rect 19168 12170 19196 12650
rect 19352 12594 19380 15506
rect 19444 13988 19472 15807
rect 19536 15570 19564 19128
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19996 17882 20024 20431
rect 20088 19446 20116 21898
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 20074 19136 20130 19145
rect 20074 19071 20130 19080
rect 20088 18970 20116 19071
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 20076 18692 20128 18698
rect 20076 18634 20128 18640
rect 20088 18601 20116 18634
rect 20074 18592 20130 18601
rect 20074 18527 20130 18536
rect 19984 17876 20036 17882
rect 19984 17818 20036 17824
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19720 17066 19748 17478
rect 19996 17105 20024 17478
rect 19982 17096 20038 17105
rect 19708 17060 19760 17066
rect 19982 17031 20038 17040
rect 19708 17002 19760 17008
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19614 16688 19670 16697
rect 19614 16623 19616 16632
rect 19668 16623 19670 16632
rect 19616 16594 19668 16600
rect 20088 16096 20116 17614
rect 19996 16068 20116 16096
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19524 15564 19576 15570
rect 19524 15506 19576 15512
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19522 15192 19578 15201
rect 19522 15127 19578 15136
rect 19536 14618 19564 15127
rect 19904 14958 19932 15302
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19536 14056 19564 14554
rect 19616 14068 19668 14074
rect 19536 14028 19616 14056
rect 19616 14010 19668 14016
rect 19444 13960 19564 13988
rect 19536 13410 19564 13960
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19996 13546 20024 16068
rect 20076 15972 20128 15978
rect 20076 15914 20128 15920
rect 20088 14482 20116 15914
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 20076 13728 20128 13734
rect 20074 13696 20076 13705
rect 20128 13696 20130 13705
rect 20074 13631 20130 13640
rect 19996 13518 20116 13546
rect 19800 13456 19852 13462
rect 19432 13388 19484 13394
rect 19536 13382 19656 13410
rect 19800 13398 19852 13404
rect 19432 13330 19484 13336
rect 19444 12866 19472 13330
rect 19444 12838 19564 12866
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19260 12566 19380 12594
rect 19260 12322 19288 12566
rect 19338 12472 19394 12481
rect 19444 12442 19472 12718
rect 19338 12407 19340 12416
rect 19392 12407 19394 12416
rect 19432 12436 19484 12442
rect 19340 12378 19392 12384
rect 19432 12378 19484 12384
rect 19260 12294 19380 12322
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19156 12164 19208 12170
rect 19156 12106 19208 12112
rect 19168 11558 19196 12106
rect 19260 12102 19288 12174
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19156 11552 19208 11558
rect 19260 11529 19288 11562
rect 19156 11494 19208 11500
rect 19246 11520 19302 11529
rect 19246 11455 19302 11464
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 18878 10160 18934 10169
rect 18788 10124 18840 10130
rect 18878 10095 18934 10104
rect 19062 10160 19118 10169
rect 19062 10095 19118 10104
rect 18788 10066 18840 10072
rect 18800 9217 18828 10066
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 18880 9988 18932 9994
rect 18880 9930 18932 9936
rect 18786 9208 18842 9217
rect 18786 9143 18788 9152
rect 18840 9143 18842 9152
rect 18788 9114 18840 9120
rect 18786 8800 18842 8809
rect 18786 8735 18842 8744
rect 18800 7206 18828 8735
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18604 6928 18656 6934
rect 18604 6870 18656 6876
rect 18616 4758 18644 6870
rect 18604 4752 18656 4758
rect 18604 4694 18656 4700
rect 18510 4312 18566 4321
rect 18510 4247 18566 4256
rect 18420 4208 18472 4214
rect 18420 4150 18472 4156
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 17960 3470 18012 3476
rect 18142 3496 18198 3505
rect 17972 3194 18000 3470
rect 18142 3431 18198 3440
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18156 3074 18184 3431
rect 17972 3046 18184 3074
rect 17972 1630 18000 3046
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 18052 2848 18104 2854
rect 18050 2816 18052 2825
rect 18104 2816 18106 2825
rect 18050 2751 18106 2760
rect 18156 2582 18184 2926
rect 18144 2576 18196 2582
rect 18144 2518 18196 2524
rect 17960 1624 18012 1630
rect 17960 1566 18012 1572
rect 18248 1442 18276 4014
rect 18616 3738 18644 4694
rect 18800 4554 18828 7142
rect 18892 4826 18920 9930
rect 18984 9586 19012 9998
rect 19076 9722 19104 9998
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 19168 9489 19196 11290
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19154 9480 19210 9489
rect 19154 9415 19210 9424
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18984 6934 19012 9318
rect 19064 8560 19116 8566
rect 19064 8502 19116 8508
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 19076 6746 19104 8502
rect 19260 8242 19288 10406
rect 19168 8214 19288 8242
rect 19168 7041 19196 8214
rect 19352 7954 19380 12294
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19444 11642 19472 12242
rect 19536 11762 19564 12838
rect 19628 12714 19656 13382
rect 19812 12986 19840 13398
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 19616 12708 19668 12714
rect 19616 12650 19668 12656
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19444 11614 19564 11642
rect 19628 11626 19656 12174
rect 19996 12073 20024 12786
rect 19982 12064 20038 12073
rect 19982 11999 20038 12008
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19444 11286 19472 11494
rect 19432 11280 19484 11286
rect 19432 11222 19484 11228
rect 19536 11234 19564 11614
rect 19616 11620 19668 11626
rect 19616 11562 19668 11568
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19536 11218 19748 11234
rect 19536 11212 19760 11218
rect 19536 11206 19708 11212
rect 19708 11154 19760 11160
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19522 11112 19578 11121
rect 19444 10810 19472 11086
rect 19522 11047 19578 11056
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19444 10470 19472 10746
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19430 10296 19486 10305
rect 19430 10231 19432 10240
rect 19484 10231 19486 10240
rect 19432 10202 19484 10208
rect 19430 9344 19486 9353
rect 19430 9279 19486 9288
rect 19444 9110 19472 9279
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19430 8936 19486 8945
rect 19430 8871 19486 8880
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19154 7032 19210 7041
rect 19154 6967 19210 6976
rect 19156 6860 19208 6866
rect 19156 6802 19208 6808
rect 18984 6718 19104 6746
rect 18984 6322 19012 6718
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 19076 6225 19104 6598
rect 19062 6216 19118 6225
rect 19062 6151 19118 6160
rect 19168 5914 19196 6802
rect 19260 6254 19288 7822
rect 19352 7546 19380 7890
rect 19444 7721 19472 8871
rect 19430 7712 19486 7721
rect 19430 7647 19486 7656
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19340 7268 19392 7274
rect 19340 7210 19392 7216
rect 19352 7177 19380 7210
rect 19444 7206 19472 7647
rect 19432 7200 19484 7206
rect 19338 7168 19394 7177
rect 19432 7142 19484 7148
rect 19338 7103 19394 7112
rect 19430 7032 19486 7041
rect 19340 6996 19392 7002
rect 19430 6967 19486 6976
rect 19340 6938 19392 6944
rect 19352 6662 19380 6938
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19444 6254 19472 6967
rect 19536 6322 19564 11047
rect 19800 11008 19852 11014
rect 19798 10976 19800 10985
rect 19852 10976 19854 10985
rect 19798 10911 19854 10920
rect 19904 10674 19932 11154
rect 19892 10668 19944 10674
rect 19892 10610 19944 10616
rect 19996 10470 20024 11698
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19996 10266 20024 10406
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19984 8968 20036 8974
rect 19614 8936 19670 8945
rect 19984 8910 20036 8916
rect 19614 8871 19616 8880
rect 19668 8871 19670 8880
rect 19616 8842 19668 8848
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19996 7936 20024 8910
rect 19812 7908 20024 7936
rect 19812 7188 19840 7908
rect 19890 7848 19946 7857
rect 19890 7783 19892 7792
rect 19944 7783 19946 7792
rect 19892 7754 19944 7760
rect 19904 7410 19932 7754
rect 19982 7440 20038 7449
rect 19892 7404 19944 7410
rect 19982 7375 20038 7384
rect 19892 7346 19944 7352
rect 19996 7342 20024 7375
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19812 7160 20024 7188
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19616 6792 19668 6798
rect 19996 6780 20024 7160
rect 19668 6752 20024 6780
rect 19616 6734 19668 6740
rect 19628 6390 19656 6734
rect 19616 6384 19668 6390
rect 19616 6326 19668 6332
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19156 5908 19208 5914
rect 19156 5850 19208 5856
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18788 4548 18840 4554
rect 18788 4490 18840 4496
rect 18696 4480 18748 4486
rect 18696 4422 18748 4428
rect 18708 4214 18736 4422
rect 18696 4208 18748 4214
rect 18696 4150 18748 4156
rect 18892 4078 18920 4762
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 18984 4282 19012 4626
rect 18972 4276 19024 4282
rect 18972 4218 19024 4224
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18418 3224 18474 3233
rect 18418 3159 18474 3168
rect 18602 3224 18658 3233
rect 18602 3159 18658 3168
rect 18788 3188 18840 3194
rect 18432 2990 18460 3159
rect 18510 3088 18566 3097
rect 18510 3023 18566 3032
rect 18524 2990 18552 3023
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 18340 1465 18368 2246
rect 18156 1414 18276 1442
rect 18326 1456 18382 1465
rect 17038 232 17094 241
rect 17038 167 17094 176
rect 17130 0 17186 480
rect 17682 0 17738 480
rect 18156 270 18184 1414
rect 18326 1391 18382 1400
rect 18432 1329 18460 2926
rect 18616 2922 18644 3159
rect 18788 3130 18840 3136
rect 18604 2916 18656 2922
rect 18604 2858 18656 2864
rect 18696 2372 18748 2378
rect 18696 2314 18748 2320
rect 18708 2009 18736 2314
rect 18694 2000 18750 2009
rect 18694 1935 18750 1944
rect 18234 1320 18290 1329
rect 18234 1255 18290 1264
rect 18418 1320 18474 1329
rect 18418 1255 18474 1264
rect 18248 480 18276 1255
rect 18800 480 18828 3130
rect 18984 2650 19012 4218
rect 19076 3738 19104 5102
rect 19154 4856 19210 4865
rect 19154 4791 19210 4800
rect 19168 4622 19196 4791
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19352 4162 19380 5510
rect 19260 4134 19380 4162
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 19260 3194 19288 4134
rect 19444 4026 19472 6054
rect 19536 5914 19564 6054
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19996 5846 20024 6258
rect 19984 5840 20036 5846
rect 19984 5782 20036 5788
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19536 5370 19564 5714
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19996 4486 20024 5306
rect 19984 4480 20036 4486
rect 19522 4448 19578 4457
rect 19984 4422 20036 4428
rect 19522 4383 19578 4392
rect 19352 3998 19472 4026
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 19352 1578 19380 3998
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19444 2689 19472 3878
rect 19536 3670 19564 4383
rect 19996 4214 20024 4422
rect 19984 4208 20036 4214
rect 19984 4150 20036 4156
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19524 3664 19576 3670
rect 19524 3606 19576 3612
rect 19996 3534 20024 4150
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 19984 3392 20036 3398
rect 19982 3360 19984 3369
rect 20036 3360 20038 3369
rect 19982 3295 20038 3304
rect 19996 3126 20024 3295
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 20088 3058 20116 13518
rect 20180 12782 20208 22034
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 20352 22024 20404 22030
rect 20352 21966 20404 21972
rect 20272 21026 20300 21966
rect 20364 21146 20392 21966
rect 20456 21554 20484 22578
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 20272 20998 20392 21026
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 20272 19553 20300 20878
rect 20258 19544 20314 19553
rect 20258 19479 20260 19488
rect 20312 19479 20314 19488
rect 20260 19450 20312 19456
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20272 18834 20300 19110
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 20272 16794 20300 18770
rect 20364 17678 20392 20998
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 20456 19718 20484 20198
rect 20444 19712 20496 19718
rect 20444 19654 20496 19660
rect 20548 19666 20576 21830
rect 20640 21593 20668 23582
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20732 22710 20760 23054
rect 20720 22704 20772 22710
rect 20718 22672 20720 22681
rect 20772 22672 20774 22681
rect 20718 22607 20774 22616
rect 20720 22568 20772 22574
rect 20720 22510 20772 22516
rect 20732 22098 20760 22510
rect 20720 22092 20772 22098
rect 20720 22034 20772 22040
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 20626 21584 20682 21593
rect 20626 21519 20682 21528
rect 20732 21457 20760 21830
rect 20718 21448 20774 21457
rect 20718 21383 20774 21392
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20640 20942 20668 21286
rect 20718 21176 20774 21185
rect 20718 21111 20774 21120
rect 20628 20936 20680 20942
rect 20628 20878 20680 20884
rect 20732 20754 20760 21111
rect 20824 21078 20852 25486
rect 20916 22964 20944 25910
rect 21008 24342 21036 25910
rect 21284 25430 21312 27520
rect 21364 26240 21416 26246
rect 21364 26182 21416 26188
rect 21272 25424 21324 25430
rect 21272 25366 21324 25372
rect 21180 25356 21232 25362
rect 21180 25298 21232 25304
rect 21086 24712 21142 24721
rect 21086 24647 21142 24656
rect 20996 24336 21048 24342
rect 20996 24278 21048 24284
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 21008 23361 21036 23462
rect 20994 23352 21050 23361
rect 20994 23287 21050 23296
rect 21008 23089 21036 23287
rect 20994 23080 21050 23089
rect 20994 23015 21050 23024
rect 20916 22936 21036 22964
rect 21008 22778 21036 22936
rect 20996 22772 21048 22778
rect 20996 22714 21048 22720
rect 21008 22574 21036 22714
rect 20996 22568 21048 22574
rect 20996 22510 21048 22516
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20916 21146 20944 21490
rect 20904 21140 20956 21146
rect 20904 21082 20956 21088
rect 20812 21072 20864 21078
rect 20812 21014 20864 21020
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20732 20726 20852 20754
rect 20718 20632 20774 20641
rect 20718 20567 20774 20576
rect 20732 20330 20760 20567
rect 20720 20324 20772 20330
rect 20720 20266 20772 20272
rect 20720 19780 20772 19786
rect 20720 19722 20772 19728
rect 20456 19378 20484 19654
rect 20548 19638 20668 19666
rect 20534 19544 20590 19553
rect 20534 19479 20590 19488
rect 20444 19372 20496 19378
rect 20444 19314 20496 19320
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20456 18630 20484 19110
rect 20444 18624 20496 18630
rect 20442 18592 20444 18601
rect 20496 18592 20498 18601
rect 20442 18527 20498 18536
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20444 17536 20496 17542
rect 20350 17504 20406 17513
rect 20444 17478 20496 17484
rect 20350 17439 20406 17448
rect 20260 16788 20312 16794
rect 20260 16730 20312 16736
rect 20364 15706 20392 17439
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20272 14929 20300 15098
rect 20258 14920 20314 14929
rect 20258 14855 20260 14864
rect 20312 14855 20314 14864
rect 20260 14826 20312 14832
rect 20456 14822 20484 17478
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20260 14340 20312 14346
rect 20260 14282 20312 14288
rect 20272 12850 20300 14282
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20364 13802 20392 14214
rect 20456 13954 20484 14758
rect 20548 14346 20576 19479
rect 20640 18698 20668 19638
rect 20732 19446 20760 19722
rect 20720 19440 20772 19446
rect 20720 19382 20772 19388
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20640 17542 20668 18634
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20628 17060 20680 17066
rect 20628 17002 20680 17008
rect 20640 16794 20668 17002
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20640 16522 20668 16730
rect 20732 16590 20760 16934
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20628 16516 20680 16522
rect 20628 16458 20680 16464
rect 20640 16250 20668 16458
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20640 15706 20668 16186
rect 20628 15700 20680 15706
rect 20628 15642 20680 15648
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20640 14414 20668 15438
rect 20824 14890 20852 20726
rect 20916 19854 20944 20878
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20916 19174 20944 19790
rect 21008 19310 21036 22374
rect 21100 21690 21128 24647
rect 21192 24614 21220 25298
rect 21180 24608 21232 24614
rect 21180 24550 21232 24556
rect 21272 24268 21324 24274
rect 21272 24210 21324 24216
rect 21284 23866 21312 24210
rect 21376 24206 21404 26182
rect 21836 25242 21864 27520
rect 22388 25514 22416 27520
rect 22928 26104 22980 26110
rect 22928 26046 22980 26052
rect 22744 25968 22796 25974
rect 22744 25910 22796 25916
rect 22204 25486 22416 25514
rect 21836 25214 21956 25242
rect 21732 25152 21784 25158
rect 21732 25094 21784 25100
rect 21744 24750 21772 25094
rect 21822 24848 21878 24857
rect 21822 24783 21878 24792
rect 21732 24744 21784 24750
rect 21732 24686 21784 24692
rect 21640 24608 21692 24614
rect 21640 24550 21692 24556
rect 21364 24200 21416 24206
rect 21364 24142 21416 24148
rect 21272 23860 21324 23866
rect 21272 23802 21324 23808
rect 21376 23594 21404 24142
rect 21548 24064 21600 24070
rect 21548 24006 21600 24012
rect 21364 23588 21416 23594
rect 21364 23530 21416 23536
rect 21272 23180 21324 23186
rect 21272 23122 21324 23128
rect 21456 23180 21508 23186
rect 21456 23122 21508 23128
rect 21178 23080 21234 23089
rect 21178 23015 21234 23024
rect 21192 22545 21220 23015
rect 21178 22536 21234 22545
rect 21178 22471 21234 22480
rect 21284 22234 21312 23122
rect 21468 22642 21496 23122
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 21272 22228 21324 22234
rect 21272 22170 21324 22176
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 21180 21480 21232 21486
rect 21180 21422 21232 21428
rect 21088 21412 21140 21418
rect 21088 21354 21140 21360
rect 20996 19304 21048 19310
rect 20996 19246 21048 19252
rect 20904 19168 20956 19174
rect 21100 19156 21128 21354
rect 21192 21146 21220 21422
rect 21180 21140 21232 21146
rect 21180 21082 21232 21088
rect 21376 20806 21404 22374
rect 21468 21622 21496 22578
rect 21560 21865 21588 24006
rect 21546 21856 21602 21865
rect 21546 21791 21602 21800
rect 21652 21706 21680 24550
rect 21744 22420 21772 24686
rect 21836 24614 21864 24783
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21824 24064 21876 24070
rect 21824 24006 21876 24012
rect 21836 23730 21864 24006
rect 21928 23866 21956 25214
rect 21916 23860 21968 23866
rect 21916 23802 21968 23808
rect 21824 23724 21876 23730
rect 21824 23666 21876 23672
rect 21916 23656 21968 23662
rect 21916 23598 21968 23604
rect 21824 23316 21876 23322
rect 21824 23258 21876 23264
rect 21836 22574 21864 23258
rect 21824 22568 21876 22574
rect 21824 22510 21876 22516
rect 21744 22392 21864 22420
rect 21732 22024 21784 22030
rect 21732 21966 21784 21972
rect 21560 21678 21680 21706
rect 21456 21616 21508 21622
rect 21456 21558 21508 21564
rect 21468 21010 21496 21558
rect 21560 21185 21588 21678
rect 21744 21350 21772 21966
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21546 21176 21602 21185
rect 21546 21111 21602 21120
rect 21548 21072 21600 21078
rect 21548 21014 21600 21020
rect 21456 21004 21508 21010
rect 21456 20946 21508 20952
rect 21364 20800 21416 20806
rect 21364 20742 21416 20748
rect 21468 20602 21496 20946
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 21560 20466 21588 21014
rect 21548 20460 21600 20466
rect 21548 20402 21600 20408
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21638 20224 21694 20233
rect 21272 19984 21324 19990
rect 21272 19926 21324 19932
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 20904 19110 20956 19116
rect 21008 19128 21128 19156
rect 20902 18864 20958 18873
rect 21008 18834 21036 19128
rect 21086 18864 21142 18873
rect 20902 18799 20958 18808
rect 20996 18828 21048 18834
rect 20916 18086 20944 18799
rect 21086 18799 21142 18808
rect 20996 18770 21048 18776
rect 21008 18154 21036 18770
rect 20996 18148 21048 18154
rect 20996 18090 21048 18096
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20996 16720 21048 16726
rect 20996 16662 21048 16668
rect 20902 16416 20958 16425
rect 20902 16351 20958 16360
rect 20916 16250 20944 16351
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 21008 15638 21036 16662
rect 20996 15632 21048 15638
rect 20996 15574 21048 15580
rect 20996 15428 21048 15434
rect 20996 15370 21048 15376
rect 20812 14884 20864 14890
rect 20812 14826 20864 14832
rect 20902 14512 20958 14521
rect 20720 14476 20772 14482
rect 21008 14498 21036 15370
rect 21100 14618 21128 18799
rect 21192 18290 21220 19314
rect 21284 19242 21312 19926
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 21468 19258 21496 19450
rect 21560 19417 21588 20198
rect 21638 20159 21694 20168
rect 21546 19408 21602 19417
rect 21546 19343 21602 19352
rect 21272 19236 21324 19242
rect 21272 19178 21324 19184
rect 21376 19230 21496 19258
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 21180 17740 21232 17746
rect 21180 17682 21232 17688
rect 21192 17513 21220 17682
rect 21178 17504 21234 17513
rect 21178 17439 21234 17448
rect 21284 16998 21312 19178
rect 21376 17338 21404 19230
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21468 18601 21496 18702
rect 21560 18630 21588 19110
rect 21652 18986 21680 20159
rect 21730 19272 21786 19281
rect 21730 19207 21786 19216
rect 21744 19174 21772 19207
rect 21732 19168 21784 19174
rect 21732 19110 21784 19116
rect 21652 18958 21772 18986
rect 21548 18624 21600 18630
rect 21454 18592 21510 18601
rect 21548 18566 21600 18572
rect 21454 18527 21510 18536
rect 21468 17882 21496 18527
rect 21638 18456 21694 18465
rect 21638 18391 21640 18400
rect 21692 18391 21694 18400
rect 21640 18362 21692 18368
rect 21640 18284 21692 18290
rect 21640 18226 21692 18232
rect 21546 17912 21602 17921
rect 21456 17876 21508 17882
rect 21546 17847 21602 17856
rect 21456 17818 21508 17824
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21362 17232 21418 17241
rect 21362 17167 21418 17176
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 21270 16824 21326 16833
rect 21270 16759 21272 16768
rect 21324 16759 21326 16768
rect 21272 16730 21324 16736
rect 21284 15706 21312 16730
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 21180 15632 21232 15638
rect 21180 15574 21232 15580
rect 21192 14872 21220 15574
rect 21192 14844 21312 14872
rect 21178 14784 21234 14793
rect 21178 14719 21234 14728
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21008 14470 21128 14498
rect 20902 14447 20958 14456
rect 20720 14418 20772 14424
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 20626 14104 20682 14113
rect 20626 14039 20682 14048
rect 20456 13926 20576 13954
rect 20640 13938 20668 14039
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 20352 13796 20404 13802
rect 20352 13738 20404 13744
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20168 12776 20220 12782
rect 20168 12718 20220 12724
rect 20168 12640 20220 12646
rect 20168 12582 20220 12588
rect 20258 12608 20314 12617
rect 20180 10810 20208 12582
rect 20364 12594 20392 13738
rect 20314 12566 20392 12594
rect 20258 12543 20314 12552
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20168 10668 20220 10674
rect 20168 10610 20220 10616
rect 20180 10198 20208 10610
rect 20168 10192 20220 10198
rect 20168 10134 20220 10140
rect 20272 9586 20300 12543
rect 20350 12064 20406 12073
rect 20350 11999 20406 12008
rect 20364 11218 20392 11999
rect 20352 11212 20404 11218
rect 20352 11154 20404 11160
rect 20350 10840 20406 10849
rect 20350 10775 20406 10784
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20272 9178 20300 9522
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 20180 8809 20208 8978
rect 20166 8800 20222 8809
rect 20166 8735 20222 8744
rect 20180 8634 20208 8735
rect 20168 8628 20220 8634
rect 20168 8570 20220 8576
rect 20258 8120 20314 8129
rect 20258 8055 20314 8064
rect 20166 7848 20222 7857
rect 20166 7783 20222 7792
rect 20180 7274 20208 7783
rect 20272 7410 20300 8055
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20168 7268 20220 7274
rect 20364 7256 20392 10775
rect 20456 10742 20484 13806
rect 20548 13682 20576 13926
rect 20628 13932 20680 13938
rect 20628 13874 20680 13880
rect 20626 13832 20682 13841
rect 20626 13767 20682 13776
rect 20640 13682 20668 13767
rect 20732 13705 20760 14418
rect 20810 14240 20866 14249
rect 20810 14175 20866 14184
rect 20824 14074 20852 14175
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20548 13654 20668 13682
rect 20640 13394 20668 13654
rect 20718 13696 20774 13705
rect 20718 13631 20774 13640
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20626 13288 20682 13297
rect 20626 13223 20682 13232
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 20444 10736 20496 10742
rect 20444 10678 20496 10684
rect 20442 10296 20498 10305
rect 20442 10231 20498 10240
rect 20456 10130 20484 10231
rect 20444 10124 20496 10130
rect 20444 10066 20496 10072
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20456 8362 20484 9658
rect 20548 9654 20576 12922
rect 20640 11098 20668 13223
rect 20732 12986 20760 13631
rect 20812 13184 20864 13190
rect 20810 13152 20812 13161
rect 20864 13152 20866 13161
rect 20810 13087 20866 13096
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20824 12850 20852 13087
rect 20916 12986 20944 14447
rect 20994 13152 21050 13161
rect 20994 13087 21050 13096
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20812 12844 20864 12850
rect 20812 12786 20864 12792
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20732 12481 20760 12582
rect 20718 12472 20774 12481
rect 20718 12407 20774 12416
rect 20732 12374 20760 12407
rect 20720 12368 20772 12374
rect 20720 12310 20772 12316
rect 20718 11792 20774 11801
rect 20718 11727 20774 11736
rect 20732 11694 20760 11727
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20718 11384 20774 11393
rect 20718 11319 20720 11328
rect 20772 11319 20774 11328
rect 20720 11290 20772 11296
rect 20640 11070 20760 11098
rect 20628 11008 20680 11014
rect 20628 10950 20680 10956
rect 20640 10674 20668 10950
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 20640 9722 20668 9998
rect 20732 9874 20760 11070
rect 20824 10266 20852 12582
rect 20916 11762 20944 12718
rect 21008 12617 21036 13087
rect 21100 12646 21128 14470
rect 21192 12782 21220 14719
rect 21284 14618 21312 14844
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 21088 12640 21140 12646
rect 20994 12608 21050 12617
rect 21088 12582 21140 12588
rect 20994 12543 21050 12552
rect 21192 12442 21220 12718
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 21088 12164 21140 12170
rect 21088 12106 21140 12112
rect 20904 11756 20956 11762
rect 20956 11716 21036 11744
rect 20904 11698 20956 11704
rect 20902 11520 20958 11529
rect 20902 11455 20958 11464
rect 20916 11354 20944 11455
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20904 10532 20956 10538
rect 20904 10474 20956 10480
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 20732 9846 20852 9874
rect 20718 9752 20774 9761
rect 20628 9716 20680 9722
rect 20718 9687 20774 9696
rect 20628 9658 20680 9664
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20548 9353 20576 9454
rect 20534 9344 20590 9353
rect 20534 9279 20590 9288
rect 20640 8974 20668 9522
rect 20732 9178 20760 9687
rect 20824 9518 20852 9846
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20812 9376 20864 9382
rect 20916 9330 20944 10474
rect 20864 9324 20944 9330
rect 20812 9318 20944 9324
rect 20824 9302 20944 9318
rect 20916 9178 20944 9302
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20444 8356 20496 8362
rect 20444 8298 20496 8304
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20168 7210 20220 7216
rect 20272 7228 20392 7256
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20180 6322 20208 6598
rect 20168 6316 20220 6322
rect 20168 6258 20220 6264
rect 20272 5930 20300 7228
rect 20272 5902 20392 5930
rect 20258 5808 20314 5817
rect 20180 5752 20258 5760
rect 20180 5732 20260 5752
rect 20180 5234 20208 5732
rect 20312 5743 20314 5752
rect 20260 5714 20312 5720
rect 20168 5228 20220 5234
rect 20168 5170 20220 5176
rect 20168 5092 20220 5098
rect 20168 5034 20220 5040
rect 20180 5001 20208 5034
rect 20166 4992 20222 5001
rect 20166 4927 20222 4936
rect 20180 4282 20208 4927
rect 20258 4856 20314 4865
rect 20258 4791 20314 4800
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 20272 4078 20300 4791
rect 20364 4078 20392 5902
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19430 2680 19486 2689
rect 19622 2672 19918 2692
rect 20088 2689 20116 2994
rect 20074 2680 20130 2689
rect 19430 2615 19486 2624
rect 20074 2615 20130 2624
rect 20088 2514 20116 2615
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 19892 2304 19944 2310
rect 19892 2246 19944 2252
rect 19352 1550 19472 1578
rect 19338 1456 19394 1465
rect 19338 1391 19394 1400
rect 19352 480 19380 1391
rect 18144 264 18196 270
rect 18144 206 18196 212
rect 18234 0 18290 480
rect 18786 0 18842 480
rect 19338 0 19394 480
rect 19444 377 19472 1550
rect 19904 480 19932 2246
rect 19430 368 19486 377
rect 19430 303 19486 312
rect 19890 0 19946 480
rect 20180 105 20208 3946
rect 20364 3738 20392 4014
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20456 480 20484 7754
rect 20548 6633 20576 8570
rect 20534 6624 20590 6633
rect 20534 6559 20590 6568
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20548 5370 20576 6258
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20640 3777 20668 8774
rect 20732 8430 20760 9114
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20824 7546 20852 8978
rect 20902 8936 20958 8945
rect 21008 8906 21036 11716
rect 21100 11150 21128 12106
rect 21284 12050 21312 14554
rect 21376 14550 21404 17167
rect 21468 16522 21496 17614
rect 21456 16516 21508 16522
rect 21456 16458 21508 16464
rect 21454 16144 21510 16153
rect 21454 16079 21510 16088
rect 21468 14600 21496 16079
rect 21560 15706 21588 17847
rect 21652 17338 21680 18226
rect 21640 17332 21692 17338
rect 21640 17274 21692 17280
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21652 16946 21680 17138
rect 21744 17066 21772 18958
rect 21732 17060 21784 17066
rect 21732 17002 21784 17008
rect 21652 16918 21772 16946
rect 21548 15700 21600 15706
rect 21548 15642 21600 15648
rect 21640 15360 21692 15366
rect 21640 15302 21692 15308
rect 21468 14572 21588 14600
rect 21364 14544 21416 14550
rect 21364 14486 21416 14492
rect 21456 14476 21508 14482
rect 21456 14418 21508 14424
rect 21468 14074 21496 14418
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21376 12170 21404 13806
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21468 12481 21496 13330
rect 21560 12918 21588 14572
rect 21548 12912 21600 12918
rect 21548 12854 21600 12860
rect 21546 12608 21602 12617
rect 21546 12543 21602 12552
rect 21454 12472 21510 12481
rect 21454 12407 21510 12416
rect 21364 12164 21416 12170
rect 21364 12106 21416 12112
rect 21468 12050 21496 12407
rect 21192 12022 21312 12050
rect 21376 12022 21496 12050
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 21100 10538 21128 11086
rect 21088 10532 21140 10538
rect 21088 10474 21140 10480
rect 20902 8871 20958 8880
rect 20996 8900 21048 8906
rect 20916 8838 20944 8871
rect 20996 8842 21048 8848
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20916 7993 20944 8774
rect 20994 8664 21050 8673
rect 20994 8599 21050 8608
rect 21008 8498 21036 8599
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 21008 8090 21036 8434
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 20902 7984 20958 7993
rect 20902 7919 20958 7928
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 20732 7313 20760 7414
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20718 7304 20774 7313
rect 20718 7239 20774 7248
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20824 6905 20852 7142
rect 20916 7041 20944 7346
rect 20902 7032 20958 7041
rect 20902 6967 20958 6976
rect 20810 6896 20866 6905
rect 20810 6831 20866 6840
rect 20902 6760 20958 6769
rect 20902 6695 20904 6704
rect 20956 6695 20958 6704
rect 20904 6666 20956 6672
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 21008 6338 21036 6598
rect 21100 6458 21128 10474
rect 21192 9586 21220 12022
rect 21270 11928 21326 11937
rect 21270 11863 21326 11872
rect 21284 11762 21312 11863
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21270 11656 21326 11665
rect 21270 11591 21326 11600
rect 21284 11354 21312 11591
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21284 10266 21312 11290
rect 21376 11121 21404 12022
rect 21454 11928 21510 11937
rect 21454 11863 21510 11872
rect 21468 11762 21496 11863
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21362 11112 21418 11121
rect 21362 11047 21418 11056
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21376 9586 21404 11047
rect 21560 10674 21588 12543
rect 21652 11898 21680 15302
rect 21744 15042 21772 16918
rect 21836 15366 21864 22392
rect 21928 21418 21956 23598
rect 22008 23588 22060 23594
rect 22008 23530 22060 23536
rect 22020 23322 22048 23530
rect 22008 23316 22060 23322
rect 22008 23258 22060 23264
rect 22008 22976 22060 22982
rect 22008 22918 22060 22924
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22020 22234 22048 22918
rect 22008 22228 22060 22234
rect 22008 22170 22060 22176
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 21916 21412 21968 21418
rect 21916 21354 21968 21360
rect 21916 20800 21968 20806
rect 21916 20742 21968 20748
rect 21928 18902 21956 20742
rect 22020 20040 22048 21830
rect 22112 21049 22140 22918
rect 22204 21729 22232 25486
rect 22376 25356 22428 25362
rect 22376 25298 22428 25304
rect 22388 24614 22416 25298
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22284 23248 22336 23254
rect 22282 23216 22284 23225
rect 22336 23216 22338 23225
rect 22282 23151 22338 23160
rect 22388 23066 22416 24550
rect 22652 24268 22704 24274
rect 22652 24210 22704 24216
rect 22558 23760 22614 23769
rect 22558 23695 22614 23704
rect 22468 23520 22520 23526
rect 22468 23462 22520 23468
rect 22296 23038 22416 23066
rect 22190 21720 22246 21729
rect 22190 21655 22246 21664
rect 22098 21040 22154 21049
rect 22098 20975 22154 20984
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 22100 20052 22152 20058
rect 22020 20012 22100 20040
rect 22100 19994 22152 20000
rect 22008 19848 22060 19854
rect 22008 19790 22060 19796
rect 22020 18970 22048 19790
rect 22204 19718 22232 20538
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 21916 18896 21968 18902
rect 21916 18838 21968 18844
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 22020 17814 22048 18022
rect 22008 17808 22060 17814
rect 21914 17776 21970 17785
rect 22008 17750 22060 17756
rect 21914 17711 21916 17720
rect 21968 17711 21970 17720
rect 21916 17682 21968 17688
rect 21928 16794 21956 17682
rect 22112 16969 22140 19246
rect 22192 18148 22244 18154
rect 22192 18090 22244 18096
rect 22204 18057 22232 18090
rect 22190 18048 22246 18057
rect 22190 17983 22246 17992
rect 22190 17096 22246 17105
rect 22190 17031 22246 17040
rect 22098 16960 22154 16969
rect 22098 16895 22154 16904
rect 21916 16788 21968 16794
rect 21916 16730 21968 16736
rect 22006 16144 22062 16153
rect 22006 16079 22062 16088
rect 22100 16108 22152 16114
rect 22020 16046 22048 16079
rect 22100 16050 22152 16056
rect 22008 16040 22060 16046
rect 22008 15982 22060 15988
rect 22006 15736 22062 15745
rect 22112 15706 22140 16050
rect 22204 15706 22232 17031
rect 22006 15671 22062 15680
rect 22100 15700 22152 15706
rect 21916 15564 21968 15570
rect 21916 15506 21968 15512
rect 21824 15360 21876 15366
rect 21824 15302 21876 15308
rect 21928 15162 21956 15506
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 21744 15014 21956 15042
rect 21824 14884 21876 14890
rect 21824 14826 21876 14832
rect 21836 13530 21864 14826
rect 21824 13524 21876 13530
rect 21824 13466 21876 13472
rect 21730 12744 21786 12753
rect 21730 12679 21732 12688
rect 21784 12679 21786 12688
rect 21732 12650 21784 12656
rect 21836 12617 21864 13466
rect 21822 12608 21878 12617
rect 21822 12543 21878 12552
rect 21732 12300 21784 12306
rect 21732 12242 21784 12248
rect 21744 12073 21772 12242
rect 21824 12096 21876 12102
rect 21730 12064 21786 12073
rect 21824 12038 21876 12044
rect 21730 11999 21786 12008
rect 21836 11898 21864 12038
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21824 11892 21876 11898
rect 21824 11834 21876 11840
rect 21822 11248 21878 11257
rect 21822 11183 21878 11192
rect 21836 11082 21864 11183
rect 21824 11076 21876 11082
rect 21824 11018 21876 11024
rect 21822 10704 21878 10713
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21548 10668 21600 10674
rect 21822 10639 21878 10648
rect 21548 10610 21600 10616
rect 21468 10062 21496 10610
rect 21560 10266 21588 10610
rect 21640 10532 21692 10538
rect 21640 10474 21692 10480
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21546 10160 21602 10169
rect 21546 10095 21602 10104
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21454 9616 21510 9625
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 21364 9580 21416 9586
rect 21454 9551 21510 9560
rect 21364 9522 21416 9528
rect 21270 9208 21326 9217
rect 21270 9143 21326 9152
rect 21178 9072 21234 9081
rect 21178 9007 21234 9016
rect 21192 8673 21220 9007
rect 21178 8664 21234 8673
rect 21178 8599 21234 8608
rect 21284 8294 21312 9143
rect 21364 9104 21416 9110
rect 21362 9072 21364 9081
rect 21416 9072 21418 9081
rect 21362 9007 21418 9016
rect 21468 8974 21496 9551
rect 21560 9450 21588 10095
rect 21652 9994 21680 10474
rect 21730 10432 21786 10441
rect 21730 10367 21786 10376
rect 21640 9988 21692 9994
rect 21640 9930 21692 9936
rect 21638 9752 21694 9761
rect 21638 9687 21694 9696
rect 21652 9518 21680 9687
rect 21640 9512 21692 9518
rect 21640 9454 21692 9460
rect 21548 9444 21600 9450
rect 21548 9386 21600 9392
rect 21744 9042 21772 10367
rect 21836 10169 21864 10639
rect 21822 10160 21878 10169
rect 21822 10095 21878 10104
rect 21928 9874 21956 15014
rect 22020 14074 22048 15671
rect 22100 15642 22152 15648
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22112 15473 22140 15642
rect 22098 15464 22154 15473
rect 22098 15399 22154 15408
rect 22098 15328 22154 15337
rect 22098 15263 22154 15272
rect 22112 15162 22140 15263
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22204 14958 22232 15642
rect 22192 14952 22244 14958
rect 22192 14894 22244 14900
rect 22190 14648 22246 14657
rect 22190 14583 22246 14592
rect 22100 14544 22152 14550
rect 22100 14486 22152 14492
rect 22008 14068 22060 14074
rect 22008 14010 22060 14016
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 22020 13841 22048 13874
rect 22006 13832 22062 13841
rect 22112 13802 22140 14486
rect 22006 13767 22062 13776
rect 22100 13796 22152 13802
rect 22020 13530 22048 13767
rect 22100 13738 22152 13744
rect 22008 13524 22060 13530
rect 22008 13466 22060 13472
rect 22008 12912 22060 12918
rect 22008 12854 22060 12860
rect 22020 11744 22048 12854
rect 22100 12708 22152 12714
rect 22100 12650 22152 12656
rect 22112 12442 22140 12650
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22100 11756 22152 11762
rect 22020 11716 22100 11744
rect 22020 11354 22048 11716
rect 22100 11698 22152 11704
rect 22204 11506 22232 14583
rect 22296 13326 22324 23038
rect 22480 22234 22508 23462
rect 22468 22228 22520 22234
rect 22468 22170 22520 22176
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22388 20466 22416 21490
rect 22468 21344 22520 21350
rect 22468 21286 22520 21292
rect 22480 20806 22508 21286
rect 22468 20800 22520 20806
rect 22468 20742 22520 20748
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22376 19236 22428 19242
rect 22376 19178 22428 19184
rect 22388 19145 22416 19178
rect 22572 19156 22600 23695
rect 22664 23526 22692 24210
rect 22652 23520 22704 23526
rect 22650 23488 22652 23497
rect 22704 23488 22706 23497
rect 22650 23423 22706 23432
rect 22756 23322 22784 25910
rect 22652 23316 22704 23322
rect 22652 23258 22704 23264
rect 22744 23316 22796 23322
rect 22744 23258 22796 23264
rect 22664 20602 22692 23258
rect 22756 22710 22784 23258
rect 22836 23180 22888 23186
rect 22836 23122 22888 23128
rect 22848 23089 22876 23122
rect 22834 23080 22890 23089
rect 22834 23015 22890 23024
rect 22848 22778 22876 23015
rect 22836 22772 22888 22778
rect 22836 22714 22888 22720
rect 22744 22704 22796 22710
rect 22744 22646 22796 22652
rect 22836 22092 22888 22098
rect 22836 22034 22888 22040
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22756 21350 22784 21966
rect 22744 21344 22796 21350
rect 22744 21286 22796 21292
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 22756 20097 22784 21286
rect 22742 20088 22798 20097
rect 22742 20023 22798 20032
rect 22756 19417 22784 20023
rect 22742 19408 22798 19417
rect 22652 19372 22704 19378
rect 22742 19343 22798 19352
rect 22652 19314 22704 19320
rect 22374 19136 22430 19145
rect 22374 19071 22430 19080
rect 22480 19128 22600 19156
rect 22480 18850 22508 19128
rect 22664 18970 22692 19314
rect 22652 18964 22704 18970
rect 22652 18906 22704 18912
rect 22388 18822 22508 18850
rect 22560 18896 22612 18902
rect 22560 18838 22612 18844
rect 22388 18086 22416 18822
rect 22466 18728 22522 18737
rect 22466 18663 22522 18672
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22480 17134 22508 18663
rect 22572 17882 22600 18838
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22664 17814 22692 18906
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22756 18426 22784 18566
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22652 17808 22704 17814
rect 22652 17750 22704 17756
rect 22664 17338 22692 17750
rect 22756 17746 22784 18362
rect 22744 17740 22796 17746
rect 22744 17682 22796 17688
rect 22756 17338 22784 17682
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 22468 17128 22520 17134
rect 22468 17070 22520 17076
rect 22480 16794 22508 17070
rect 22560 17060 22612 17066
rect 22560 17002 22612 17008
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22468 16244 22520 16250
rect 22468 16186 22520 16192
rect 22376 15564 22428 15570
rect 22376 15506 22428 15512
rect 22388 15094 22416 15506
rect 22480 15502 22508 16186
rect 22468 15496 22520 15502
rect 22468 15438 22520 15444
rect 22572 15162 22600 17002
rect 22652 16992 22704 16998
rect 22652 16934 22704 16940
rect 22664 16697 22692 16934
rect 22650 16688 22706 16697
rect 22756 16658 22784 17274
rect 22650 16623 22706 16632
rect 22744 16652 22796 16658
rect 22744 16594 22796 16600
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22664 16289 22692 16390
rect 22650 16280 22706 16289
rect 22756 16250 22784 16594
rect 22650 16215 22706 16224
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22376 15088 22428 15094
rect 22376 15030 22428 15036
rect 22388 14618 22416 15030
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 22376 14000 22428 14006
rect 22376 13942 22428 13948
rect 22388 13841 22416 13942
rect 22374 13832 22430 13841
rect 22374 13767 22430 13776
rect 22284 13320 22336 13326
rect 22284 13262 22336 13268
rect 22284 13184 22336 13190
rect 22282 13152 22284 13161
rect 22336 13152 22338 13161
rect 22282 13087 22338 13096
rect 22376 12912 22428 12918
rect 22374 12880 22376 12889
rect 22428 12880 22430 12889
rect 22374 12815 22430 12824
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 22296 11898 22324 12174
rect 22374 11928 22430 11937
rect 22284 11892 22336 11898
rect 22374 11863 22430 11872
rect 22284 11834 22336 11840
rect 22388 11762 22416 11863
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22204 11478 22324 11506
rect 22190 11384 22246 11393
rect 22008 11348 22060 11354
rect 22190 11319 22246 11328
rect 22008 11290 22060 11296
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22020 10674 22048 11086
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 22020 10266 22048 10610
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 21928 9846 22048 9874
rect 21822 9616 21878 9625
rect 21822 9551 21878 9560
rect 21916 9580 21968 9586
rect 21732 9036 21784 9042
rect 21732 8978 21784 8984
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21376 8838 21404 8910
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 21272 8288 21324 8294
rect 21178 8256 21234 8265
rect 21272 8230 21324 8236
rect 21178 8191 21234 8200
rect 21192 7546 21220 8191
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21284 7002 21312 8230
rect 21376 7585 21404 8774
rect 21468 8634 21496 8910
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 21732 8424 21784 8430
rect 21836 8401 21864 9551
rect 21916 9522 21968 9528
rect 21928 9178 21956 9522
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 21916 8900 21968 8906
rect 21916 8842 21968 8848
rect 21732 8366 21784 8372
rect 21822 8392 21878 8401
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21362 7576 21418 7585
rect 21362 7511 21418 7520
rect 21560 7449 21588 7686
rect 21546 7440 21602 7449
rect 21652 7410 21680 8230
rect 21744 7970 21772 8366
rect 21822 8327 21878 8336
rect 21928 8022 21956 8842
rect 21916 8016 21968 8022
rect 21744 7942 21864 7970
rect 21916 7958 21968 7964
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21546 7375 21602 7384
rect 21640 7404 21692 7410
rect 21560 7342 21588 7375
rect 21640 7346 21692 7352
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21652 7177 21680 7346
rect 21744 7206 21772 7822
rect 21836 7313 21864 7942
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 21822 7304 21878 7313
rect 21822 7239 21878 7248
rect 21732 7200 21784 7206
rect 21638 7168 21694 7177
rect 21732 7142 21784 7148
rect 21638 7103 21694 7112
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21180 6792 21232 6798
rect 21178 6760 21180 6769
rect 21232 6760 21234 6769
rect 21178 6695 21234 6704
rect 21178 6488 21234 6497
rect 21088 6452 21140 6458
rect 21178 6423 21234 6432
rect 21088 6394 21140 6400
rect 21008 6322 21128 6338
rect 21008 6316 21140 6322
rect 21008 6310 21088 6316
rect 21088 6258 21140 6264
rect 20810 6080 20866 6089
rect 20810 6015 20866 6024
rect 20718 5128 20774 5137
rect 20718 5063 20774 5072
rect 20732 4826 20760 5063
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20732 4049 20760 4558
rect 20718 4040 20774 4049
rect 20718 3975 20774 3984
rect 20626 3768 20682 3777
rect 20626 3703 20682 3712
rect 20732 3194 20760 3975
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 20824 2990 20852 6015
rect 20994 5400 21050 5409
rect 20994 5335 20996 5344
rect 21048 5335 21050 5344
rect 20996 5306 21048 5312
rect 20996 4072 21048 4078
rect 20996 4014 21048 4020
rect 21008 3942 21036 4014
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 21008 3505 21036 3878
rect 20994 3496 21050 3505
rect 20994 3431 21050 3440
rect 20994 3224 21050 3233
rect 21100 3210 21128 6258
rect 21192 6118 21220 6423
rect 21284 6390 21312 6938
rect 21454 6896 21510 6905
rect 21454 6831 21510 6840
rect 21364 6792 21416 6798
rect 21468 6780 21496 6831
rect 21416 6752 21496 6780
rect 21364 6734 21416 6740
rect 21272 6384 21324 6390
rect 21272 6326 21324 6332
rect 21270 6216 21326 6225
rect 21270 6151 21326 6160
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 21284 5953 21312 6151
rect 21270 5944 21326 5953
rect 21270 5879 21326 5888
rect 21364 5908 21416 5914
rect 21284 5846 21312 5879
rect 21364 5850 21416 5856
rect 21272 5840 21324 5846
rect 21376 5817 21404 5850
rect 21272 5782 21324 5788
rect 21362 5808 21418 5817
rect 21362 5743 21418 5752
rect 21468 5574 21496 6752
rect 21546 6352 21602 6361
rect 21546 6287 21602 6296
rect 21560 6254 21588 6287
rect 21548 6248 21600 6254
rect 21744 6225 21772 7142
rect 21548 6190 21600 6196
rect 21730 6216 21786 6225
rect 21560 5914 21588 6190
rect 21730 6151 21786 6160
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 21822 5672 21878 5681
rect 21548 5636 21600 5642
rect 21548 5578 21600 5584
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21468 5098 21496 5510
rect 21560 5166 21588 5578
rect 21640 5228 21692 5234
rect 21640 5170 21692 5176
rect 21548 5160 21600 5166
rect 21652 5137 21680 5170
rect 21548 5102 21600 5108
rect 21638 5128 21694 5137
rect 21456 5092 21508 5098
rect 21638 5063 21694 5072
rect 21456 5034 21508 5040
rect 21180 5024 21232 5030
rect 21180 4966 21232 4972
rect 21192 4457 21220 4966
rect 21744 4826 21772 5646
rect 21822 5607 21878 5616
rect 21836 5574 21864 5607
rect 21824 5568 21876 5574
rect 21824 5510 21876 5516
rect 21928 5386 21956 7686
rect 22020 7206 22048 9846
rect 22112 9042 22140 10746
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 22204 8537 22232 11319
rect 22296 10713 22324 11478
rect 22388 11286 22416 11698
rect 22480 11354 22508 15098
rect 22572 14056 22600 15098
rect 22756 15094 22784 16186
rect 22848 15366 22876 22034
rect 22940 21078 22968 26046
rect 23032 25498 23060 27520
rect 23296 26512 23348 26518
rect 23296 26454 23348 26460
rect 23202 25936 23258 25945
rect 23202 25871 23258 25880
rect 23020 25492 23072 25498
rect 23020 25434 23072 25440
rect 23216 25294 23244 25871
rect 23204 25288 23256 25294
rect 23110 25256 23166 25265
rect 23204 25230 23256 25236
rect 23110 25191 23166 25200
rect 23018 24168 23074 24177
rect 23018 24103 23074 24112
rect 23032 22234 23060 24103
rect 23020 22228 23072 22234
rect 23020 22170 23072 22176
rect 23032 21690 23060 22170
rect 23020 21684 23072 21690
rect 23020 21626 23072 21632
rect 23032 21486 23060 21626
rect 23020 21480 23072 21486
rect 23020 21422 23072 21428
rect 22928 21072 22980 21078
rect 22928 21014 22980 21020
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 22836 15360 22888 15366
rect 22836 15302 22888 15308
rect 22744 15088 22796 15094
rect 22744 15030 22796 15036
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22664 14521 22692 14758
rect 22650 14512 22706 14521
rect 22650 14447 22706 14456
rect 22756 14362 22784 15030
rect 22664 14334 22784 14362
rect 22664 14278 22692 14334
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22756 14074 22784 14334
rect 22744 14068 22796 14074
rect 22572 14028 22692 14056
rect 22664 13734 22692 14028
rect 22744 14010 22796 14016
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 22756 13546 22784 14010
rect 22664 13518 22784 13546
rect 22664 13462 22692 13518
rect 22652 13456 22704 13462
rect 22652 13398 22704 13404
rect 22744 13388 22796 13394
rect 22744 13330 22796 13336
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22376 11280 22428 11286
rect 22376 11222 22428 11228
rect 22572 10810 22600 13262
rect 22756 13025 22784 13330
rect 22742 13016 22798 13025
rect 22742 12951 22744 12960
rect 22796 12951 22798 12960
rect 22744 12922 22796 12928
rect 22756 12891 22784 12922
rect 22848 12850 22876 15302
rect 22836 12844 22888 12850
rect 22836 12786 22888 12792
rect 22650 12744 22706 12753
rect 22940 12730 22968 20538
rect 23020 20392 23072 20398
rect 23020 20334 23072 20340
rect 23032 18834 23060 20334
rect 23124 19990 23152 25191
rect 23204 23112 23256 23118
rect 23204 23054 23256 23060
rect 23216 22438 23244 23054
rect 23204 22432 23256 22438
rect 23204 22374 23256 22380
rect 23308 22386 23336 26454
rect 23480 25696 23532 25702
rect 23480 25638 23532 25644
rect 23492 23066 23520 25638
rect 23584 24857 23612 27520
rect 23768 26858 23796 27639
rect 24122 27520 24178 28000
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25870 27520 25926 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 23756 26852 23808 26858
rect 23756 26794 23808 26800
rect 23754 26616 23810 26625
rect 23754 26551 23810 26560
rect 23768 26314 23796 26551
rect 23756 26308 23808 26314
rect 23756 26250 23808 26256
rect 23756 25900 23808 25906
rect 23756 25842 23808 25848
rect 23570 24848 23626 24857
rect 23570 24783 23626 24792
rect 23572 24608 23624 24614
rect 23572 24550 23624 24556
rect 23400 23038 23520 23066
rect 23400 22556 23428 23038
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23492 22681 23520 22918
rect 23478 22672 23534 22681
rect 23478 22607 23534 22616
rect 23400 22528 23520 22556
rect 23112 19984 23164 19990
rect 23112 19926 23164 19932
rect 23112 19712 23164 19718
rect 23112 19654 23164 19660
rect 23124 19446 23152 19654
rect 23112 19440 23164 19446
rect 23112 19382 23164 19388
rect 23112 19304 23164 19310
rect 23112 19246 23164 19252
rect 23124 18902 23152 19246
rect 23112 18896 23164 18902
rect 23112 18838 23164 18844
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 23018 18728 23074 18737
rect 23018 18663 23074 18672
rect 23032 18426 23060 18663
rect 23020 18420 23072 18426
rect 23020 18362 23072 18368
rect 23032 18222 23060 18362
rect 23020 18216 23072 18222
rect 23020 18158 23072 18164
rect 23112 17876 23164 17882
rect 23112 17818 23164 17824
rect 23124 16998 23152 17818
rect 23112 16992 23164 16998
rect 23018 16960 23074 16969
rect 23112 16934 23164 16940
rect 23018 16895 23074 16904
rect 22650 12679 22706 12688
rect 22848 12702 22968 12730
rect 22664 12374 22692 12679
rect 22652 12368 22704 12374
rect 22652 12310 22704 12316
rect 22744 11212 22796 11218
rect 22744 11154 22796 11160
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22282 10704 22338 10713
rect 22282 10639 22338 10648
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22296 10130 22324 10406
rect 22284 10124 22336 10130
rect 22284 10066 22336 10072
rect 22296 9722 22324 10066
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22190 8528 22246 8537
rect 22190 8463 22192 8472
rect 22244 8463 22246 8472
rect 22192 8434 22244 8440
rect 22204 8403 22232 8434
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 22112 6848 22140 7142
rect 22020 6820 22140 6848
rect 22020 6730 22048 6820
rect 22296 6746 22324 8774
rect 22388 8072 22416 10610
rect 22560 10600 22612 10606
rect 22466 10568 22522 10577
rect 22560 10542 22612 10548
rect 22466 10503 22522 10512
rect 22480 10266 22508 10503
rect 22468 10260 22520 10266
rect 22468 10202 22520 10208
rect 22388 8044 22508 8072
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22388 7750 22416 7890
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22388 7002 22416 7686
rect 22376 6996 22428 7002
rect 22376 6938 22428 6944
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 22008 6724 22060 6730
rect 22008 6666 22060 6672
rect 22204 6718 22324 6746
rect 22020 6089 22048 6666
rect 22006 6080 22062 6089
rect 22006 6015 22062 6024
rect 22204 5930 22232 6718
rect 22284 6656 22336 6662
rect 22282 6624 22284 6633
rect 22336 6624 22338 6633
rect 22282 6559 22338 6568
rect 22388 6304 22416 6802
rect 22020 5902 22232 5930
rect 22296 6276 22416 6304
rect 22020 5642 22048 5902
rect 22008 5636 22060 5642
rect 22008 5578 22060 5584
rect 22098 5400 22154 5409
rect 21928 5358 22098 5386
rect 22098 5335 22154 5344
rect 22192 5296 22244 5302
rect 22192 5238 22244 5244
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 21270 4720 21326 4729
rect 21270 4655 21272 4664
rect 21324 4655 21326 4664
rect 21272 4626 21324 4632
rect 21178 4448 21234 4457
rect 21178 4383 21234 4392
rect 21284 4026 21312 4626
rect 21916 4480 21968 4486
rect 21916 4422 21968 4428
rect 21732 4140 21784 4146
rect 21732 4082 21784 4088
rect 21284 3998 21496 4026
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 21362 3904 21418 3913
rect 21192 3233 21220 3878
rect 21362 3839 21418 3848
rect 21376 3738 21404 3839
rect 21364 3732 21416 3738
rect 21364 3674 21416 3680
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 21284 3369 21312 3538
rect 21270 3360 21326 3369
rect 21270 3295 21326 3304
rect 21050 3182 21128 3210
rect 21178 3224 21234 3233
rect 20994 3159 21050 3168
rect 21178 3159 21234 3168
rect 21284 2990 21312 3295
rect 20812 2984 20864 2990
rect 20718 2952 20774 2961
rect 21272 2984 21324 2990
rect 20812 2926 20864 2932
rect 21086 2952 21142 2961
rect 20718 2887 20720 2896
rect 20772 2887 20774 2896
rect 20996 2916 21048 2922
rect 20720 2858 20772 2864
rect 21272 2926 21324 2932
rect 21086 2887 21142 2896
rect 20996 2858 21048 2864
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 20534 2408 20590 2417
rect 20534 2343 20536 2352
rect 20588 2343 20590 2352
rect 20536 2314 20588 2320
rect 20916 2310 20944 2518
rect 20904 2304 20956 2310
rect 20902 2272 20904 2281
rect 20956 2272 20958 2281
rect 20902 2207 20958 2216
rect 21008 2009 21036 2858
rect 20994 2000 21050 2009
rect 20994 1935 21050 1944
rect 21100 1034 21128 2887
rect 21376 2854 21404 3674
rect 21468 3670 21496 3998
rect 21546 3768 21602 3777
rect 21546 3703 21602 3712
rect 21456 3664 21508 3670
rect 21456 3606 21508 3612
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21008 1006 21128 1034
rect 21008 480 21036 1006
rect 21560 480 21588 3703
rect 21744 3534 21772 4082
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21744 3058 21772 3470
rect 21732 3052 21784 3058
rect 21732 2994 21784 3000
rect 21744 2446 21772 2994
rect 21928 2553 21956 4422
rect 22112 4010 22140 5170
rect 22204 5137 22232 5238
rect 22190 5128 22246 5137
rect 22190 5063 22246 5072
rect 22100 4004 22152 4010
rect 22100 3946 22152 3952
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 22008 3528 22060 3534
rect 22008 3470 22060 3476
rect 22020 3194 22048 3470
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22112 2666 22140 3538
rect 22020 2650 22140 2666
rect 22008 2644 22140 2650
rect 22060 2638 22140 2644
rect 22008 2586 22060 2592
rect 21914 2544 21970 2553
rect 21914 2479 21970 2488
rect 21732 2440 21784 2446
rect 21732 2382 21784 2388
rect 22204 1442 22232 3946
rect 22296 3194 22324 6276
rect 22480 6236 22508 8044
rect 22572 7410 22600 10542
rect 22664 10062 22692 10746
rect 22756 10674 22784 11154
rect 22744 10668 22796 10674
rect 22744 10610 22796 10616
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22664 9722 22692 9998
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22652 8832 22704 8838
rect 22652 8774 22704 8780
rect 22560 7404 22612 7410
rect 22560 7346 22612 7352
rect 22664 6905 22692 8774
rect 22848 8634 22876 12702
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 22940 10606 22968 11086
rect 22928 10600 22980 10606
rect 22928 10542 22980 10548
rect 22928 10192 22980 10198
rect 22926 10160 22928 10169
rect 22980 10160 22982 10169
rect 22926 10095 22982 10104
rect 22928 9648 22980 9654
rect 22926 9616 22928 9625
rect 22980 9616 22982 9625
rect 22926 9551 22982 9560
rect 23032 9382 23060 16895
rect 23124 12782 23152 16934
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 23110 12608 23166 12617
rect 23110 12543 23166 12552
rect 23124 11014 23152 12543
rect 23216 11150 23244 22374
rect 23308 22358 23428 22386
rect 23296 22024 23348 22030
rect 23296 21966 23348 21972
rect 23308 21622 23336 21966
rect 23296 21616 23348 21622
rect 23296 21558 23348 21564
rect 23400 21298 23428 22358
rect 23308 21270 23428 21298
rect 23308 17882 23336 21270
rect 23386 19680 23442 19689
rect 23386 19615 23442 19624
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 23296 16720 23348 16726
rect 23296 16662 23348 16668
rect 23308 16250 23336 16662
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 23308 12918 23336 15846
rect 23400 14657 23428 19615
rect 23492 17490 23520 22528
rect 23584 18873 23612 24550
rect 23662 23760 23718 23769
rect 23662 23695 23718 23704
rect 23676 23497 23704 23695
rect 23662 23488 23718 23497
rect 23662 23423 23718 23432
rect 23662 22944 23718 22953
rect 23662 22879 23718 22888
rect 23676 22574 23704 22879
rect 23664 22568 23716 22574
rect 23664 22510 23716 22516
rect 23768 22273 23796 25842
rect 24030 24712 24086 24721
rect 24030 24647 24086 24656
rect 24044 24614 24072 24647
rect 24032 24608 24084 24614
rect 24032 24550 24084 24556
rect 24136 24410 24164 27520
rect 24780 27282 24808 27520
rect 24596 27254 24808 27282
rect 24596 25770 24624 27254
rect 24766 27160 24822 27169
rect 24766 27095 24822 27104
rect 24780 26722 24808 27095
rect 24768 26716 24820 26722
rect 24768 26658 24820 26664
rect 25044 26172 25096 26178
rect 25044 26114 25096 26120
rect 24584 25764 24636 25770
rect 24584 25706 24636 25712
rect 24766 25392 24822 25401
rect 24216 25356 24268 25362
rect 24766 25327 24822 25336
rect 24216 25298 24268 25304
rect 24228 24596 24256 25298
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24780 24886 24808 25327
rect 24768 24880 24820 24886
rect 24768 24822 24820 24828
rect 24400 24608 24452 24614
rect 24228 24568 24400 24596
rect 24400 24550 24452 24556
rect 24124 24404 24176 24410
rect 24124 24346 24176 24352
rect 24412 24313 24440 24550
rect 24674 24440 24730 24449
rect 24674 24375 24676 24384
rect 24728 24375 24730 24384
rect 24676 24346 24728 24352
rect 24398 24304 24454 24313
rect 24124 24268 24176 24274
rect 24398 24239 24454 24248
rect 24124 24210 24176 24216
rect 23846 23760 23902 23769
rect 24136 23730 24164 24210
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24766 23896 24822 23905
rect 24766 23831 24768 23840
rect 24820 23831 24822 23840
rect 24768 23802 24820 23808
rect 23846 23695 23902 23704
rect 24124 23724 24176 23730
rect 23860 22778 23888 23695
rect 24124 23666 24176 23672
rect 24032 23520 24084 23526
rect 24032 23462 24084 23468
rect 23848 22772 23900 22778
rect 23848 22714 23900 22720
rect 23754 22264 23810 22273
rect 23754 22199 23810 22208
rect 24044 22098 24072 23462
rect 24032 22092 24084 22098
rect 24032 22034 24084 22040
rect 24136 22030 24164 23666
rect 24766 23488 24822 23497
rect 24766 23423 24822 23432
rect 24780 23322 24808 23423
rect 24768 23316 24820 23322
rect 24768 23258 24820 23264
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22506 24716 23122
rect 24676 22500 24728 22506
rect 24676 22442 24728 22448
rect 24124 22024 24176 22030
rect 23846 21992 23902 22001
rect 24124 21966 24176 21972
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 23846 21927 23902 21936
rect 23940 21956 23992 21962
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23768 21622 23796 21830
rect 23756 21616 23808 21622
rect 23756 21558 23808 21564
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23676 20262 23704 20742
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23570 18864 23626 18873
rect 23570 18799 23626 18808
rect 23570 18728 23626 18737
rect 23570 18663 23626 18672
rect 23584 18358 23612 18663
rect 23676 18601 23704 20198
rect 23662 18592 23718 18601
rect 23662 18527 23718 18536
rect 23572 18352 23624 18358
rect 23572 18294 23624 18300
rect 23662 17640 23718 17649
rect 23662 17575 23718 17584
rect 23492 17462 23612 17490
rect 23478 17368 23534 17377
rect 23478 17303 23480 17312
rect 23532 17303 23534 17312
rect 23480 17274 23532 17280
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23492 14958 23520 15302
rect 23480 14952 23532 14958
rect 23478 14920 23480 14929
rect 23532 14920 23534 14929
rect 23478 14855 23534 14864
rect 23386 14648 23442 14657
rect 23386 14583 23442 14592
rect 23480 14612 23532 14618
rect 23480 14554 23532 14560
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 23400 13954 23428 14418
rect 23492 14074 23520 14554
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23400 13926 23520 13954
rect 23386 13560 23442 13569
rect 23386 13495 23442 13504
rect 23400 13326 23428 13495
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23400 12986 23428 13262
rect 23492 13258 23520 13926
rect 23480 13252 23532 13258
rect 23480 13194 23532 13200
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23296 12912 23348 12918
rect 23296 12854 23348 12860
rect 23296 12776 23348 12782
rect 23296 12718 23348 12724
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 23112 11008 23164 11014
rect 23112 10950 23164 10956
rect 23216 10810 23244 11086
rect 23204 10804 23256 10810
rect 23204 10746 23256 10752
rect 23308 10690 23336 12718
rect 23492 12714 23520 13194
rect 23480 12708 23532 12714
rect 23480 12650 23532 12656
rect 23386 12472 23442 12481
rect 23386 12407 23388 12416
rect 23440 12407 23442 12416
rect 23388 12378 23440 12384
rect 23492 12374 23520 12650
rect 23584 12617 23612 17462
rect 23676 17338 23704 17575
rect 23664 17332 23716 17338
rect 23664 17274 23716 17280
rect 23664 17128 23716 17134
rect 23664 17070 23716 17076
rect 23676 16250 23704 17070
rect 23768 17066 23796 21286
rect 23756 17060 23808 17066
rect 23756 17002 23808 17008
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23664 16244 23716 16250
rect 23664 16186 23716 16192
rect 23664 14816 23716 14822
rect 23664 14758 23716 14764
rect 23570 12608 23626 12617
rect 23570 12543 23626 12552
rect 23480 12368 23532 12374
rect 23480 12310 23532 12316
rect 23492 12238 23520 12310
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23570 12200 23626 12209
rect 23570 12135 23626 12144
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 23124 10662 23336 10690
rect 23020 9376 23072 9382
rect 23020 9318 23072 9324
rect 23020 9036 23072 9042
rect 23020 8978 23072 8984
rect 22928 8832 22980 8838
rect 22928 8774 22980 8780
rect 22836 8628 22888 8634
rect 22836 8570 22888 8576
rect 22742 8528 22798 8537
rect 22742 8463 22798 8472
rect 22756 8294 22784 8463
rect 22744 8288 22796 8294
rect 22744 8230 22796 8236
rect 22848 8090 22876 8570
rect 22940 8401 22968 8774
rect 23032 8634 23060 8978
rect 23020 8628 23072 8634
rect 23020 8570 23072 8576
rect 22926 8392 22982 8401
rect 22926 8327 22982 8336
rect 22836 8084 22888 8090
rect 22888 8044 22968 8072
rect 22836 8026 22888 8032
rect 22834 7984 22890 7993
rect 22744 7948 22796 7954
rect 22834 7919 22890 7928
rect 22744 7890 22796 7896
rect 22756 7274 22784 7890
rect 22744 7268 22796 7274
rect 22744 7210 22796 7216
rect 22848 7002 22876 7919
rect 22940 7546 22968 8044
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 23032 7206 23060 7822
rect 23020 7200 23072 7206
rect 23020 7142 23072 7148
rect 22926 7032 22982 7041
rect 22836 6996 22888 7002
rect 22926 6967 22982 6976
rect 22836 6938 22888 6944
rect 22650 6896 22706 6905
rect 22650 6831 22706 6840
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22572 6458 22600 6734
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22388 6208 22508 6236
rect 22560 6248 22612 6254
rect 22388 4162 22416 6208
rect 22560 6190 22612 6196
rect 22468 6112 22520 6118
rect 22468 6054 22520 6060
rect 22480 5914 22508 6054
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 22466 4584 22522 4593
rect 22572 4570 22600 6190
rect 22756 5778 22784 6802
rect 22848 6458 22876 6938
rect 22836 6452 22888 6458
rect 22836 6394 22888 6400
rect 22940 5914 22968 6967
rect 22928 5908 22980 5914
rect 22928 5850 22980 5856
rect 22744 5772 22796 5778
rect 22744 5714 22796 5720
rect 22756 5370 22784 5714
rect 22940 5370 22968 5850
rect 23020 5704 23072 5710
rect 23020 5646 23072 5652
rect 22744 5364 22796 5370
rect 22744 5306 22796 5312
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 23032 5273 23060 5646
rect 23018 5264 23074 5273
rect 23018 5199 23074 5208
rect 22652 5092 22704 5098
rect 22652 5034 22704 5040
rect 22664 4593 22692 5034
rect 23032 4826 23060 5199
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 23124 4758 23152 10662
rect 23296 10056 23348 10062
rect 23294 10024 23296 10033
rect 23348 10024 23350 10033
rect 23204 9988 23256 9994
rect 23400 10010 23428 11494
rect 23492 11150 23520 11698
rect 23584 11286 23612 12135
rect 23572 11280 23624 11286
rect 23572 11222 23624 11228
rect 23480 11144 23532 11150
rect 23478 11112 23480 11121
rect 23532 11112 23534 11121
rect 23478 11047 23534 11056
rect 23480 11008 23532 11014
rect 23480 10950 23532 10956
rect 23492 10169 23520 10950
rect 23570 10704 23626 10713
rect 23570 10639 23626 10648
rect 23478 10160 23534 10169
rect 23478 10095 23534 10104
rect 23584 10033 23612 10639
rect 23676 10130 23704 14758
rect 23768 12442 23796 16594
rect 23860 13190 23888 21927
rect 23940 21898 23992 21904
rect 23952 21729 23980 21898
rect 24032 21888 24084 21894
rect 24030 21856 24032 21865
rect 24124 21888 24176 21894
rect 24084 21856 24086 21865
rect 24124 21830 24176 21836
rect 24030 21791 24086 21800
rect 23938 21720 23994 21729
rect 23938 21655 23994 21664
rect 23938 21584 23994 21593
rect 24044 21554 24072 21791
rect 23938 21519 23994 21528
rect 24032 21548 24084 21554
rect 23952 21418 23980 21519
rect 24032 21490 24084 21496
rect 23940 21412 23992 21418
rect 23940 21354 23992 21360
rect 23952 21010 23980 21354
rect 23940 21004 23992 21010
rect 23940 20946 23992 20952
rect 24136 20890 24164 21830
rect 24228 21321 24256 21966
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21672 24716 22442
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24320 21644 24716 21672
rect 24214 21312 24270 21321
rect 24214 21247 24270 21256
rect 24320 21162 24348 21644
rect 24400 21548 24452 21554
rect 24400 21490 24452 21496
rect 23952 20862 24164 20890
rect 24228 21134 24348 21162
rect 23952 16658 23980 20862
rect 24032 20800 24084 20806
rect 24030 20768 24032 20777
rect 24124 20800 24176 20806
rect 24084 20768 24086 20777
rect 24124 20742 24176 20748
rect 24030 20703 24086 20712
rect 24032 20256 24084 20262
rect 24032 20198 24084 20204
rect 24044 19854 24072 20198
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 24044 19446 24072 19790
rect 24032 19440 24084 19446
rect 24032 19382 24084 19388
rect 24136 19310 24164 20742
rect 24124 19304 24176 19310
rect 24124 19246 24176 19252
rect 24228 19258 24256 21134
rect 24412 20874 24440 21490
rect 24584 21344 24636 21350
rect 24582 21312 24584 21321
rect 24636 21312 24638 21321
rect 24582 21247 24638 21256
rect 24780 21146 24808 22374
rect 24950 22128 25006 22137
rect 24860 22092 24912 22098
rect 24950 22063 25006 22072
rect 24860 22034 24912 22040
rect 24872 21690 24900 22034
rect 24860 21684 24912 21690
rect 24860 21626 24912 21632
rect 24768 21140 24820 21146
rect 24820 21100 24900 21128
rect 24768 21082 24820 21088
rect 24676 21072 24728 21078
rect 24676 21014 24728 21020
rect 24400 20868 24452 20874
rect 24400 20810 24452 20816
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20058 24716 21014
rect 24768 20800 24820 20806
rect 24768 20742 24820 20748
rect 24676 20052 24728 20058
rect 24676 19994 24728 20000
rect 24584 19984 24636 19990
rect 24636 19932 24716 19938
rect 24584 19926 24716 19932
rect 24596 19910 24716 19926
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24490 19408 24546 19417
rect 24490 19343 24546 19352
rect 24136 18970 24164 19246
rect 24228 19230 24348 19258
rect 24216 19168 24268 19174
rect 24216 19110 24268 19116
rect 24124 18964 24176 18970
rect 24124 18906 24176 18912
rect 24124 18828 24176 18834
rect 24124 18770 24176 18776
rect 24030 18592 24086 18601
rect 24030 18527 24086 18536
rect 24044 18290 24072 18527
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 24136 18222 24164 18770
rect 24228 18630 24256 19110
rect 24320 18834 24348 19230
rect 24308 18828 24360 18834
rect 24308 18770 24360 18776
rect 24504 18737 24532 19343
rect 24490 18728 24546 18737
rect 24490 18663 24546 18672
rect 24216 18624 24268 18630
rect 24216 18566 24268 18572
rect 24228 18426 24256 18566
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24216 18420 24268 18426
rect 24216 18362 24268 18368
rect 24400 18352 24452 18358
rect 24400 18294 24452 18300
rect 24124 18216 24176 18222
rect 24030 18184 24086 18193
rect 24124 18158 24176 18164
rect 24030 18119 24086 18128
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 23940 16516 23992 16522
rect 23940 16458 23992 16464
rect 23952 15978 23980 16458
rect 24044 16114 24072 18119
rect 24124 18080 24176 18086
rect 24124 18022 24176 18028
rect 24032 16108 24084 16114
rect 24032 16050 24084 16056
rect 23940 15972 23992 15978
rect 23940 15914 23992 15920
rect 23952 15337 23980 15914
rect 24032 15904 24084 15910
rect 24032 15846 24084 15852
rect 24044 15745 24072 15846
rect 24030 15736 24086 15745
rect 24030 15671 24032 15680
rect 24084 15671 24086 15680
rect 24032 15642 24084 15648
rect 24044 15611 24072 15642
rect 24136 15450 24164 18022
rect 24412 17882 24440 18294
rect 24688 18154 24716 19910
rect 24780 18193 24808 20742
rect 24872 20058 24900 21100
rect 24860 20052 24912 20058
rect 24860 19994 24912 20000
rect 24964 19938 24992 22063
rect 24872 19910 24992 19938
rect 24872 18222 24900 19910
rect 24952 19712 25004 19718
rect 24952 19654 25004 19660
rect 24964 19514 24992 19654
rect 24952 19508 25004 19514
rect 24952 19450 25004 19456
rect 24952 18828 25004 18834
rect 24952 18770 25004 18776
rect 24964 18358 24992 18770
rect 24952 18352 25004 18358
rect 24950 18320 24952 18329
rect 25004 18320 25006 18329
rect 24950 18255 25006 18264
rect 24860 18216 24912 18222
rect 24766 18184 24822 18193
rect 24676 18148 24728 18154
rect 24860 18158 24912 18164
rect 24766 18119 24822 18128
rect 24676 18090 24728 18096
rect 24216 17876 24268 17882
rect 24216 17818 24268 17824
rect 24400 17876 24452 17882
rect 24400 17818 24452 17824
rect 24228 16726 24256 17818
rect 24766 17776 24822 17785
rect 25056 17762 25084 26114
rect 25226 24848 25282 24857
rect 25226 24783 25282 24792
rect 25240 23361 25268 24783
rect 25332 23769 25360 27520
rect 25778 26208 25834 26217
rect 25778 26143 25834 26152
rect 25792 24596 25820 26143
rect 25884 24721 25912 27520
rect 26146 25800 26202 25809
rect 26146 25735 26202 25744
rect 26056 25152 26108 25158
rect 26056 25094 26108 25100
rect 25870 24712 25926 24721
rect 25870 24647 25926 24656
rect 25792 24568 25912 24596
rect 25318 23760 25374 23769
rect 25318 23695 25374 23704
rect 25320 23656 25372 23662
rect 25320 23598 25372 23604
rect 25226 23352 25282 23361
rect 25226 23287 25282 23296
rect 25134 22536 25190 22545
rect 25134 22471 25190 22480
rect 25148 20058 25176 22471
rect 25240 22098 25268 23287
rect 25228 22092 25280 22098
rect 25228 22034 25280 22040
rect 25226 21312 25282 21321
rect 25226 21247 25282 21256
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 25134 19816 25190 19825
rect 25134 19751 25190 19760
rect 25148 19446 25176 19751
rect 25136 19440 25188 19446
rect 25136 19382 25188 19388
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 25148 17921 25176 19246
rect 25240 18970 25268 21247
rect 25228 18964 25280 18970
rect 25228 18906 25280 18912
rect 25226 18456 25282 18465
rect 25226 18391 25282 18400
rect 25134 17912 25190 17921
rect 25134 17847 25190 17856
rect 24766 17711 24822 17720
rect 24952 17740 25004 17746
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 17134 24716 17478
rect 24676 17128 24728 17134
rect 24676 17070 24728 17076
rect 24676 16788 24728 16794
rect 24676 16730 24728 16736
rect 24216 16720 24268 16726
rect 24216 16662 24268 16668
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24044 15422 24164 15450
rect 23938 15328 23994 15337
rect 23938 15263 23994 15272
rect 24044 15094 24072 15422
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 24032 15088 24084 15094
rect 24032 15030 24084 15036
rect 24136 15026 24164 15302
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 24044 14346 24072 14758
rect 24136 14618 24164 14962
rect 24124 14612 24176 14618
rect 24124 14554 24176 14560
rect 24032 14340 24084 14346
rect 24032 14282 24084 14288
rect 24044 14074 24072 14282
rect 24124 14272 24176 14278
rect 24124 14214 24176 14220
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 24136 13938 24164 14214
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24308 13932 24360 13938
rect 24308 13874 24360 13880
rect 24032 13728 24084 13734
rect 24032 13670 24084 13676
rect 24044 13530 24072 13670
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 23848 13184 23900 13190
rect 23848 13126 23900 13132
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 23848 12912 23900 12918
rect 23848 12854 23900 12860
rect 24044 12866 24072 13126
rect 24136 12986 24164 13874
rect 24320 13394 24348 13874
rect 24688 13682 24716 16730
rect 24780 16266 24808 17711
rect 25056 17734 25176 17762
rect 24952 17682 25004 17688
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 24872 17241 24900 17478
rect 24858 17232 24914 17241
rect 24858 17167 24914 17176
rect 24964 16998 24992 17682
rect 24952 16992 25004 16998
rect 24952 16934 25004 16940
rect 25042 16824 25098 16833
rect 25042 16759 25044 16768
rect 25096 16759 25098 16768
rect 25044 16730 25096 16736
rect 24780 16250 24900 16266
rect 24780 16244 24912 16250
rect 24780 16238 24860 16244
rect 24860 16186 24912 16192
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24766 14920 24822 14929
rect 24766 14855 24822 14864
rect 24596 13654 24716 13682
rect 24596 13530 24624 13654
rect 24674 13560 24730 13569
rect 24584 13524 24636 13530
rect 24674 13495 24730 13504
rect 24584 13466 24636 13472
rect 24308 13388 24360 13394
rect 24308 13330 24360 13336
rect 24214 13288 24270 13297
rect 24214 13223 24270 13232
rect 24124 12980 24176 12986
rect 24124 12922 24176 12928
rect 23860 12442 23888 12854
rect 24044 12838 24164 12866
rect 24032 12776 24084 12782
rect 24032 12718 24084 12724
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 23768 10810 23796 12378
rect 23860 11354 23888 12378
rect 24044 12238 24072 12718
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 23938 12064 23994 12073
rect 23938 11999 23994 12008
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23756 10804 23808 10810
rect 23756 10746 23808 10752
rect 23754 10568 23810 10577
rect 23754 10503 23810 10512
rect 23768 10266 23796 10503
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23664 10124 23716 10130
rect 23664 10066 23716 10072
rect 23570 10024 23626 10033
rect 23400 9982 23520 10010
rect 23294 9959 23350 9968
rect 23204 9930 23256 9936
rect 23216 8650 23244 9930
rect 23294 9888 23350 9897
rect 23294 9823 23350 9832
rect 23308 9178 23336 9823
rect 23388 9376 23440 9382
rect 23492 9353 23520 9982
rect 23570 9959 23626 9968
rect 23676 9722 23704 10066
rect 23860 9722 23888 10406
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23848 9716 23900 9722
rect 23848 9658 23900 9664
rect 23662 9616 23718 9625
rect 23662 9551 23718 9560
rect 23848 9580 23900 9586
rect 23676 9518 23704 9551
rect 23848 9522 23900 9528
rect 23664 9512 23716 9518
rect 23570 9480 23626 9489
rect 23664 9454 23716 9460
rect 23570 9415 23626 9424
rect 23388 9318 23440 9324
rect 23478 9344 23534 9353
rect 23296 9172 23348 9178
rect 23296 9114 23348 9120
rect 23216 8622 23336 8650
rect 23204 8560 23256 8566
rect 23204 8502 23256 8508
rect 23112 4752 23164 4758
rect 23112 4694 23164 4700
rect 22836 4684 22888 4690
rect 22836 4626 22888 4632
rect 22522 4542 22600 4570
rect 22650 4584 22706 4593
rect 22466 4519 22522 4528
rect 22650 4519 22706 4528
rect 22650 4448 22706 4457
rect 22650 4383 22706 4392
rect 22466 4176 22522 4185
rect 22388 4134 22466 4162
rect 22466 4111 22522 4120
rect 22284 3188 22336 3194
rect 22284 3130 22336 3136
rect 22296 2990 22324 3130
rect 22480 2990 22508 4111
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 22284 2984 22336 2990
rect 22284 2926 22336 2932
rect 22468 2984 22520 2990
rect 22468 2926 22520 2932
rect 22282 2680 22338 2689
rect 22282 2615 22284 2624
rect 22336 2615 22338 2624
rect 22284 2586 22336 2592
rect 22572 2582 22600 4014
rect 22560 2576 22612 2582
rect 22560 2518 22612 2524
rect 22112 1414 22232 1442
rect 22112 480 22140 1414
rect 22664 480 22692 4383
rect 22742 4176 22798 4185
rect 22742 4111 22798 4120
rect 22756 2514 22784 4111
rect 22848 3942 22876 4626
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 22756 2417 22784 2450
rect 22742 2408 22798 2417
rect 22742 2343 22798 2352
rect 22848 1737 22876 3878
rect 22928 3528 22980 3534
rect 22928 3470 22980 3476
rect 22940 2446 22968 3470
rect 23032 3466 23060 4558
rect 23124 4282 23152 4694
rect 23112 4276 23164 4282
rect 23112 4218 23164 4224
rect 23020 3460 23072 3466
rect 23020 3402 23072 3408
rect 23032 2514 23060 3402
rect 23112 2848 23164 2854
rect 23112 2790 23164 2796
rect 23124 2689 23152 2790
rect 23110 2680 23166 2689
rect 23110 2615 23166 2624
rect 23020 2508 23072 2514
rect 23020 2450 23072 2456
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 22928 2304 22980 2310
rect 22928 2246 22980 2252
rect 22834 1728 22890 1737
rect 22834 1663 22890 1672
rect 22940 1465 22968 2246
rect 22926 1456 22982 1465
rect 22926 1391 22982 1400
rect 23216 480 23244 8502
rect 23308 7721 23336 8622
rect 23400 7970 23428 9318
rect 23478 9279 23534 9288
rect 23492 9178 23520 9279
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23478 9072 23534 9081
rect 23478 9007 23534 9016
rect 23492 8634 23520 9007
rect 23584 8906 23612 9415
rect 23754 9072 23810 9081
rect 23754 9007 23810 9016
rect 23572 8900 23624 8906
rect 23572 8842 23624 8848
rect 23664 8832 23716 8838
rect 23662 8800 23664 8809
rect 23716 8800 23718 8809
rect 23662 8735 23718 8744
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23492 8401 23520 8434
rect 23664 8424 23716 8430
rect 23478 8392 23534 8401
rect 23664 8366 23716 8372
rect 23478 8327 23534 8336
rect 23676 8265 23704 8366
rect 23662 8256 23718 8265
rect 23662 8191 23718 8200
rect 23662 7984 23718 7993
rect 23400 7954 23520 7970
rect 23400 7948 23532 7954
rect 23400 7942 23480 7948
rect 23662 7919 23718 7928
rect 23480 7890 23532 7896
rect 23388 7812 23440 7818
rect 23388 7754 23440 7760
rect 23294 7712 23350 7721
rect 23294 7647 23350 7656
rect 23296 7200 23348 7206
rect 23296 7142 23348 7148
rect 23308 6798 23336 7142
rect 23296 6792 23348 6798
rect 23296 6734 23348 6740
rect 23296 6180 23348 6186
rect 23296 6122 23348 6128
rect 23308 5681 23336 6122
rect 23400 5778 23428 7754
rect 23480 7744 23532 7750
rect 23480 7686 23532 7692
rect 23572 7744 23624 7750
rect 23572 7686 23624 7692
rect 23492 7449 23520 7686
rect 23478 7440 23534 7449
rect 23478 7375 23534 7384
rect 23478 7168 23534 7177
rect 23478 7103 23534 7112
rect 23388 5772 23440 5778
rect 23388 5714 23440 5720
rect 23294 5672 23350 5681
rect 23492 5642 23520 7103
rect 23584 5846 23612 7686
rect 23676 7002 23704 7919
rect 23664 6996 23716 7002
rect 23664 6938 23716 6944
rect 23768 6882 23796 9007
rect 23860 8809 23888 9522
rect 23952 9042 23980 11999
rect 24044 11898 24072 12174
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 24032 11552 24084 11558
rect 24030 11520 24032 11529
rect 24084 11520 24086 11529
rect 24030 11455 24086 11464
rect 24044 11150 24072 11455
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 24032 11008 24084 11014
rect 24032 10950 24084 10956
rect 24044 10538 24072 10950
rect 24032 10532 24084 10538
rect 24032 10474 24084 10480
rect 24044 10266 24072 10474
rect 24032 10260 24084 10266
rect 24032 10202 24084 10208
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 24044 9761 24072 9862
rect 24030 9752 24086 9761
rect 24030 9687 24086 9696
rect 23940 9036 23992 9042
rect 23992 8996 24072 9024
rect 23940 8978 23992 8984
rect 23940 8832 23992 8838
rect 23846 8800 23902 8809
rect 23940 8774 23992 8780
rect 23846 8735 23902 8744
rect 23952 8673 23980 8774
rect 23938 8664 23994 8673
rect 24044 8634 24072 8996
rect 23938 8599 23994 8608
rect 24032 8628 24084 8634
rect 24032 8570 24084 8576
rect 23848 8288 23900 8294
rect 23848 8230 23900 8236
rect 23860 7342 23888 8230
rect 24136 8090 24164 12838
rect 24228 12764 24256 13223
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24492 12912 24544 12918
rect 24492 12854 24544 12860
rect 24308 12776 24360 12782
rect 24228 12736 24308 12764
rect 24308 12718 24360 12724
rect 24214 12608 24270 12617
rect 24214 12543 24270 12552
rect 24228 11354 24256 12543
rect 24504 12442 24532 12854
rect 24688 12594 24716 13495
rect 24780 13002 24808 14855
rect 24872 13530 24900 15982
rect 24952 15564 25004 15570
rect 24952 15506 25004 15512
rect 24964 15162 24992 15506
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24872 13297 24900 13330
rect 24858 13288 24914 13297
rect 24858 13223 24914 13232
rect 24964 13190 24992 14350
rect 25044 14340 25096 14346
rect 25044 14282 25096 14288
rect 25056 14006 25084 14282
rect 25044 14000 25096 14006
rect 25044 13942 25096 13948
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 24780 12986 24900 13002
rect 24780 12980 24912 12986
rect 24780 12974 24860 12980
rect 24860 12922 24912 12928
rect 24688 12566 24808 12594
rect 24492 12436 24544 12442
rect 24780 12424 24808 12566
rect 24964 12481 24992 13126
rect 25056 12918 25084 13330
rect 25044 12912 25096 12918
rect 25044 12854 25096 12860
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 24950 12472 25006 12481
rect 24860 12436 24912 12442
rect 24780 12396 24860 12424
rect 24492 12378 24544 12384
rect 24950 12407 25006 12416
rect 24860 12378 24912 12384
rect 24858 12336 24914 12345
rect 24858 12271 24914 12280
rect 24952 12300 25004 12306
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24766 11928 24822 11937
rect 24766 11863 24822 11872
rect 24674 11656 24730 11665
rect 24674 11591 24730 11600
rect 24400 11552 24452 11558
rect 24400 11494 24452 11500
rect 24216 11348 24268 11354
rect 24216 11290 24268 11296
rect 24216 11212 24268 11218
rect 24216 11154 24268 11160
rect 24228 10470 24256 11154
rect 24412 11082 24440 11494
rect 24400 11076 24452 11082
rect 24400 11018 24452 11024
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24584 10736 24636 10742
rect 24584 10678 24636 10684
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 24216 10192 24268 10198
rect 24216 10134 24268 10140
rect 24124 8084 24176 8090
rect 24124 8026 24176 8032
rect 24032 7948 24084 7954
rect 24032 7890 24084 7896
rect 24044 7546 24072 7890
rect 24032 7540 24084 7546
rect 24032 7482 24084 7488
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 23940 7268 23992 7274
rect 23940 7210 23992 7216
rect 23676 6854 23796 6882
rect 23676 6254 23704 6854
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23768 6662 23796 6734
rect 23756 6656 23808 6662
rect 23756 6598 23808 6604
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23768 6322 23796 6598
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 23756 6180 23808 6186
rect 23756 6122 23808 6128
rect 23664 6112 23716 6118
rect 23664 6054 23716 6060
rect 23676 5914 23704 6054
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 23572 5840 23624 5846
rect 23572 5782 23624 5788
rect 23294 5607 23350 5616
rect 23480 5636 23532 5642
rect 23480 5578 23532 5584
rect 23662 5400 23718 5409
rect 23662 5335 23664 5344
rect 23716 5335 23718 5344
rect 23664 5306 23716 5312
rect 23664 4616 23716 4622
rect 23664 4558 23716 4564
rect 23296 4548 23348 4554
rect 23296 4490 23348 4496
rect 23388 4548 23440 4554
rect 23388 4490 23440 4496
rect 20166 96 20222 105
rect 20166 31 20222 40
rect 20442 0 20498 480
rect 20994 0 21050 480
rect 21546 0 21602 480
rect 22098 0 22154 480
rect 22650 0 22706 480
rect 23202 0 23258 480
rect 23308 377 23336 4490
rect 23400 4185 23428 4490
rect 23572 4480 23624 4486
rect 23572 4422 23624 4428
rect 23386 4176 23442 4185
rect 23386 4111 23442 4120
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23388 3936 23440 3942
rect 23492 3924 23520 4082
rect 23440 3896 23520 3924
rect 23388 3878 23440 3884
rect 23400 785 23428 3878
rect 23584 3738 23612 4422
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 23480 3664 23532 3670
rect 23478 3632 23480 3641
rect 23532 3632 23534 3641
rect 23676 3618 23704 4558
rect 23768 4078 23796 6122
rect 23860 4457 23888 6598
rect 23952 6089 23980 7210
rect 24044 7002 24072 7482
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 24032 6996 24084 7002
rect 24032 6938 24084 6944
rect 24032 6860 24084 6866
rect 24032 6802 24084 6808
rect 24044 6769 24072 6802
rect 24030 6760 24086 6769
rect 24030 6695 24086 6704
rect 24044 6458 24072 6695
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 23938 6080 23994 6089
rect 23938 6015 23994 6024
rect 24044 5930 24072 6258
rect 23952 5902 24072 5930
rect 23952 5710 23980 5902
rect 23940 5704 23992 5710
rect 23940 5646 23992 5652
rect 23952 5234 23980 5646
rect 24030 5400 24086 5409
rect 24030 5335 24086 5344
rect 23940 5228 23992 5234
rect 23940 5170 23992 5176
rect 24044 5166 24072 5335
rect 24032 5160 24084 5166
rect 24032 5102 24084 5108
rect 24044 4826 24072 5102
rect 24032 4820 24084 4826
rect 24032 4762 24084 4768
rect 23846 4448 23902 4457
rect 23846 4383 23902 4392
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 23940 4004 23992 4010
rect 23940 3946 23992 3952
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23478 3567 23534 3576
rect 23584 3590 23704 3618
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23492 2582 23520 3334
rect 23584 3126 23612 3590
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 23676 3194 23704 3470
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 23572 3120 23624 3126
rect 23572 3062 23624 3068
rect 23768 2990 23796 3878
rect 23848 3392 23900 3398
rect 23848 3334 23900 3340
rect 23860 3097 23888 3334
rect 23846 3088 23902 3097
rect 23846 3023 23902 3032
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23756 2984 23808 2990
rect 23756 2926 23808 2932
rect 23480 2576 23532 2582
rect 23480 2518 23532 2524
rect 23584 1465 23612 2926
rect 23756 2848 23808 2854
rect 23756 2790 23808 2796
rect 23570 1456 23626 1465
rect 23570 1391 23626 1400
rect 23386 776 23442 785
rect 23386 711 23442 720
rect 23768 480 23796 2790
rect 23952 2650 23980 3946
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 24044 3466 24072 3878
rect 24032 3460 24084 3466
rect 24032 3402 24084 3408
rect 24030 3224 24086 3233
rect 24030 3159 24086 3168
rect 24044 3058 24072 3159
rect 24032 3052 24084 3058
rect 24032 2994 24084 3000
rect 24030 2816 24086 2825
rect 24030 2751 24086 2760
rect 23940 2644 23992 2650
rect 23940 2586 23992 2592
rect 23938 2272 23994 2281
rect 23938 2207 23994 2216
rect 23952 1737 23980 2207
rect 23938 1728 23994 1737
rect 23938 1663 23994 1672
rect 24044 1057 24072 2751
rect 24030 1048 24086 1057
rect 24030 983 24086 992
rect 24136 898 24164 7142
rect 24228 4622 24256 10134
rect 24596 10130 24624 10678
rect 24584 10124 24636 10130
rect 24584 10066 24636 10072
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24308 9444 24360 9450
rect 24308 9386 24360 9392
rect 24320 9178 24348 9386
rect 24308 9172 24360 9178
rect 24308 9114 24360 9120
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24308 6248 24360 6254
rect 24308 6190 24360 6196
rect 24582 6216 24638 6225
rect 24320 5846 24348 6190
rect 24582 6151 24638 6160
rect 24308 5840 24360 5846
rect 24308 5782 24360 5788
rect 24596 5710 24624 6151
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24308 5228 24360 5234
rect 24308 5170 24360 5176
rect 24320 4826 24348 5170
rect 24308 4820 24360 4826
rect 24308 4762 24360 4768
rect 24688 4690 24716 11591
rect 24780 10810 24808 11863
rect 24872 11354 24900 12271
rect 24952 12242 25004 12248
rect 24964 11898 24992 12242
rect 24952 11892 25004 11898
rect 24952 11834 25004 11840
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 25056 11064 25084 12718
rect 24964 11036 25084 11064
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24768 10600 24820 10606
rect 24768 10542 24820 10548
rect 24780 10266 24808 10542
rect 24768 10260 24820 10266
rect 24768 10202 24820 10208
rect 24964 10198 24992 11036
rect 25042 10976 25098 10985
rect 25042 10911 25098 10920
rect 25056 10266 25084 10911
rect 25044 10260 25096 10266
rect 25044 10202 25096 10208
rect 24952 10192 25004 10198
rect 24952 10134 25004 10140
rect 24768 10124 24820 10130
rect 24768 10066 24820 10072
rect 24780 9722 24808 10066
rect 24768 9716 24820 9722
rect 24768 9658 24820 9664
rect 25042 9616 25098 9625
rect 25042 9551 25098 9560
rect 24860 9512 24912 9518
rect 24860 9454 24912 9460
rect 24766 8392 24822 8401
rect 24766 8327 24822 8336
rect 24780 7426 24808 8327
rect 24872 8129 24900 9454
rect 25056 9178 25084 9551
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 25148 8634 25176 17734
rect 25240 15706 25268 18391
rect 25332 17066 25360 23598
rect 25410 23080 25466 23089
rect 25410 23015 25466 23024
rect 25424 21690 25452 23015
rect 25686 21856 25742 21865
rect 25686 21791 25742 21800
rect 25412 21684 25464 21690
rect 25412 21626 25464 21632
rect 25502 20632 25558 20641
rect 25502 20567 25558 20576
rect 25410 20088 25466 20097
rect 25410 20023 25466 20032
rect 25424 17882 25452 20023
rect 25516 18426 25544 20567
rect 25596 19372 25648 19378
rect 25596 19314 25648 19320
rect 25504 18420 25556 18426
rect 25504 18362 25556 18368
rect 25502 18320 25558 18329
rect 25502 18255 25558 18264
rect 25412 17876 25464 17882
rect 25412 17818 25464 17824
rect 25412 17536 25464 17542
rect 25412 17478 25464 17484
rect 25320 17060 25372 17066
rect 25320 17002 25372 17008
rect 25320 16652 25372 16658
rect 25320 16594 25372 16600
rect 25332 15978 25360 16594
rect 25320 15972 25372 15978
rect 25320 15914 25372 15920
rect 25424 15858 25452 17478
rect 25516 16250 25544 18255
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25332 15830 25452 15858
rect 25228 15700 25280 15706
rect 25228 15642 25280 15648
rect 25332 15552 25360 15830
rect 25410 15736 25466 15745
rect 25410 15671 25466 15680
rect 25240 15524 25360 15552
rect 25240 14006 25268 15524
rect 25318 15464 25374 15473
rect 25318 15399 25374 15408
rect 25228 14000 25280 14006
rect 25228 13942 25280 13948
rect 25228 13864 25280 13870
rect 25226 13832 25228 13841
rect 25280 13832 25282 13841
rect 25226 13767 25282 13776
rect 25332 13530 25360 15399
rect 25424 14074 25452 15671
rect 25504 15632 25556 15638
rect 25502 15600 25504 15609
rect 25556 15600 25558 15609
rect 25502 15535 25558 15544
rect 25504 14476 25556 14482
rect 25504 14418 25556 14424
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25412 13932 25464 13938
rect 25412 13874 25464 13880
rect 25320 13524 25372 13530
rect 25320 13466 25372 13472
rect 25424 13410 25452 13874
rect 25240 13382 25452 13410
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 24858 8120 24914 8129
rect 24858 8055 24914 8064
rect 25042 8120 25098 8129
rect 25042 8055 25044 8064
rect 25096 8055 25098 8064
rect 25044 8026 25096 8032
rect 25240 7954 25268 13382
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25332 12646 25360 13262
rect 25516 13190 25544 14418
rect 25504 13184 25556 13190
rect 25410 13152 25466 13161
rect 25504 13126 25556 13132
rect 25410 13087 25466 13096
rect 25320 12640 25372 12646
rect 25320 12582 25372 12588
rect 25424 11898 25452 13087
rect 25516 12753 25544 13126
rect 25502 12744 25558 12753
rect 25502 12679 25558 12688
rect 25608 12628 25636 19314
rect 25700 19174 25728 21791
rect 25780 21344 25832 21350
rect 25780 21286 25832 21292
rect 25792 20262 25820 21286
rect 25780 20256 25832 20262
rect 25780 20198 25832 20204
rect 25778 19544 25834 19553
rect 25778 19479 25834 19488
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25686 19000 25742 19009
rect 25686 18935 25742 18944
rect 25700 16794 25728 18935
rect 25792 17338 25820 19479
rect 25780 17332 25832 17338
rect 25780 17274 25832 17280
rect 25688 16788 25740 16794
rect 25688 16730 25740 16736
rect 25884 16402 25912 24568
rect 25964 20392 26016 20398
rect 25962 20360 25964 20369
rect 26016 20360 26018 20369
rect 25962 20295 26018 20304
rect 25964 20256 26016 20262
rect 25964 20198 26016 20204
rect 25976 17542 26004 20198
rect 25964 17536 26016 17542
rect 25964 17478 26016 17484
rect 25962 17232 26018 17241
rect 25962 17167 26018 17176
rect 25516 12600 25636 12628
rect 25700 16374 25912 16402
rect 25412 11892 25464 11898
rect 25412 11834 25464 11840
rect 25318 10024 25374 10033
rect 25318 9959 25374 9968
rect 25228 7948 25280 7954
rect 25228 7890 25280 7896
rect 25136 7744 25188 7750
rect 25136 7686 25188 7692
rect 24780 7398 24900 7426
rect 24768 7336 24820 7342
rect 24768 7278 24820 7284
rect 24780 7002 24808 7278
rect 24768 6996 24820 7002
rect 24768 6938 24820 6944
rect 24872 6882 24900 7398
rect 24780 6854 24900 6882
rect 25042 6896 25098 6905
rect 24780 6254 24808 6854
rect 25042 6831 25098 6840
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24780 5370 24808 5646
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 24216 4616 24268 4622
rect 24216 4558 24268 4564
rect 24216 4480 24268 4486
rect 24216 4422 24268 4428
rect 24228 3913 24256 4422
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24688 4282 24716 4626
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 24214 3904 24270 3913
rect 24214 3839 24270 3848
rect 24780 3738 24808 4422
rect 24768 3732 24820 3738
rect 24768 3674 24820 3680
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24688 3194 24716 3470
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24216 3120 24268 3126
rect 24688 3074 24716 3130
rect 24216 3062 24268 3068
rect 24228 2854 24256 3062
rect 24308 3052 24360 3058
rect 24308 2994 24360 3000
rect 24596 3046 24716 3074
rect 24216 2848 24268 2854
rect 24216 2790 24268 2796
rect 24320 2514 24348 2994
rect 24490 2544 24546 2553
rect 24308 2508 24360 2514
rect 24490 2479 24492 2488
rect 24308 2450 24360 2456
rect 24544 2479 24546 2488
rect 24492 2450 24544 2456
rect 24596 2446 24624 3046
rect 24676 2984 24728 2990
rect 24676 2926 24728 2932
rect 24688 2514 24716 2926
rect 24780 2582 24808 3334
rect 24768 2576 24820 2582
rect 24768 2518 24820 2524
rect 24676 2508 24728 2514
rect 24676 2450 24728 2456
rect 24584 2440 24636 2446
rect 24636 2388 24716 2394
rect 24584 2382 24716 2388
rect 24596 2366 24716 2382
rect 24596 2317 24624 2366
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24688 1601 24716 2366
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 24674 1592 24730 1601
rect 24674 1527 24730 1536
rect 24136 870 24348 898
rect 24320 480 24348 870
rect 24780 649 24808 2246
rect 24766 640 24822 649
rect 24766 575 24822 584
rect 24872 480 24900 6598
rect 25056 6458 25084 6831
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 25056 6254 25084 6394
rect 25044 6248 25096 6254
rect 25044 6190 25096 6196
rect 25044 5772 25096 5778
rect 25044 5714 25096 5720
rect 24952 5636 25004 5642
rect 24952 5578 25004 5584
rect 24964 5001 24992 5578
rect 25056 5370 25084 5714
rect 25044 5364 25096 5370
rect 25044 5306 25096 5312
rect 24950 4992 25006 5001
rect 24950 4927 25006 4936
rect 25044 4752 25096 4758
rect 25042 4720 25044 4729
rect 25096 4720 25098 4729
rect 25042 4655 25098 4664
rect 24950 4176 25006 4185
rect 24950 4111 24952 4120
rect 25004 4111 25006 4120
rect 24952 4082 25004 4088
rect 25044 4072 25096 4078
rect 25042 4040 25044 4049
rect 25096 4040 25098 4049
rect 25042 3975 25098 3984
rect 25148 3040 25176 7686
rect 25240 7546 25268 7890
rect 25332 7834 25360 9959
rect 25410 9616 25466 9625
rect 25410 9551 25466 9560
rect 25424 9178 25452 9551
rect 25412 9172 25464 9178
rect 25412 9114 25464 9120
rect 25332 7806 25452 7834
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25228 7540 25280 7546
rect 25228 7482 25280 7488
rect 25228 6792 25280 6798
rect 25228 6734 25280 6740
rect 25240 5302 25268 6734
rect 25228 5296 25280 5302
rect 25228 5238 25280 5244
rect 25228 5024 25280 5030
rect 25228 4966 25280 4972
rect 25240 4282 25268 4966
rect 25228 4276 25280 4282
rect 25228 4218 25280 4224
rect 25332 4049 25360 7686
rect 25424 5778 25452 7806
rect 25516 7546 25544 12600
rect 25594 12336 25650 12345
rect 25594 12271 25596 12280
rect 25648 12271 25650 12280
rect 25596 12242 25648 12248
rect 25594 10976 25650 10985
rect 25594 10911 25650 10920
rect 25608 10810 25636 10911
rect 25596 10804 25648 10810
rect 25596 10746 25648 10752
rect 25700 8634 25728 16374
rect 25780 16244 25832 16250
rect 25780 16186 25832 16192
rect 25792 14906 25820 16186
rect 25872 15972 25924 15978
rect 25872 15914 25924 15920
rect 25884 15042 25912 15914
rect 25976 15162 26004 17167
rect 25964 15156 26016 15162
rect 25964 15098 26016 15104
rect 25884 15014 26004 15042
rect 25792 14878 25912 14906
rect 25780 14272 25832 14278
rect 25780 14214 25832 14220
rect 25792 13977 25820 14214
rect 25778 13968 25834 13977
rect 25884 13938 25912 14878
rect 25778 13903 25834 13912
rect 25872 13932 25924 13938
rect 25872 13874 25924 13880
rect 25872 13796 25924 13802
rect 25872 13738 25924 13744
rect 25884 13530 25912 13738
rect 25872 13524 25924 13530
rect 25872 13466 25924 13472
rect 25778 13424 25834 13433
rect 25778 13359 25834 13368
rect 25792 12238 25820 13359
rect 25870 13288 25926 13297
rect 25870 13223 25926 13232
rect 25780 12232 25832 12238
rect 25780 12174 25832 12180
rect 25778 10432 25834 10441
rect 25778 10367 25834 10376
rect 25792 10266 25820 10367
rect 25780 10260 25832 10266
rect 25780 10202 25832 10208
rect 25778 9480 25834 9489
rect 25778 9415 25834 9424
rect 25792 9178 25820 9415
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 25688 8628 25740 8634
rect 25688 8570 25740 8576
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25504 7540 25556 7546
rect 25504 7482 25556 7488
rect 25700 7041 25728 7686
rect 25686 7032 25742 7041
rect 25686 6967 25742 6976
rect 25780 6724 25832 6730
rect 25780 6666 25832 6672
rect 25792 6458 25820 6666
rect 25780 6452 25832 6458
rect 25780 6394 25832 6400
rect 25688 6112 25740 6118
rect 25688 6054 25740 6060
rect 25412 5772 25464 5778
rect 25412 5714 25464 5720
rect 25412 5568 25464 5574
rect 25412 5510 25464 5516
rect 25424 4865 25452 5510
rect 25502 4992 25558 5001
rect 25502 4927 25558 4936
rect 25410 4856 25466 4865
rect 25410 4791 25466 4800
rect 25318 4040 25374 4049
rect 25318 3975 25374 3984
rect 25412 3936 25464 3942
rect 25412 3878 25464 3884
rect 25226 3768 25282 3777
rect 25226 3703 25282 3712
rect 24964 3012 25176 3040
rect 24964 610 24992 3012
rect 25134 2952 25190 2961
rect 25134 2887 25190 2896
rect 25148 2854 25176 2887
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 25136 2848 25188 2854
rect 25240 2825 25268 3703
rect 25424 3505 25452 3878
rect 25410 3496 25466 3505
rect 25410 3431 25466 3440
rect 25136 2790 25188 2796
rect 25226 2816 25282 2825
rect 25056 1329 25084 2790
rect 25226 2751 25282 2760
rect 25516 2310 25544 4927
rect 25700 2922 25728 6054
rect 25780 5772 25832 5778
rect 25780 5714 25832 5720
rect 25792 2990 25820 5714
rect 25884 5370 25912 13223
rect 25976 10577 26004 15014
rect 26068 11898 26096 25094
rect 26160 17338 26188 25735
rect 26528 24449 26556 27520
rect 26608 26036 26660 26042
rect 26608 25978 26660 25984
rect 26514 24440 26570 24449
rect 26514 24375 26570 24384
rect 26332 19780 26384 19786
rect 26332 19722 26384 19728
rect 26148 17332 26200 17338
rect 26148 17274 26200 17280
rect 26148 17060 26200 17066
rect 26148 17002 26200 17008
rect 26056 11892 26108 11898
rect 26056 11834 26108 11840
rect 25962 10568 26018 10577
rect 25962 10503 26018 10512
rect 25962 9616 26018 9625
rect 25962 9551 26018 9560
rect 25976 8634 26004 9551
rect 26056 9376 26108 9382
rect 26056 9318 26108 9324
rect 26068 8974 26096 9318
rect 26056 8968 26108 8974
rect 26056 8910 26108 8916
rect 25964 8628 26016 8634
rect 25964 8570 26016 8576
rect 26160 8566 26188 17002
rect 26240 16040 26292 16046
rect 26238 16008 26240 16017
rect 26292 16008 26294 16017
rect 26238 15943 26294 15952
rect 26240 15088 26292 15094
rect 26238 15056 26240 15065
rect 26292 15056 26294 15065
rect 26238 14991 26294 15000
rect 26240 14408 26292 14414
rect 26238 14376 26240 14385
rect 26292 14376 26294 14385
rect 26238 14311 26294 14320
rect 26238 13696 26294 13705
rect 26238 13631 26294 13640
rect 26252 13530 26280 13631
rect 26240 13524 26292 13530
rect 26240 13466 26292 13472
rect 26240 11824 26292 11830
rect 26238 11792 26240 11801
rect 26292 11792 26294 11801
rect 26238 11727 26294 11736
rect 26238 9208 26294 9217
rect 26238 9143 26240 9152
rect 26292 9143 26294 9152
rect 26240 9114 26292 9120
rect 26344 8634 26372 19722
rect 26620 14074 26648 25978
rect 27080 23497 27108 27520
rect 27632 23905 27660 27520
rect 27618 23896 27674 23905
rect 27618 23831 27674 23840
rect 27066 23488 27122 23497
rect 27066 23423 27122 23432
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26424 9376 26476 9382
rect 26424 9318 26476 9324
rect 26436 8945 26464 9318
rect 26422 8936 26478 8945
rect 26422 8871 26478 8880
rect 26332 8628 26384 8634
rect 26332 8570 26384 8576
rect 26148 8560 26200 8566
rect 26148 8502 26200 8508
rect 26056 7880 26108 7886
rect 26054 7848 26056 7857
rect 26108 7848 26110 7857
rect 26054 7783 26110 7792
rect 25964 7200 26016 7206
rect 25964 7142 26016 7148
rect 26148 7200 26200 7206
rect 26424 7200 26476 7206
rect 26148 7142 26200 7148
rect 26422 7168 26424 7177
rect 26476 7168 26478 7177
rect 25872 5364 25924 5370
rect 25872 5306 25924 5312
rect 25884 5166 25912 5306
rect 25872 5160 25924 5166
rect 25872 5102 25924 5108
rect 25780 2984 25832 2990
rect 25780 2926 25832 2932
rect 25688 2916 25740 2922
rect 25688 2858 25740 2864
rect 25504 2304 25556 2310
rect 25504 2246 25556 2252
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 25792 1873 25820 2246
rect 25778 1864 25834 1873
rect 25778 1799 25834 1808
rect 25042 1320 25098 1329
rect 25042 1255 25098 1264
rect 24952 604 25004 610
rect 24952 546 25004 552
rect 25412 604 25464 610
rect 25412 546 25464 552
rect 25424 480 25452 546
rect 25976 480 26004 7142
rect 26056 6656 26108 6662
rect 26056 6598 26108 6604
rect 26068 513 26096 6598
rect 26160 1737 26188 7142
rect 26422 7103 26478 7112
rect 26240 6112 26292 6118
rect 26240 6054 26292 6060
rect 26252 5953 26280 6054
rect 26238 5944 26294 5953
rect 26238 5879 26294 5888
rect 26240 5840 26292 5846
rect 26238 5808 26240 5817
rect 26292 5808 26294 5817
rect 26238 5743 26294 5752
rect 26240 4480 26292 4486
rect 26240 4422 26292 4428
rect 26252 4214 26280 4422
rect 26240 4208 26292 4214
rect 26240 4150 26292 4156
rect 27066 4040 27122 4049
rect 27066 3975 27122 3984
rect 26514 3904 26570 3913
rect 26514 3839 26570 3848
rect 26238 3088 26294 3097
rect 26238 3023 26240 3032
rect 26292 3023 26294 3032
rect 26240 2994 26292 3000
rect 26422 2544 26478 2553
rect 26422 2479 26424 2488
rect 26476 2479 26478 2488
rect 26424 2450 26476 2456
rect 26146 1728 26202 1737
rect 26146 1663 26202 1672
rect 26054 504 26110 513
rect 23294 368 23350 377
rect 23294 303 23350 312
rect 23754 0 23810 480
rect 24306 0 24362 480
rect 24858 0 24914 480
rect 25410 0 25466 480
rect 25962 0 26018 480
rect 26528 480 26556 3839
rect 27080 480 27108 3975
rect 27618 3496 27674 3505
rect 27618 3431 27674 3440
rect 27632 480 27660 3431
rect 26054 439 26110 448
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 1122 27648 1178 27704
rect 662 27104 718 27160
rect 662 24384 718 24440
rect 570 20032 626 20088
rect 1030 25880 1086 25936
rect 938 24792 994 24848
rect 23754 27648 23810 27704
rect 1306 26560 1362 26616
rect 1214 24112 1270 24168
rect 1398 18944 1454 19000
rect 1582 18264 1638 18320
rect 1950 23704 2006 23760
rect 2134 24556 2136 24576
rect 2136 24556 2188 24576
rect 2188 24556 2190 24576
rect 2134 24520 2190 24556
rect 2226 24268 2282 24304
rect 2226 24248 2228 24268
rect 2228 24248 2280 24268
rect 2280 24248 2282 24268
rect 1858 22072 1914 22128
rect 18 12280 74 12336
rect 1950 17040 2006 17096
rect 1766 16088 1822 16144
rect 1674 15272 1730 15328
rect 1582 15000 1638 15056
rect 1582 14864 1638 14920
rect 1490 10920 1546 10976
rect 2134 17312 2190 17368
rect 2042 16496 2098 16552
rect 1766 12300 1822 12336
rect 1766 12280 1768 12300
rect 1768 12280 1820 12300
rect 1820 12280 1822 12300
rect 2410 24692 2412 24712
rect 2412 24692 2464 24712
rect 2464 24692 2466 24712
rect 2410 24656 2466 24692
rect 2410 20712 2466 20768
rect 2410 20304 2466 20360
rect 2502 17448 2558 17504
rect 2410 16632 2466 16688
rect 2410 16396 2412 16416
rect 2412 16396 2464 16416
rect 2464 16396 2466 16416
rect 2410 16360 2466 16396
rect 2778 25336 2834 25392
rect 3238 24656 3294 24712
rect 2870 21256 2926 21312
rect 2870 20168 2926 20224
rect 3514 23044 3570 23080
rect 3514 23024 3516 23044
rect 3516 23024 3568 23044
rect 3568 23024 3570 23044
rect 3330 22380 3332 22400
rect 3332 22380 3384 22400
rect 3384 22380 3386 22400
rect 3330 22344 3386 22380
rect 3422 21664 3478 21720
rect 3238 21528 3294 21584
rect 3422 21392 3478 21448
rect 3238 20984 3294 21040
rect 2778 18964 2834 19000
rect 2778 18944 2780 18964
rect 2780 18944 2832 18964
rect 2832 18944 2834 18964
rect 2410 15136 2466 15192
rect 2410 14612 2466 14648
rect 2410 14592 2412 14612
rect 2412 14592 2464 14612
rect 2464 14592 2466 14612
rect 2042 13096 2098 13152
rect 1950 12008 2006 12064
rect 1858 11600 1914 11656
rect 2410 12416 2466 12472
rect 2778 16904 2834 16960
rect 2962 17176 3018 17232
rect 3514 20440 3570 20496
rect 3790 24792 3846 24848
rect 3882 23704 3938 23760
rect 3974 23568 4030 23624
rect 3698 21800 3754 21856
rect 4066 23432 4122 23488
rect 4250 23840 4306 23896
rect 4250 23568 4306 23624
rect 4066 22480 4122 22536
rect 4342 22888 4398 22944
rect 4342 22616 4398 22672
rect 3054 16632 3110 16688
rect 3146 16496 3202 16552
rect 3146 15816 3202 15872
rect 2226 11736 2282 11792
rect 2042 11192 2098 11248
rect 2042 10532 2098 10568
rect 2042 10512 2044 10532
rect 2044 10512 2096 10532
rect 2096 10512 2098 10532
rect 1398 9968 1454 10024
rect 1398 9560 1454 9616
rect 1766 9596 1768 9616
rect 1768 9596 1820 9616
rect 1820 9596 1822 9616
rect 1766 9560 1822 9596
rect 662 3032 718 3088
rect 202 1672 258 1728
rect 2410 12164 2466 12200
rect 2410 12144 2412 12164
rect 2412 12144 2464 12164
rect 2464 12144 2466 12164
rect 2318 10240 2374 10296
rect 2134 9444 2190 9480
rect 2134 9424 2136 9444
rect 2136 9424 2188 9444
rect 2188 9424 2190 9444
rect 2042 9288 2098 9344
rect 1950 8744 2006 8800
rect 1858 8472 1914 8528
rect 2410 9172 2466 9208
rect 2410 9152 2412 9172
rect 2412 9152 2464 9172
rect 2464 9152 2466 9172
rect 2134 9016 2190 9072
rect 2042 7404 2098 7440
rect 2042 7384 2044 7404
rect 2044 7384 2096 7404
rect 2096 7384 2098 7404
rect 1582 6976 1638 7032
rect 1858 6160 1914 6216
rect 2686 12280 2742 12336
rect 2870 11464 2926 11520
rect 3698 17584 3754 17640
rect 3790 16124 3792 16144
rect 3792 16124 3844 16144
rect 3844 16124 3846 16144
rect 3790 16088 3846 16124
rect 4158 18828 4214 18864
rect 4158 18808 4160 18828
rect 4160 18808 4212 18828
rect 4212 18808 4214 18828
rect 4066 18264 4122 18320
rect 4158 17448 4214 17504
rect 4342 18300 4344 18320
rect 4344 18300 4396 18320
rect 4396 18300 4398 18320
rect 4342 18264 4398 18300
rect 4250 16768 4306 16824
rect 4066 16632 4122 16688
rect 4066 15952 4122 16008
rect 3974 15408 4030 15464
rect 3790 15136 3846 15192
rect 3790 13504 3846 13560
rect 3790 13368 3846 13424
rect 4250 14884 4306 14920
rect 4250 14864 4252 14884
rect 4252 14864 4304 14884
rect 4304 14864 4306 14884
rect 4250 13640 4306 13696
rect 3698 12552 3754 12608
rect 3606 12416 3662 12472
rect 3606 11600 3662 11656
rect 3514 10920 3570 10976
rect 3514 10376 3570 10432
rect 2870 8916 2872 8936
rect 2872 8916 2924 8936
rect 2924 8916 2926 8936
rect 2870 8880 2926 8916
rect 2502 8064 2558 8120
rect 2410 7692 2412 7712
rect 2412 7692 2464 7712
rect 2464 7692 2466 7712
rect 2410 7656 2466 7692
rect 2410 6724 2466 6760
rect 2410 6704 2412 6724
rect 2412 6704 2464 6724
rect 2464 6704 2466 6724
rect 1858 4392 1914 4448
rect 2318 5208 2374 5264
rect 2594 6196 2596 6216
rect 2596 6196 2648 6216
rect 2648 6196 2650 6216
rect 2594 6160 2650 6196
rect 3238 9696 3294 9752
rect 3146 8472 3202 8528
rect 2962 7792 3018 7848
rect 2686 6024 2742 6080
rect 2226 4120 2282 4176
rect 2778 4664 2834 4720
rect 1582 2252 1584 2272
rect 1584 2252 1636 2272
rect 1636 2252 1638 2272
rect 1582 2216 1638 2252
rect 1490 720 1546 776
rect 1950 1808 2006 1864
rect 3422 9152 3478 9208
rect 3330 8608 3386 8664
rect 3330 8472 3386 8528
rect 3054 5208 3110 5264
rect 3422 7520 3478 7576
rect 3790 12416 3846 12472
rect 3974 12960 4030 13016
rect 4066 12844 4122 12880
rect 4066 12824 4068 12844
rect 4068 12824 4120 12844
rect 4120 12824 4122 12844
rect 4066 12708 4122 12744
rect 4066 12688 4068 12708
rect 4068 12688 4120 12708
rect 4120 12688 4122 12708
rect 3974 12144 4030 12200
rect 3974 11872 4030 11928
rect 3698 9560 3754 9616
rect 3790 8880 3846 8936
rect 3698 7828 3700 7848
rect 3700 7828 3752 7848
rect 3752 7828 3754 7848
rect 3698 7792 3754 7828
rect 3514 6840 3570 6896
rect 3422 5888 3478 5944
rect 3146 3168 3202 3224
rect 4158 9560 4214 9616
rect 4066 8880 4122 8936
rect 4066 6996 4122 7032
rect 4066 6976 4068 6996
rect 4068 6976 4120 6996
rect 4120 6976 4122 6996
rect 4158 4664 4214 4720
rect 4066 4528 4122 4584
rect 3882 4004 3938 4040
rect 3882 3984 3884 4004
rect 3884 3984 3936 4004
rect 3936 3984 3938 4004
rect 2962 2896 3018 2952
rect 2502 1264 2558 1320
rect 4158 3712 4214 3768
rect 3790 2896 3846 2952
rect 3698 2524 3700 2544
rect 3700 2524 3752 2544
rect 3752 2524 3754 2544
rect 3698 2488 3754 2524
rect 4066 1944 4122 2000
rect 4066 1536 4122 1592
rect 4802 24656 4858 24712
rect 4618 12044 4620 12064
rect 4620 12044 4672 12064
rect 4672 12044 4674 12064
rect 4618 12008 4674 12044
rect 5170 24792 5226 24848
rect 4894 22072 4950 22128
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 6366 26016 6422 26072
rect 6182 24284 6184 24304
rect 6184 24284 6236 24304
rect 6236 24284 6238 24304
rect 6182 24248 6238 24284
rect 5170 17856 5226 17912
rect 4802 14456 4858 14512
rect 4802 11620 4858 11656
rect 4802 11600 4804 11620
rect 4804 11600 4856 11620
rect 4856 11600 4858 11620
rect 4526 9696 4582 9752
rect 4710 9560 4766 9616
rect 5078 17720 5134 17776
rect 4986 16768 5042 16824
rect 4986 13948 4988 13968
rect 4988 13948 5040 13968
rect 5040 13948 5042 13968
rect 4986 13912 5042 13948
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5630 22380 5632 22400
rect 5632 22380 5684 22400
rect 5684 22380 5686 22400
rect 5630 22344 5686 22380
rect 6366 23840 6422 23896
rect 6182 22752 6238 22808
rect 6366 22888 6422 22944
rect 5998 21936 6054 21992
rect 5998 21800 6054 21856
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5998 21392 6054 21448
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5814 20340 5816 20360
rect 5816 20340 5868 20360
rect 5868 20340 5870 20360
rect 5814 20304 5870 20340
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 6090 20168 6146 20224
rect 5998 18672 6054 18728
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5630 17720 5686 17776
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5170 15952 5226 16008
rect 5170 13096 5226 13152
rect 5170 12552 5226 12608
rect 5170 10684 5172 10704
rect 5172 10684 5224 10704
rect 5224 10684 5226 10704
rect 5170 10648 5226 10684
rect 4710 8608 4766 8664
rect 5078 8472 5134 8528
rect 4434 7656 4490 7712
rect 4526 3732 4582 3768
rect 4526 3712 4528 3732
rect 4528 3712 4580 3732
rect 4580 3712 4582 3732
rect 4342 1400 4398 1456
rect 4066 856 4122 912
rect 3882 312 3938 368
rect 4986 6568 5042 6624
rect 5446 16768 5502 16824
rect 5354 16360 5410 16416
rect 6182 19624 6238 19680
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5446 15680 5502 15736
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5354 13776 5410 13832
rect 5446 13232 5502 13288
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 6642 24248 6698 24304
rect 6826 23704 6882 23760
rect 7010 23468 7012 23488
rect 7012 23468 7064 23488
rect 7064 23468 7066 23488
rect 7010 23432 7066 23468
rect 7286 23704 7342 23760
rect 7470 23296 7526 23352
rect 6274 15544 6330 15600
rect 6458 17584 6514 17640
rect 6366 14764 6368 14784
rect 6368 14764 6420 14784
rect 6420 14764 6422 14784
rect 5998 13640 6054 13696
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5722 12416 5778 12472
rect 6366 14728 6422 14764
rect 6182 14612 6238 14648
rect 6182 14592 6184 14612
rect 6184 14592 6236 14612
rect 6236 14592 6238 14612
rect 6366 14592 6422 14648
rect 5446 12280 5502 12336
rect 5538 12144 5594 12200
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5538 10140 5540 10160
rect 5540 10140 5592 10160
rect 5592 10140 5594 10160
rect 5538 10104 5594 10140
rect 5906 10376 5962 10432
rect 5814 10124 5870 10160
rect 5814 10104 5816 10124
rect 5816 10104 5868 10124
rect 5868 10104 5870 10124
rect 5354 9832 5410 9888
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5906 9152 5962 9208
rect 5814 9052 5816 9072
rect 5816 9052 5868 9072
rect 5868 9052 5870 9072
rect 5170 7404 5226 7440
rect 5170 7384 5172 7404
rect 5172 7384 5224 7404
rect 5224 7384 5226 7404
rect 5814 9016 5870 9052
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5630 8472 5686 8528
rect 5538 8200 5594 8256
rect 5354 7520 5410 7576
rect 5354 7112 5410 7168
rect 5262 6840 5318 6896
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5170 5752 5226 5808
rect 5354 6024 5410 6080
rect 6090 12008 6146 12064
rect 6090 11872 6146 11928
rect 6366 12552 6422 12608
rect 6550 12824 6606 12880
rect 6458 12144 6514 12200
rect 6458 10260 6514 10296
rect 6458 10240 6460 10260
rect 6460 10240 6512 10260
rect 6512 10240 6514 10260
rect 6366 9832 6422 9888
rect 6182 9424 6238 9480
rect 6182 9152 6238 9208
rect 6182 8880 6238 8936
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 6090 6724 6146 6760
rect 6090 6704 6092 6724
rect 6092 6704 6144 6724
rect 6144 6704 6146 6724
rect 6182 5752 6238 5808
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5722 5228 5778 5264
rect 5722 5208 5724 5228
rect 5724 5208 5776 5228
rect 5776 5208 5778 5228
rect 5170 3576 5226 3632
rect 4894 1400 4950 1456
rect 4066 176 4122 232
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 5998 2080 6054 2136
rect 6090 1264 6146 1320
rect 6366 4120 6422 4176
rect 6458 3576 6514 3632
rect 6734 21120 6790 21176
rect 6918 20168 6974 20224
rect 6734 20032 6790 20088
rect 6918 17992 6974 18048
rect 7194 20304 7250 20360
rect 7378 18808 7434 18864
rect 7378 18536 7434 18592
rect 7746 25064 7802 25120
rect 7470 18400 7526 18456
rect 7470 18028 7472 18048
rect 7472 18028 7524 18048
rect 7524 18028 7526 18048
rect 7470 17992 7526 18028
rect 6918 16904 6974 16960
rect 7194 16904 7250 16960
rect 7010 16632 7066 16688
rect 6734 15000 6790 15056
rect 7010 15272 7066 15328
rect 6918 14340 6974 14376
rect 6918 14320 6920 14340
rect 6920 14320 6972 14340
rect 6972 14320 6974 14340
rect 6734 13368 6790 13424
rect 6734 13096 6790 13152
rect 6734 12552 6790 12608
rect 6734 11600 6790 11656
rect 6826 11464 6882 11520
rect 4986 312 5042 368
rect 6274 448 6330 504
rect 6918 7928 6974 7984
rect 6826 6840 6882 6896
rect 7102 7420 7104 7440
rect 7104 7420 7156 7440
rect 7156 7420 7158 7440
rect 7102 7384 7158 7420
rect 7654 17176 7710 17232
rect 8022 23044 8078 23080
rect 8022 23024 8024 23044
rect 8024 23024 8076 23044
rect 8076 23024 8078 23044
rect 7838 20984 7894 21040
rect 7930 19780 7986 19816
rect 7930 19760 7932 19780
rect 7932 19760 7984 19780
rect 7984 19760 7986 19780
rect 7838 17992 7894 18048
rect 8482 22888 8538 22944
rect 8390 21120 8446 21176
rect 8206 20712 8262 20768
rect 8298 20052 8354 20088
rect 8298 20032 8300 20052
rect 8300 20032 8352 20052
rect 8352 20032 8354 20052
rect 8666 24012 8668 24032
rect 8668 24012 8720 24032
rect 8720 24012 8722 24032
rect 8666 23976 8722 24012
rect 8850 24520 8906 24576
rect 8758 21528 8814 21584
rect 9218 25336 9274 25392
rect 9126 24384 9182 24440
rect 9034 24112 9090 24168
rect 8666 18264 8722 18320
rect 8942 18400 8998 18456
rect 7562 15680 7618 15736
rect 7286 10804 7342 10840
rect 7286 10784 7288 10804
rect 7288 10784 7340 10804
rect 7340 10784 7342 10804
rect 7194 7248 7250 7304
rect 7194 6296 7250 6352
rect 6826 3068 6828 3088
rect 6828 3068 6880 3088
rect 6880 3068 6882 3088
rect 6826 3032 6882 3068
rect 7194 5480 7250 5536
rect 7746 15428 7802 15464
rect 7746 15408 7748 15428
rect 7748 15408 7800 15428
rect 7800 15408 7802 15428
rect 7746 15136 7802 15192
rect 7746 11192 7802 11248
rect 7654 10648 7710 10704
rect 7654 9988 7710 10024
rect 7654 9968 7656 9988
rect 7656 9968 7708 9988
rect 7708 9968 7710 9988
rect 7562 9696 7618 9752
rect 7654 9016 7710 9072
rect 7378 7268 7434 7304
rect 7378 7248 7380 7268
rect 7380 7248 7432 7268
rect 7432 7248 7434 7268
rect 7562 7520 7618 7576
rect 7470 5480 7526 5536
rect 7562 4664 7618 4720
rect 7562 3848 7618 3904
rect 7194 856 7250 912
rect 7470 584 7526 640
rect 8022 17040 8078 17096
rect 8022 16088 8078 16144
rect 8022 15408 8078 15464
rect 8574 17332 8630 17368
rect 8574 17312 8576 17332
rect 8576 17312 8628 17332
rect 8628 17312 8630 17332
rect 8482 16224 8538 16280
rect 8390 16088 8446 16144
rect 8574 15680 8630 15736
rect 8022 14320 8078 14376
rect 8206 14048 8262 14104
rect 8758 15680 8814 15736
rect 8942 17584 8998 17640
rect 9402 24928 9458 24984
rect 9494 24792 9550 24848
rect 9494 24384 9550 24440
rect 10046 26424 10102 26480
rect 9218 21120 9274 21176
rect 8666 15272 8722 15328
rect 8850 15272 8906 15328
rect 8574 14592 8630 14648
rect 8390 13776 8446 13832
rect 8390 12860 8392 12880
rect 8392 12860 8444 12880
rect 8444 12860 8446 12880
rect 8390 12824 8446 12860
rect 8298 12280 8354 12336
rect 8298 12008 8354 12064
rect 8022 11736 8078 11792
rect 8206 11736 8262 11792
rect 8206 11600 8262 11656
rect 8298 11192 8354 11248
rect 7930 10648 7986 10704
rect 8022 9560 8078 9616
rect 7930 7828 7932 7848
rect 7932 7828 7984 7848
rect 7984 7828 7986 7848
rect 7930 7792 7986 7828
rect 7930 6976 7986 7032
rect 9034 13912 9090 13968
rect 8942 13504 8998 13560
rect 9126 13812 9128 13832
rect 9128 13812 9180 13832
rect 9180 13812 9182 13832
rect 9126 13776 9182 13812
rect 9126 13640 9182 13696
rect 8666 12280 8722 12336
rect 8114 6452 8170 6488
rect 8114 6432 8116 6452
rect 8116 6432 8168 6452
rect 8168 6432 8170 6452
rect 8022 5208 8078 5264
rect 8022 3576 8078 3632
rect 7838 3460 7894 3496
rect 7838 3440 7840 3460
rect 7840 3440 7892 3460
rect 7892 3440 7894 3460
rect 8298 5752 8354 5808
rect 8298 3712 8354 3768
rect 7930 2796 7932 2816
rect 7932 2796 7984 2816
rect 7984 2796 7986 2816
rect 7930 2760 7986 2796
rect 8850 11736 8906 11792
rect 8574 7520 8630 7576
rect 9494 22924 9496 22944
rect 9496 22924 9548 22944
rect 9548 22924 9550 22944
rect 9494 22888 9550 22924
rect 9310 20848 9366 20904
rect 9310 20576 9366 20632
rect 9678 20168 9734 20224
rect 9494 19352 9550 19408
rect 9678 18828 9734 18864
rect 9678 18808 9680 18828
rect 9680 18808 9732 18828
rect 9732 18808 9734 18828
rect 9402 17176 9458 17232
rect 9678 17876 9734 17912
rect 9678 17856 9680 17876
rect 9680 17856 9732 17876
rect 9732 17856 9734 17876
rect 9402 15136 9458 15192
rect 9310 13912 9366 13968
rect 9678 13776 9734 13832
rect 8850 6976 8906 7032
rect 9218 7248 9274 7304
rect 8758 6160 8814 6216
rect 8850 5908 8906 5944
rect 8850 5888 8852 5908
rect 8852 5888 8904 5908
rect 8904 5888 8906 5908
rect 8574 4392 8630 4448
rect 8482 3848 8538 3904
rect 8942 4936 8998 4992
rect 8574 3304 8630 3360
rect 8574 2896 8630 2952
rect 8758 2896 8814 2952
rect 9218 4528 9274 4584
rect 9218 4256 9274 4312
rect 8942 3032 8998 3088
rect 9678 11464 9734 11520
rect 9586 11328 9642 11384
rect 9494 9560 9550 9616
rect 9402 8744 9458 8800
rect 9678 9444 9734 9480
rect 9678 9424 9680 9444
rect 9680 9424 9732 9444
rect 9732 9424 9734 9444
rect 9862 23160 9918 23216
rect 11334 26560 11390 26616
rect 11610 26560 11666 26616
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10138 24656 10194 24712
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10690 24112 10746 24168
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10782 23840 10838 23896
rect 11058 24828 11060 24848
rect 11060 24828 11112 24848
rect 11112 24828 11114 24848
rect 11058 24792 11114 24828
rect 11426 24792 11482 24848
rect 11426 24248 11482 24304
rect 10966 23976 11022 24032
rect 11334 23704 11390 23760
rect 10782 23024 10838 23080
rect 10690 22616 10746 22672
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10690 20984 10746 21040
rect 10138 20848 10194 20904
rect 10046 20712 10102 20768
rect 10046 20204 10048 20224
rect 10048 20204 10100 20224
rect 10100 20204 10102 20224
rect 10046 20168 10102 20204
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 9954 16360 10010 16416
rect 9862 15816 9918 15872
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10782 20576 10838 20632
rect 10690 18808 10746 18864
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10874 17876 10930 17912
rect 10874 17856 10876 17876
rect 10876 17856 10928 17876
rect 10928 17856 10930 17876
rect 11058 23180 11114 23216
rect 11058 23160 11060 23180
rect 11060 23160 11112 23180
rect 11112 23160 11114 23180
rect 11242 23024 11298 23080
rect 11150 22888 11206 22944
rect 11242 22752 11298 22808
rect 11058 20984 11114 21040
rect 11426 23160 11482 23216
rect 11610 24520 11666 24576
rect 11610 24248 11666 24304
rect 11610 23568 11666 23624
rect 11242 20576 11298 20632
rect 11058 17992 11114 18048
rect 11242 17856 11298 17912
rect 11242 17312 11298 17368
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 9954 13368 10010 13424
rect 10598 14456 10654 14512
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10230 13368 10286 13424
rect 10046 12824 10102 12880
rect 9678 8336 9734 8392
rect 9494 4800 9550 4856
rect 9494 3576 9550 3632
rect 8666 2488 8722 2544
rect 9218 2624 9274 2680
rect 9770 4392 9826 4448
rect 9678 4120 9734 4176
rect 9954 12008 10010 12064
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10138 11192 10194 11248
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10138 9832 10194 9888
rect 10598 9832 10654 9888
rect 10598 9696 10654 9752
rect 10598 9424 10654 9480
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 11242 16496 11298 16552
rect 10874 15000 10930 15056
rect 11334 15136 11390 15192
rect 10966 14592 11022 14648
rect 10966 13776 11022 13832
rect 10874 13504 10930 13560
rect 10782 12552 10838 12608
rect 10874 12300 10930 12336
rect 10874 12280 10876 12300
rect 10876 12280 10928 12300
rect 10928 12280 10930 12300
rect 11242 14356 11244 14376
rect 11244 14356 11296 14376
rect 11296 14356 11298 14376
rect 11242 14320 11298 14356
rect 11334 14184 11390 14240
rect 11886 23568 11942 23624
rect 12530 24384 12586 24440
rect 12438 23976 12494 24032
rect 12070 22752 12126 22808
rect 11702 22072 11758 22128
rect 11886 22072 11942 22128
rect 12070 20304 12126 20360
rect 11702 19796 11704 19816
rect 11704 19796 11756 19816
rect 11756 19796 11758 19816
rect 11702 19760 11758 19796
rect 11518 15408 11574 15464
rect 11242 13776 11298 13832
rect 11150 12960 11206 13016
rect 11150 12688 11206 12744
rect 10874 12144 10930 12200
rect 10874 11600 10930 11656
rect 10782 11328 10838 11384
rect 10782 11192 10838 11248
rect 10966 11056 11022 11112
rect 11058 10648 11114 10704
rect 10874 10412 10876 10432
rect 10876 10412 10928 10432
rect 10928 10412 10930 10432
rect 10874 10376 10930 10412
rect 11058 10240 11114 10296
rect 10966 9832 11022 9888
rect 10690 8200 10746 8256
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 11058 9152 11114 9208
rect 11058 8472 11114 8528
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10414 6704 10470 6760
rect 10598 6704 10654 6760
rect 9954 6452 10010 6488
rect 9954 6432 9956 6452
rect 9956 6432 10008 6452
rect 10008 6432 10010 6452
rect 9954 6160 10010 6216
rect 9586 3304 9642 3360
rect 9770 3304 9826 3360
rect 9770 2796 9772 2816
rect 9772 2796 9824 2816
rect 9824 2796 9826 2816
rect 9770 2760 9826 2796
rect 9586 2216 9642 2272
rect 9770 992 9826 1048
rect 10506 6432 10562 6488
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10322 5480 10378 5536
rect 10506 5480 10562 5536
rect 10966 7112 11022 7168
rect 11886 16496 11942 16552
rect 11794 15544 11850 15600
rect 11794 15272 11850 15328
rect 11702 13232 11758 13288
rect 11610 12688 11666 12744
rect 11518 12416 11574 12472
rect 11426 11872 11482 11928
rect 11426 11192 11482 11248
rect 11334 9988 11390 10024
rect 11334 9968 11336 9988
rect 11336 9968 11388 9988
rect 11388 9968 11390 9988
rect 10874 5072 10930 5128
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10322 4428 10324 4448
rect 10324 4428 10376 4448
rect 10376 4428 10378 4448
rect 10322 4392 10378 4428
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 11058 4256 11114 4312
rect 10782 3168 10838 3224
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10690 2624 10746 2680
rect 10598 2352 10654 2408
rect 10782 2352 10838 2408
rect 10966 1944 11022 2000
rect 11242 3032 11298 3088
rect 11058 1672 11114 1728
rect 10598 1128 10654 1184
rect 11242 2488 11298 2544
rect 11702 12280 11758 12336
rect 11610 10240 11666 10296
rect 11518 5208 11574 5264
rect 11610 4800 11666 4856
rect 11518 3984 11574 4040
rect 11242 1672 11298 1728
rect 11426 1128 11482 1184
rect 11978 14184 12034 14240
rect 11886 12280 11942 12336
rect 11886 10804 11942 10840
rect 11886 10784 11888 10804
rect 11888 10784 11940 10804
rect 11940 10784 11942 10804
rect 12438 23432 12494 23488
rect 12990 24656 13046 24712
rect 12806 22924 12808 22944
rect 12808 22924 12860 22944
rect 12860 22924 12862 22944
rect 12806 22888 12862 22924
rect 13358 24248 13414 24304
rect 13358 23704 13414 23760
rect 12990 22208 13046 22264
rect 12254 21528 12310 21584
rect 12714 21004 12770 21040
rect 12714 20984 12716 21004
rect 12716 20984 12768 21004
rect 12768 20984 12770 21004
rect 12990 20984 13046 21040
rect 12806 20848 12862 20904
rect 12898 20052 12954 20088
rect 12898 20032 12900 20052
rect 12900 20032 12952 20052
rect 12952 20032 12954 20052
rect 12162 17992 12218 18048
rect 12438 17992 12494 18048
rect 12438 17176 12494 17232
rect 13910 25472 13966 25528
rect 13910 24248 13966 24304
rect 14830 26288 14886 26344
rect 14462 26016 14518 26072
rect 14646 26016 14702 26072
rect 14462 25472 14518 25528
rect 14278 24792 14334 24848
rect 14646 25064 14702 25120
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15106 24792 15162 24848
rect 13634 21800 13690 21856
rect 13634 21140 13690 21176
rect 13634 21120 13636 21140
rect 13636 21120 13688 21140
rect 13688 21120 13690 21140
rect 14002 21972 14004 21992
rect 14004 21972 14056 21992
rect 14056 21972 14058 21992
rect 14002 21936 14058 21972
rect 13910 21120 13966 21176
rect 13910 20576 13966 20632
rect 13450 20032 13506 20088
rect 12346 16244 12402 16280
rect 12346 16224 12348 16244
rect 12348 16224 12400 16244
rect 12400 16224 12402 16244
rect 12162 15700 12218 15736
rect 12162 15680 12164 15700
rect 12164 15680 12216 15700
rect 12216 15680 12218 15700
rect 12070 13096 12126 13152
rect 12070 12552 12126 12608
rect 12070 12416 12126 12472
rect 11886 5788 11888 5808
rect 11888 5788 11940 5808
rect 11940 5788 11942 5808
rect 11886 5752 11942 5788
rect 12162 10104 12218 10160
rect 12622 14864 12678 14920
rect 12530 10920 12586 10976
rect 12530 10784 12586 10840
rect 12070 8472 12126 8528
rect 11794 3848 11850 3904
rect 11794 3440 11850 3496
rect 12438 9152 12494 9208
rect 12162 7520 12218 7576
rect 12070 4936 12126 4992
rect 12070 4120 12126 4176
rect 12438 7420 12440 7440
rect 12440 7420 12492 7440
rect 12492 7420 12494 7440
rect 12438 7384 12494 7420
rect 12530 6432 12586 6488
rect 12898 16088 12954 16144
rect 12898 14456 12954 14512
rect 13082 17312 13138 17368
rect 13174 16496 13230 16552
rect 12990 14320 13046 14376
rect 13542 16360 13598 16416
rect 13450 15816 13506 15872
rect 13450 15544 13506 15600
rect 13542 15444 13544 15464
rect 13544 15444 13596 15464
rect 13596 15444 13598 15464
rect 13542 15408 13598 15444
rect 14370 23976 14426 24032
rect 14278 23296 14334 23352
rect 14186 21664 14242 21720
rect 13910 16632 13966 16688
rect 13818 15680 13874 15736
rect 13726 15408 13782 15464
rect 13634 15136 13690 15192
rect 13358 14864 13414 14920
rect 13174 14320 13230 14376
rect 12714 11736 12770 11792
rect 12714 10648 12770 10704
rect 13174 13096 13230 13152
rect 13358 13096 13414 13152
rect 13174 12688 13230 12744
rect 13818 14592 13874 14648
rect 14278 20304 14334 20360
rect 14922 24676 14978 24712
rect 14922 24656 14924 24676
rect 14924 24656 14976 24676
rect 14976 24656 14978 24676
rect 15290 24656 15346 24712
rect 15382 24384 15438 24440
rect 14738 24112 14794 24168
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14738 22752 14794 22808
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15106 21256 15162 21312
rect 14830 20848 14886 20904
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14830 20168 14886 20224
rect 14738 19080 14794 19136
rect 14370 18128 14426 18184
rect 14186 17756 14188 17776
rect 14188 17756 14240 17776
rect 14240 17756 14242 17776
rect 14186 17720 14242 17756
rect 14370 17076 14372 17096
rect 14372 17076 14424 17096
rect 14424 17076 14426 17096
rect 14370 17040 14426 17076
rect 14370 16088 14426 16144
rect 14278 15952 14334 16008
rect 13818 13504 13874 13560
rect 14186 15272 14242 15328
rect 14002 13504 14058 13560
rect 14278 15136 14334 15192
rect 14554 17448 14610 17504
rect 14646 15408 14702 15464
rect 14370 14184 14426 14240
rect 14462 13776 14518 13832
rect 14370 13640 14426 13696
rect 13542 12960 13598 13016
rect 13082 11464 13138 11520
rect 12990 11192 13046 11248
rect 12898 9832 12954 9888
rect 12898 8472 12954 8528
rect 12806 5616 12862 5672
rect 12990 5616 13046 5672
rect 13450 11328 13506 11384
rect 13910 12144 13966 12200
rect 13634 11192 13690 11248
rect 13634 10920 13690 10976
rect 13542 10648 13598 10704
rect 13174 9016 13230 9072
rect 13818 10376 13874 10432
rect 13726 9016 13782 9072
rect 13726 8472 13782 8528
rect 13174 7112 13230 7168
rect 12530 3984 12586 4040
rect 12070 3304 12126 3360
rect 12254 3304 12310 3360
rect 11978 2080 12034 2136
rect 11886 720 11942 776
rect 13082 5072 13138 5128
rect 13358 6740 13360 6760
rect 13360 6740 13412 6760
rect 13412 6740 13414 6760
rect 13358 6704 13414 6740
rect 13266 5480 13322 5536
rect 13266 1808 13322 1864
rect 14002 9424 14058 9480
rect 15382 20576 15438 20632
rect 15382 20168 15438 20224
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15566 22480 15622 22536
rect 16118 23568 16174 23624
rect 15934 21936 15990 21992
rect 15842 20032 15898 20088
rect 15842 19624 15898 19680
rect 15842 19352 15898 19408
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 15106 18128 15162 18184
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14922 16768 14978 16824
rect 14830 16668 14832 16688
rect 14832 16668 14884 16688
rect 14884 16668 14886 16688
rect 14830 16632 14886 16668
rect 15106 16652 15162 16688
rect 15106 16632 15108 16652
rect 15108 16632 15160 16652
rect 15160 16632 15162 16652
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14922 15972 14978 16008
rect 14922 15952 14924 15972
rect 14924 15952 14976 15972
rect 14976 15952 14978 15972
rect 14922 15408 14978 15464
rect 15106 15444 15108 15464
rect 15108 15444 15160 15464
rect 15160 15444 15162 15464
rect 15106 15408 15162 15444
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14922 15000 14978 15056
rect 15658 18536 15714 18592
rect 15290 14356 15292 14376
rect 15292 14356 15344 14376
rect 15344 14356 15346 14376
rect 15290 14320 15346 14356
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14922 13268 14924 13288
rect 14924 13268 14976 13288
rect 14976 13268 14978 13288
rect 14922 13232 14978 13268
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14186 11600 14242 11656
rect 14278 11348 14334 11384
rect 14278 11328 14280 11348
rect 14280 11328 14332 11348
rect 14332 11328 14334 11348
rect 14186 10104 14242 10160
rect 14554 12416 14610 12472
rect 14554 12280 14610 12336
rect 14462 10784 14518 10840
rect 14462 10376 14518 10432
rect 14278 9288 14334 9344
rect 14094 8880 14150 8936
rect 13818 8200 13874 8256
rect 14002 7520 14058 7576
rect 13634 7248 13690 7304
rect 13726 5752 13782 5808
rect 14186 7112 14242 7168
rect 13910 5616 13966 5672
rect 14094 6296 14150 6352
rect 13634 2796 13636 2816
rect 13636 2796 13688 2816
rect 13688 2796 13690 2816
rect 13634 2760 13690 2796
rect 13542 2624 13598 2680
rect 13726 1808 13782 1864
rect 14094 4564 14096 4584
rect 14096 4564 14148 4584
rect 14148 4564 14150 4584
rect 14094 4528 14150 4564
rect 14278 6976 14334 7032
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 15382 12144 15438 12200
rect 14830 11328 14886 11384
rect 15290 11328 15346 11384
rect 14738 11092 14740 11112
rect 14740 11092 14792 11112
rect 14792 11092 14794 11112
rect 14738 11056 14794 11092
rect 14554 7248 14610 7304
rect 14738 6976 14794 7032
rect 14738 6432 14794 6488
rect 14278 4392 14334 4448
rect 14554 4528 14610 4584
rect 14554 4392 14610 4448
rect 14278 3576 14334 3632
rect 14646 4120 14702 4176
rect 14370 3440 14426 3496
rect 14002 2916 14058 2952
rect 14002 2896 14004 2916
rect 14004 2896 14056 2916
rect 14056 2896 14058 2916
rect 14554 3304 14610 3360
rect 14462 3168 14518 3224
rect 14554 3032 14610 3088
rect 14554 2352 14610 2408
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15290 10240 15346 10296
rect 15658 15272 15714 15328
rect 15842 17312 15898 17368
rect 15474 12008 15530 12064
rect 15474 11464 15530 11520
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14922 9288 14978 9344
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15658 10920 15714 10976
rect 15750 10648 15806 10704
rect 15658 10376 15714 10432
rect 15658 10240 15714 10296
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 16026 21664 16082 21720
rect 16026 21120 16082 21176
rect 16210 19488 16266 19544
rect 16210 18672 16266 18728
rect 16118 17856 16174 17912
rect 16026 15408 16082 15464
rect 15934 13132 15936 13152
rect 15936 13132 15988 13152
rect 15988 13132 15990 13152
rect 15934 13096 15990 13132
rect 17038 26288 17094 26344
rect 16946 24148 16948 24168
rect 16948 24148 17000 24168
rect 17000 24148 17002 24168
rect 16946 24112 17002 24148
rect 16578 23160 16634 23216
rect 16394 21120 16450 21176
rect 17222 25608 17278 25664
rect 17222 25200 17278 25256
rect 17130 24520 17186 24576
rect 17038 23840 17094 23896
rect 17222 23024 17278 23080
rect 16486 20576 16542 20632
rect 16394 20476 16396 20496
rect 16396 20476 16448 20496
rect 16448 20476 16450 20496
rect 16394 20440 16450 20476
rect 16394 20304 16450 20360
rect 16578 19508 16634 19544
rect 16578 19488 16580 19508
rect 16580 19488 16632 19508
rect 16632 19488 16634 19508
rect 16486 18028 16488 18048
rect 16488 18028 16540 18048
rect 16540 18028 16542 18048
rect 16486 17992 16542 18028
rect 17222 22344 17278 22400
rect 17038 22072 17094 22128
rect 17038 21292 17040 21312
rect 17040 21292 17092 21312
rect 17092 21292 17094 21312
rect 17038 21256 17094 21292
rect 17038 20032 17094 20088
rect 16946 19252 16948 19272
rect 16948 19252 17000 19272
rect 17000 19252 17002 19272
rect 16946 19216 17002 19252
rect 17130 18672 17186 18728
rect 16670 17312 16726 17368
rect 16486 17196 16542 17232
rect 16486 17176 16488 17196
rect 16488 17176 16540 17196
rect 16540 17176 16542 17196
rect 16118 12980 16174 13016
rect 16118 12960 16120 12980
rect 16120 12960 16172 12980
rect 16172 12960 16174 12980
rect 16210 12688 16266 12744
rect 16118 12280 16174 12336
rect 16026 10784 16082 10840
rect 16026 10240 16082 10296
rect 16026 10104 16082 10160
rect 15750 9016 15806 9072
rect 15750 8628 15806 8664
rect 15750 8608 15752 8628
rect 15752 8608 15804 8628
rect 15804 8608 15806 8628
rect 16394 11872 16450 11928
rect 16210 11736 16266 11792
rect 16210 10548 16212 10568
rect 16212 10548 16264 10568
rect 16264 10548 16266 10568
rect 16210 10512 16266 10548
rect 16210 10376 16266 10432
rect 16394 9968 16450 10024
rect 16302 9016 16358 9072
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15474 6060 15476 6080
rect 15476 6060 15528 6080
rect 15528 6060 15530 6080
rect 15474 6024 15530 6060
rect 15290 5908 15346 5944
rect 15290 5888 15292 5908
rect 15292 5888 15344 5908
rect 15344 5888 15346 5908
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15290 4664 15346 4720
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15014 4156 15016 4176
rect 15016 4156 15068 4176
rect 15068 4156 15070 4176
rect 15014 4120 15070 4156
rect 15658 4664 15714 4720
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15750 3984 15806 4040
rect 16210 8492 16266 8528
rect 16210 8472 16212 8492
rect 16212 8472 16264 8492
rect 16264 8472 16266 8492
rect 16578 12300 16634 12336
rect 16578 12280 16580 12300
rect 16580 12280 16632 12300
rect 16632 12280 16634 12300
rect 17314 22072 17370 22128
rect 17498 23704 17554 23760
rect 17774 23296 17830 23352
rect 17682 23160 17738 23216
rect 17498 22888 17554 22944
rect 17682 21800 17738 21856
rect 17682 20848 17738 20904
rect 18234 23432 18290 23488
rect 18234 22208 18290 22264
rect 17774 19116 17776 19136
rect 17776 19116 17828 19136
rect 17828 19116 17830 19136
rect 17774 19080 17830 19116
rect 16854 14864 16910 14920
rect 16670 12180 16672 12200
rect 16672 12180 16724 12200
rect 16724 12180 16726 12200
rect 16670 12144 16726 12180
rect 16762 11328 16818 11384
rect 16762 10532 16818 10568
rect 16762 10512 16764 10532
rect 16764 10512 16816 10532
rect 16816 10512 16818 10532
rect 17958 17584 18014 17640
rect 18234 21256 18290 21312
rect 18142 21120 18198 21176
rect 18694 23432 18750 23488
rect 18418 23024 18474 23080
rect 18326 18300 18328 18320
rect 18328 18300 18380 18320
rect 18380 18300 18382 18320
rect 18326 18264 18382 18300
rect 18234 17876 18290 17912
rect 18234 17856 18236 17876
rect 18236 17856 18288 17876
rect 18288 17856 18290 17876
rect 18142 17584 18198 17640
rect 17774 16904 17830 16960
rect 17406 14184 17462 14240
rect 17314 13404 17316 13424
rect 17316 13404 17368 13424
rect 17368 13404 17370 13424
rect 17314 13368 17370 13404
rect 17498 13252 17554 13288
rect 17498 13232 17500 13252
rect 17500 13232 17552 13252
rect 17552 13232 17554 13252
rect 17498 12860 17500 12880
rect 17500 12860 17552 12880
rect 17552 12860 17554 12880
rect 17498 12824 17554 12860
rect 17130 11056 17186 11112
rect 16946 10240 17002 10296
rect 16854 9868 16856 9888
rect 16856 9868 16908 9888
rect 16908 9868 16910 9888
rect 16854 9832 16910 9868
rect 15382 3712 15438 3768
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15106 1572 15108 1592
rect 15108 1572 15160 1592
rect 15160 1572 15162 1592
rect 15106 1536 15162 1572
rect 15198 1264 15254 1320
rect 14830 212 14832 232
rect 14832 212 14884 232
rect 14884 212 14886 232
rect 14830 176 14886 212
rect 15842 3032 15898 3088
rect 16854 6976 16910 7032
rect 16578 6296 16634 6352
rect 16762 6568 16818 6624
rect 16302 3732 16358 3768
rect 16302 3712 16304 3732
rect 16304 3712 16356 3732
rect 16356 3712 16358 3732
rect 16210 3168 16266 3224
rect 16762 3848 16818 3904
rect 17130 4664 17186 4720
rect 17314 8608 17370 8664
rect 17314 8336 17370 8392
rect 17498 8744 17554 8800
rect 16854 1808 16910 1864
rect 17038 584 17094 640
rect 15198 312 15254 368
rect 17406 2896 17462 2952
rect 17866 16124 17868 16144
rect 17868 16124 17920 16144
rect 17920 16124 17922 16144
rect 17866 16088 17922 16124
rect 18142 16360 18198 16416
rect 17958 14048 18014 14104
rect 18234 15428 18290 15464
rect 18234 15408 18236 15428
rect 18236 15408 18288 15428
rect 18288 15408 18290 15428
rect 18510 22752 18566 22808
rect 18602 22208 18658 22264
rect 18970 22208 19026 22264
rect 18786 20032 18842 20088
rect 18510 18808 18566 18864
rect 18602 18128 18658 18184
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19329 25336 19385 25392
rect 19154 24248 19210 24304
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 20258 25744 20314 25800
rect 20258 25472 20314 25528
rect 20350 25336 20406 25392
rect 20534 25744 20590 25800
rect 20534 24792 20590 24848
rect 20074 23840 20130 23896
rect 19246 22344 19302 22400
rect 19982 23568 20038 23624
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19430 22480 19486 22536
rect 19798 22516 19800 22536
rect 19800 22516 19852 22536
rect 19852 22516 19854 22536
rect 19798 22480 19854 22516
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19154 20032 19210 20088
rect 20442 23024 20498 23080
rect 19798 21800 19854 21856
rect 19706 21684 19762 21720
rect 19706 21664 19708 21684
rect 19708 21664 19760 21684
rect 19760 21664 19762 21684
rect 19890 21664 19946 21720
rect 19329 19780 19385 19816
rect 19329 19760 19340 19780
rect 19340 19760 19385 19780
rect 19062 18400 19118 18456
rect 18878 17720 18934 17776
rect 18694 17448 18750 17504
rect 18970 16360 19026 16416
rect 18510 15272 18566 15328
rect 18694 14592 18750 14648
rect 18602 14456 18658 14512
rect 18510 13640 18566 13696
rect 18510 12824 18566 12880
rect 18234 12416 18290 12472
rect 18050 11600 18106 11656
rect 17958 11192 18014 11248
rect 17866 10376 17922 10432
rect 18326 11192 18382 11248
rect 18050 9968 18106 10024
rect 17958 6860 18014 6896
rect 17958 6840 17960 6860
rect 17960 6840 18012 6860
rect 18012 6840 18014 6860
rect 18050 6432 18106 6488
rect 17682 4528 17738 4584
rect 17866 4528 17922 4584
rect 17314 2488 17370 2544
rect 17498 2488 17554 2544
rect 17314 2216 17370 2272
rect 17314 1128 17370 1184
rect 17498 1844 17500 1864
rect 17500 1844 17552 1864
rect 17552 1844 17554 1864
rect 17498 1808 17554 1844
rect 17406 856 17462 912
rect 17314 720 17370 776
rect 18050 3712 18106 3768
rect 17774 3612 17776 3632
rect 17776 3612 17828 3632
rect 17828 3612 17830 3632
rect 17774 3576 17830 3612
rect 18418 9696 18474 9752
rect 18326 8608 18382 8664
rect 18234 6316 18290 6352
rect 18234 6296 18236 6316
rect 18236 6296 18288 6316
rect 18288 6296 18290 6316
rect 18234 5636 18290 5672
rect 18234 5616 18236 5636
rect 18236 5616 18288 5636
rect 18288 5616 18290 5636
rect 18418 6976 18474 7032
rect 18418 5888 18474 5944
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19982 20440 20038 20496
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19246 16788 19302 16824
rect 19246 16768 19248 16788
rect 19248 16768 19300 16788
rect 19300 16768 19302 16788
rect 19430 16904 19486 16960
rect 19062 15272 19118 15328
rect 19430 15816 19486 15872
rect 18786 12960 18842 13016
rect 18878 12552 18934 12608
rect 19062 12416 19118 12472
rect 18786 11464 18842 11520
rect 18970 10804 19026 10840
rect 18970 10784 18972 10804
rect 18972 10784 19024 10804
rect 19024 10784 19026 10804
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 20074 19080 20130 19136
rect 20074 18536 20130 18592
rect 19982 17040 20038 17096
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19614 16652 19670 16688
rect 19614 16632 19616 16652
rect 19616 16632 19668 16652
rect 19668 16632 19670 16652
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19522 15136 19578 15192
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 20074 13676 20076 13696
rect 20076 13676 20128 13696
rect 20128 13676 20130 13696
rect 20074 13640 20130 13676
rect 19338 12436 19394 12472
rect 19338 12416 19340 12436
rect 19340 12416 19392 12436
rect 19392 12416 19394 12436
rect 19246 11464 19302 11520
rect 18878 10104 18934 10160
rect 19062 10104 19118 10160
rect 18786 9172 18842 9208
rect 18786 9152 18788 9172
rect 18788 9152 18840 9172
rect 18840 9152 18842 9172
rect 18786 8744 18842 8800
rect 18510 4256 18566 4312
rect 18142 3440 18198 3496
rect 18050 2796 18052 2816
rect 18052 2796 18104 2816
rect 18104 2796 18106 2816
rect 18050 2760 18106 2796
rect 19154 9424 19210 9480
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19982 12008 20038 12064
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19522 11056 19578 11112
rect 19430 10260 19486 10296
rect 19430 10240 19432 10260
rect 19432 10240 19484 10260
rect 19484 10240 19486 10260
rect 19430 9288 19486 9344
rect 19430 8880 19486 8936
rect 19154 6976 19210 7032
rect 19062 6160 19118 6216
rect 19430 7656 19486 7712
rect 19338 7112 19394 7168
rect 19430 6976 19486 7032
rect 19798 10956 19800 10976
rect 19800 10956 19852 10976
rect 19852 10956 19854 10976
rect 19798 10920 19854 10956
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19614 8900 19670 8936
rect 19614 8880 19616 8900
rect 19616 8880 19668 8900
rect 19668 8880 19670 8900
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19890 7812 19946 7848
rect 19890 7792 19892 7812
rect 19892 7792 19944 7812
rect 19944 7792 19946 7812
rect 19982 7384 20038 7440
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 18418 3168 18474 3224
rect 18602 3168 18658 3224
rect 18510 3032 18566 3088
rect 17038 176 17094 232
rect 18326 1400 18382 1456
rect 18694 1944 18750 2000
rect 18234 1264 18290 1320
rect 18418 1264 18474 1320
rect 19154 4800 19210 4856
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19522 4392 19578 4448
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19982 3340 19984 3360
rect 19984 3340 20036 3360
rect 20036 3340 20038 3360
rect 19982 3304 20038 3340
rect 20258 19508 20314 19544
rect 20258 19488 20260 19508
rect 20260 19488 20312 19508
rect 20312 19488 20314 19508
rect 20718 22652 20720 22672
rect 20720 22652 20772 22672
rect 20772 22652 20774 22672
rect 20718 22616 20774 22652
rect 20626 21528 20682 21584
rect 20718 21392 20774 21448
rect 20718 21120 20774 21176
rect 21086 24656 21142 24712
rect 20994 23296 21050 23352
rect 20994 23024 21050 23080
rect 20718 20576 20774 20632
rect 20534 19488 20590 19544
rect 20442 18572 20444 18592
rect 20444 18572 20496 18592
rect 20496 18572 20498 18592
rect 20442 18536 20498 18572
rect 20350 17448 20406 17504
rect 20258 14884 20314 14920
rect 20258 14864 20260 14884
rect 20260 14864 20312 14884
rect 20312 14864 20314 14884
rect 21822 24792 21878 24848
rect 21178 23024 21234 23080
rect 21178 22480 21234 22536
rect 21546 21800 21602 21856
rect 21546 21120 21602 21176
rect 20902 18808 20958 18864
rect 21086 18808 21142 18864
rect 20902 16360 20958 16416
rect 20902 14456 20958 14512
rect 21638 20168 21694 20224
rect 21546 19352 21602 19408
rect 21178 17448 21234 17504
rect 21730 19216 21786 19272
rect 21454 18536 21510 18592
rect 21638 18420 21694 18456
rect 21638 18400 21640 18420
rect 21640 18400 21692 18420
rect 21692 18400 21694 18420
rect 21546 17856 21602 17912
rect 21362 17176 21418 17232
rect 21270 16788 21326 16824
rect 21270 16768 21272 16788
rect 21272 16768 21324 16788
rect 21324 16768 21326 16788
rect 21178 14728 21234 14784
rect 20626 14048 20682 14104
rect 20258 12552 20314 12608
rect 20350 12008 20406 12064
rect 20350 10784 20406 10840
rect 20166 8744 20222 8800
rect 20258 8064 20314 8120
rect 20166 7792 20222 7848
rect 20626 13776 20682 13832
rect 20810 14184 20866 14240
rect 20718 13640 20774 13696
rect 20626 13232 20682 13288
rect 20442 10240 20498 10296
rect 20810 13132 20812 13152
rect 20812 13132 20864 13152
rect 20864 13132 20866 13152
rect 20810 13096 20866 13132
rect 20994 13096 21050 13152
rect 20718 12416 20774 12472
rect 20718 11736 20774 11792
rect 20718 11348 20774 11384
rect 20718 11328 20720 11348
rect 20720 11328 20772 11348
rect 20772 11328 20774 11348
rect 20994 12552 21050 12608
rect 20902 11464 20958 11520
rect 20718 9696 20774 9752
rect 20534 9288 20590 9344
rect 20258 5772 20314 5808
rect 20258 5752 20260 5772
rect 20260 5752 20312 5772
rect 20312 5752 20314 5772
rect 20166 4936 20222 4992
rect 20258 4800 20314 4856
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 19430 2624 19486 2680
rect 20074 2624 20130 2680
rect 19338 1400 19394 1456
rect 19430 312 19486 368
rect 20534 6568 20590 6624
rect 20902 8880 20958 8936
rect 21454 16088 21510 16144
rect 21546 12552 21602 12608
rect 21454 12416 21510 12472
rect 20994 8608 21050 8664
rect 20902 7928 20958 7984
rect 20718 7248 20774 7304
rect 20902 6976 20958 7032
rect 20810 6840 20866 6896
rect 20902 6724 20958 6760
rect 20902 6704 20904 6724
rect 20904 6704 20956 6724
rect 20956 6704 20958 6724
rect 21270 11872 21326 11928
rect 21270 11600 21326 11656
rect 21454 11872 21510 11928
rect 21362 11056 21418 11112
rect 22282 23196 22284 23216
rect 22284 23196 22336 23216
rect 22336 23196 22338 23216
rect 22282 23160 22338 23196
rect 22558 23704 22614 23760
rect 22190 21664 22246 21720
rect 22098 20984 22154 21040
rect 21914 17740 21970 17776
rect 21914 17720 21916 17740
rect 21916 17720 21968 17740
rect 21968 17720 21970 17740
rect 22190 17992 22246 18048
rect 22190 17040 22246 17096
rect 22098 16904 22154 16960
rect 22006 16088 22062 16144
rect 22006 15680 22062 15736
rect 21730 12708 21786 12744
rect 21730 12688 21732 12708
rect 21732 12688 21784 12708
rect 21784 12688 21786 12708
rect 21822 12552 21878 12608
rect 21730 12008 21786 12064
rect 21822 11192 21878 11248
rect 21822 10648 21878 10704
rect 21546 10104 21602 10160
rect 21454 9560 21510 9616
rect 21270 9152 21326 9208
rect 21178 9016 21234 9072
rect 21178 8608 21234 8664
rect 21362 9052 21364 9072
rect 21364 9052 21416 9072
rect 21416 9052 21418 9072
rect 21362 9016 21418 9052
rect 21730 10376 21786 10432
rect 21638 9696 21694 9752
rect 21822 10104 21878 10160
rect 22098 15408 22154 15464
rect 22098 15272 22154 15328
rect 22190 14592 22246 14648
rect 22006 13776 22062 13832
rect 22650 23468 22652 23488
rect 22652 23468 22704 23488
rect 22704 23468 22706 23488
rect 22650 23432 22706 23468
rect 22834 23024 22890 23080
rect 22742 20032 22798 20088
rect 22742 19352 22798 19408
rect 22374 19080 22430 19136
rect 22466 18672 22522 18728
rect 22650 16632 22706 16688
rect 22650 16224 22706 16280
rect 22374 13776 22430 13832
rect 22282 13132 22284 13152
rect 22284 13132 22336 13152
rect 22336 13132 22338 13152
rect 22282 13096 22338 13132
rect 22374 12860 22376 12880
rect 22376 12860 22428 12880
rect 22428 12860 22430 12880
rect 22374 12824 22430 12860
rect 22374 11872 22430 11928
rect 22190 11328 22246 11384
rect 21822 9560 21878 9616
rect 21178 8200 21234 8256
rect 21362 7520 21418 7576
rect 21546 7384 21602 7440
rect 21822 8336 21878 8392
rect 21822 7248 21878 7304
rect 21638 7112 21694 7168
rect 21178 6740 21180 6760
rect 21180 6740 21232 6760
rect 21232 6740 21234 6760
rect 21178 6704 21234 6740
rect 21178 6432 21234 6488
rect 20810 6024 20866 6080
rect 20718 5072 20774 5128
rect 20718 3984 20774 4040
rect 20626 3712 20682 3768
rect 20994 5364 21050 5400
rect 20994 5344 20996 5364
rect 20996 5344 21048 5364
rect 21048 5344 21050 5364
rect 20994 3440 21050 3496
rect 20994 3168 21050 3224
rect 21454 6840 21510 6896
rect 21270 6160 21326 6216
rect 21270 5888 21326 5944
rect 21362 5752 21418 5808
rect 21546 6296 21602 6352
rect 21730 6160 21786 6216
rect 21638 5072 21694 5128
rect 21822 5616 21878 5672
rect 23202 25880 23258 25936
rect 23110 25200 23166 25256
rect 23018 24112 23074 24168
rect 22650 14456 22706 14512
rect 22742 12980 22798 13016
rect 22742 12960 22744 12980
rect 22744 12960 22796 12980
rect 22796 12960 22798 12980
rect 22650 12688 22706 12744
rect 23754 26560 23810 26616
rect 23570 24792 23626 24848
rect 23478 22616 23534 22672
rect 23018 18672 23074 18728
rect 23018 16904 23074 16960
rect 22282 10648 22338 10704
rect 22190 8492 22246 8528
rect 22190 8472 22192 8492
rect 22192 8472 22244 8492
rect 22244 8472 22246 8492
rect 22466 10512 22522 10568
rect 22006 6024 22062 6080
rect 22282 6604 22284 6624
rect 22284 6604 22336 6624
rect 22336 6604 22338 6624
rect 22282 6568 22338 6604
rect 22098 5344 22154 5400
rect 21270 4684 21326 4720
rect 21270 4664 21272 4684
rect 21272 4664 21324 4684
rect 21324 4664 21326 4684
rect 21178 4392 21234 4448
rect 21362 3848 21418 3904
rect 21270 3304 21326 3360
rect 21178 3168 21234 3224
rect 20718 2916 20774 2952
rect 20718 2896 20720 2916
rect 20720 2896 20772 2916
rect 20772 2896 20774 2916
rect 21086 2896 21142 2952
rect 20534 2372 20590 2408
rect 20534 2352 20536 2372
rect 20536 2352 20588 2372
rect 20588 2352 20590 2372
rect 20902 2252 20904 2272
rect 20904 2252 20956 2272
rect 20956 2252 20958 2272
rect 20902 2216 20958 2252
rect 20994 1944 21050 2000
rect 21546 3712 21602 3768
rect 22190 5072 22246 5128
rect 21914 2488 21970 2544
rect 22926 10140 22928 10160
rect 22928 10140 22980 10160
rect 22980 10140 22982 10160
rect 22926 10104 22982 10140
rect 22926 9596 22928 9616
rect 22928 9596 22980 9616
rect 22980 9596 22982 9616
rect 22926 9560 22982 9596
rect 23110 12552 23166 12608
rect 23386 19624 23442 19680
rect 23662 23704 23718 23760
rect 23662 23432 23718 23488
rect 23662 22888 23718 22944
rect 24030 24656 24086 24712
rect 24766 27104 24822 27160
rect 24766 25336 24822 25392
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24674 24404 24730 24440
rect 24674 24384 24676 24404
rect 24676 24384 24728 24404
rect 24728 24384 24730 24404
rect 24398 24248 24454 24304
rect 23846 23704 23902 23760
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24766 23860 24822 23896
rect 24766 23840 24768 23860
rect 24768 23840 24820 23860
rect 24820 23840 24822 23860
rect 23754 22208 23810 22264
rect 24766 23432 24822 23488
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 23846 21936 23902 21992
rect 23570 18808 23626 18864
rect 23570 18672 23626 18728
rect 23662 18536 23718 18592
rect 23662 17584 23718 17640
rect 23478 17332 23534 17368
rect 23478 17312 23480 17332
rect 23480 17312 23532 17332
rect 23532 17312 23534 17332
rect 23478 14900 23480 14920
rect 23480 14900 23532 14920
rect 23532 14900 23534 14920
rect 23478 14864 23534 14900
rect 23386 14592 23442 14648
rect 23386 13504 23442 13560
rect 23386 12436 23442 12472
rect 23386 12416 23388 12436
rect 23388 12416 23440 12436
rect 23440 12416 23442 12436
rect 23570 12552 23626 12608
rect 23570 12144 23626 12200
rect 22742 8472 22798 8528
rect 22926 8336 22982 8392
rect 22834 7928 22890 7984
rect 22926 6976 22982 7032
rect 22650 6840 22706 6896
rect 22466 4528 22522 4584
rect 23018 5208 23074 5264
rect 23294 10004 23296 10024
rect 23296 10004 23348 10024
rect 23348 10004 23350 10024
rect 23294 9968 23350 10004
rect 23478 11092 23480 11112
rect 23480 11092 23532 11112
rect 23532 11092 23534 11112
rect 23478 11056 23534 11092
rect 23570 10648 23626 10704
rect 23478 10104 23534 10160
rect 24030 21836 24032 21856
rect 24032 21836 24084 21856
rect 24084 21836 24086 21856
rect 24030 21800 24086 21836
rect 23938 21664 23994 21720
rect 23938 21528 23994 21584
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24214 21256 24270 21312
rect 24030 20748 24032 20768
rect 24032 20748 24084 20768
rect 24084 20748 24086 20768
rect 24030 20712 24086 20748
rect 24582 21292 24584 21312
rect 24584 21292 24636 21312
rect 24636 21292 24638 21312
rect 24582 21256 24638 21292
rect 24950 22072 25006 22128
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24490 19352 24546 19408
rect 24030 18536 24086 18592
rect 24490 18672 24546 18728
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24030 18128 24086 18184
rect 24030 15700 24086 15736
rect 24030 15680 24032 15700
rect 24032 15680 24084 15700
rect 24084 15680 24086 15700
rect 24950 18300 24952 18320
rect 24952 18300 25004 18320
rect 25004 18300 25006 18320
rect 24950 18264 25006 18300
rect 24766 18128 24822 18184
rect 24766 17720 24822 17776
rect 25226 24792 25282 24848
rect 25778 26152 25834 26208
rect 26146 25744 26202 25800
rect 25870 24656 25926 24712
rect 25318 23704 25374 23760
rect 25226 23296 25282 23352
rect 25134 22480 25190 22536
rect 25226 21256 25282 21312
rect 25134 19760 25190 19816
rect 25226 18400 25282 18456
rect 25134 17856 25190 17912
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 23938 15272 23994 15328
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24858 17176 24914 17232
rect 25042 16788 25098 16824
rect 25042 16768 25044 16788
rect 25044 16768 25096 16788
rect 25096 16768 25098 16788
rect 24766 14864 24822 14920
rect 24674 13504 24730 13560
rect 24214 13232 24270 13288
rect 23938 12008 23994 12064
rect 23754 10512 23810 10568
rect 23294 9832 23350 9888
rect 23570 9968 23626 10024
rect 23662 9560 23718 9616
rect 23570 9424 23626 9480
rect 22650 4528 22706 4584
rect 22650 4392 22706 4448
rect 22466 4120 22522 4176
rect 22282 2644 22338 2680
rect 22282 2624 22284 2644
rect 22284 2624 22336 2644
rect 22336 2624 22338 2644
rect 22742 4120 22798 4176
rect 22742 2352 22798 2408
rect 23110 2624 23166 2680
rect 22834 1672 22890 1728
rect 22926 1400 22982 1456
rect 23478 9288 23534 9344
rect 23478 9016 23534 9072
rect 23754 9016 23810 9072
rect 23662 8780 23664 8800
rect 23664 8780 23716 8800
rect 23716 8780 23718 8800
rect 23662 8744 23718 8780
rect 23478 8336 23534 8392
rect 23662 8200 23718 8256
rect 23662 7928 23718 7984
rect 23294 7656 23350 7712
rect 23478 7384 23534 7440
rect 23478 7112 23534 7168
rect 23294 5616 23350 5672
rect 24030 11500 24032 11520
rect 24032 11500 24084 11520
rect 24084 11500 24086 11520
rect 24030 11464 24086 11500
rect 24030 9696 24086 9752
rect 23846 8744 23902 8800
rect 23938 8608 23994 8664
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24214 12552 24270 12608
rect 24858 13232 24914 13288
rect 24950 12416 25006 12472
rect 24858 12280 24914 12336
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24766 11872 24822 11928
rect 24674 11600 24730 11656
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 23662 5364 23718 5400
rect 23662 5344 23664 5364
rect 23664 5344 23716 5364
rect 23716 5344 23718 5364
rect 20166 40 20222 96
rect 23386 4120 23442 4176
rect 23478 3612 23480 3632
rect 23480 3612 23532 3632
rect 23532 3612 23534 3632
rect 24030 6704 24086 6760
rect 23938 6024 23994 6080
rect 24030 5344 24086 5400
rect 23846 4392 23902 4448
rect 23478 3576 23534 3612
rect 23846 3032 23902 3088
rect 23570 1400 23626 1456
rect 23386 720 23442 776
rect 24030 3168 24086 3224
rect 24030 2760 24086 2816
rect 23938 2216 23994 2272
rect 23938 1672 23994 1728
rect 24030 992 24086 1048
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24582 6160 24638 6216
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 25042 10920 25098 10976
rect 25042 9560 25098 9616
rect 24766 8336 24822 8392
rect 25410 23024 25466 23080
rect 25686 21800 25742 21856
rect 25502 20576 25558 20632
rect 25410 20032 25466 20088
rect 25502 18264 25558 18320
rect 25410 15680 25466 15736
rect 25318 15408 25374 15464
rect 25226 13812 25228 13832
rect 25228 13812 25280 13832
rect 25280 13812 25282 13832
rect 25226 13776 25282 13812
rect 25502 15580 25504 15600
rect 25504 15580 25556 15600
rect 25556 15580 25558 15600
rect 25502 15544 25558 15580
rect 24858 8064 24914 8120
rect 25042 8084 25098 8120
rect 25042 8064 25044 8084
rect 25044 8064 25096 8084
rect 25096 8064 25098 8084
rect 25410 13096 25466 13152
rect 25502 12688 25558 12744
rect 25778 19488 25834 19544
rect 25686 18944 25742 19000
rect 25962 20340 25964 20360
rect 25964 20340 26016 20360
rect 26016 20340 26018 20360
rect 25962 20304 26018 20340
rect 25962 17176 26018 17232
rect 25318 9968 25374 10024
rect 25042 6840 25098 6896
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24214 3848 24270 3904
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24490 2508 24546 2544
rect 24490 2488 24492 2508
rect 24492 2488 24544 2508
rect 24544 2488 24546 2508
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24674 1536 24730 1592
rect 24766 584 24822 640
rect 24950 4936 25006 4992
rect 25042 4700 25044 4720
rect 25044 4700 25096 4720
rect 25096 4700 25098 4720
rect 25042 4664 25098 4700
rect 24950 4140 25006 4176
rect 24950 4120 24952 4140
rect 24952 4120 25004 4140
rect 25004 4120 25006 4140
rect 25042 4020 25044 4040
rect 25044 4020 25096 4040
rect 25096 4020 25098 4040
rect 25042 3984 25098 4020
rect 25410 9560 25466 9616
rect 25594 12300 25650 12336
rect 25594 12280 25596 12300
rect 25596 12280 25648 12300
rect 25648 12280 25650 12300
rect 25594 10920 25650 10976
rect 25778 13912 25834 13968
rect 25778 13368 25834 13424
rect 25870 13232 25926 13288
rect 25778 10376 25834 10432
rect 25778 9424 25834 9480
rect 25686 6976 25742 7032
rect 25502 4936 25558 4992
rect 25410 4800 25466 4856
rect 25318 3984 25374 4040
rect 25226 3712 25282 3768
rect 25134 2896 25190 2952
rect 25410 3440 25466 3496
rect 25226 2760 25282 2816
rect 26514 24384 26570 24440
rect 25962 10512 26018 10568
rect 25962 9560 26018 9616
rect 26238 15988 26240 16008
rect 26240 15988 26292 16008
rect 26292 15988 26294 16008
rect 26238 15952 26294 15988
rect 26238 15036 26240 15056
rect 26240 15036 26292 15056
rect 26292 15036 26294 15056
rect 26238 15000 26294 15036
rect 26238 14356 26240 14376
rect 26240 14356 26292 14376
rect 26292 14356 26294 14376
rect 26238 14320 26294 14356
rect 26238 13640 26294 13696
rect 26238 11772 26240 11792
rect 26240 11772 26292 11792
rect 26292 11772 26294 11792
rect 26238 11736 26294 11772
rect 26238 9172 26294 9208
rect 26238 9152 26240 9172
rect 26240 9152 26292 9172
rect 26292 9152 26294 9172
rect 27618 23840 27674 23896
rect 27066 23432 27122 23488
rect 26422 8880 26478 8936
rect 26054 7828 26056 7848
rect 26056 7828 26108 7848
rect 26108 7828 26110 7848
rect 26054 7792 26110 7828
rect 26422 7148 26424 7168
rect 26424 7148 26476 7168
rect 26476 7148 26478 7168
rect 25778 1808 25834 1864
rect 25042 1264 25098 1320
rect 26422 7112 26478 7148
rect 26238 5888 26294 5944
rect 26238 5788 26240 5808
rect 26240 5788 26292 5808
rect 26292 5788 26294 5808
rect 26238 5752 26294 5788
rect 27066 3984 27122 4040
rect 26514 3848 26570 3904
rect 26238 3052 26294 3088
rect 26238 3032 26240 3052
rect 26240 3032 26292 3052
rect 26292 3032 26294 3052
rect 26422 2508 26478 2544
rect 26422 2488 26424 2508
rect 26424 2488 26476 2508
rect 26476 2488 26478 2508
rect 26146 1672 26202 1728
rect 23294 312 23350 368
rect 26054 448 26110 504
rect 27618 3440 27674 3496
<< metal3 >>
rect 0 27706 480 27736
rect 1117 27706 1183 27709
rect 0 27704 1183 27706
rect 0 27648 1122 27704
rect 1178 27648 1183 27704
rect 0 27646 1183 27648
rect 0 27616 480 27646
rect 1117 27643 1183 27646
rect 23749 27706 23815 27709
rect 27520 27706 28000 27736
rect 23749 27704 28000 27706
rect 23749 27648 23754 27704
rect 23810 27648 28000 27704
rect 23749 27646 28000 27648
rect 23749 27643 23815 27646
rect 27520 27616 28000 27646
rect 0 27162 480 27192
rect 657 27162 723 27165
rect 0 27160 723 27162
rect 0 27104 662 27160
rect 718 27104 723 27160
rect 0 27102 723 27104
rect 0 27072 480 27102
rect 657 27099 723 27102
rect 24761 27162 24827 27165
rect 27520 27162 28000 27192
rect 24761 27160 28000 27162
rect 24761 27104 24766 27160
rect 24822 27104 28000 27160
rect 24761 27102 28000 27104
rect 24761 27099 24827 27102
rect 27520 27072 28000 27102
rect 0 26618 480 26648
rect 1301 26618 1367 26621
rect 0 26616 1367 26618
rect 0 26560 1306 26616
rect 1362 26560 1367 26616
rect 0 26558 1367 26560
rect 0 26528 480 26558
rect 1301 26555 1367 26558
rect 11329 26618 11395 26621
rect 11605 26618 11671 26621
rect 21950 26618 21956 26620
rect 11329 26616 21956 26618
rect 11329 26560 11334 26616
rect 11390 26560 11610 26616
rect 11666 26560 21956 26616
rect 11329 26558 21956 26560
rect 11329 26555 11395 26558
rect 11605 26555 11671 26558
rect 21950 26556 21956 26558
rect 22020 26556 22026 26620
rect 23749 26618 23815 26621
rect 27520 26618 28000 26648
rect 23749 26616 28000 26618
rect 23749 26560 23754 26616
rect 23810 26560 28000 26616
rect 23749 26558 28000 26560
rect 23749 26555 23815 26558
rect 27520 26528 28000 26558
rect 10041 26482 10107 26485
rect 21030 26482 21036 26484
rect 10041 26480 21036 26482
rect 10041 26424 10046 26480
rect 10102 26424 21036 26480
rect 10041 26422 21036 26424
rect 10041 26419 10107 26422
rect 21030 26420 21036 26422
rect 21100 26420 21106 26484
rect 12934 26284 12940 26348
rect 13004 26346 13010 26348
rect 14825 26346 14891 26349
rect 13004 26344 14891 26346
rect 13004 26288 14830 26344
rect 14886 26288 14891 26344
rect 13004 26286 14891 26288
rect 13004 26284 13010 26286
rect 14825 26283 14891 26286
rect 17033 26346 17099 26349
rect 23606 26346 23612 26348
rect 17033 26344 23612 26346
rect 17033 26288 17038 26344
rect 17094 26288 23612 26344
rect 17033 26286 23612 26288
rect 17033 26283 17099 26286
rect 23606 26284 23612 26286
rect 23676 26284 23682 26348
rect 2998 26148 3004 26212
rect 3068 26210 3074 26212
rect 25773 26210 25839 26213
rect 3068 26208 25839 26210
rect 3068 26152 25778 26208
rect 25834 26152 25839 26208
rect 3068 26150 25839 26152
rect 3068 26148 3074 26150
rect 25773 26147 25839 26150
rect 6361 26074 6427 26077
rect 14457 26074 14523 26077
rect 6361 26072 14523 26074
rect 6361 26016 6366 26072
rect 6422 26016 14462 26072
rect 14518 26016 14523 26072
rect 6361 26014 14523 26016
rect 6361 26011 6427 26014
rect 14457 26011 14523 26014
rect 14641 26074 14707 26077
rect 25078 26074 25084 26076
rect 14641 26072 25084 26074
rect 14641 26016 14646 26072
rect 14702 26016 25084 26072
rect 14641 26014 25084 26016
rect 14641 26011 14707 26014
rect 25078 26012 25084 26014
rect 25148 26012 25154 26076
rect 0 25938 480 25968
rect 1025 25938 1091 25941
rect 0 25936 1091 25938
rect 0 25880 1030 25936
rect 1086 25880 1091 25936
rect 0 25878 1091 25880
rect 0 25848 480 25878
rect 1025 25875 1091 25878
rect 3734 25876 3740 25940
rect 3804 25938 3810 25940
rect 22318 25938 22324 25940
rect 3804 25878 22324 25938
rect 3804 25876 3810 25878
rect 22318 25876 22324 25878
rect 22388 25876 22394 25940
rect 23197 25938 23263 25941
rect 27520 25938 28000 25968
rect 23197 25936 28000 25938
rect 23197 25880 23202 25936
rect 23258 25880 28000 25936
rect 23197 25878 28000 25880
rect 23197 25875 23263 25878
rect 27520 25848 28000 25878
rect 2446 25740 2452 25804
rect 2516 25802 2522 25804
rect 20253 25802 20319 25805
rect 2516 25800 20319 25802
rect 2516 25744 20258 25800
rect 20314 25744 20319 25800
rect 2516 25742 20319 25744
rect 2516 25740 2522 25742
rect 20253 25739 20319 25742
rect 20529 25802 20595 25805
rect 26141 25802 26207 25805
rect 20529 25800 26207 25802
rect 20529 25744 20534 25800
rect 20590 25744 26146 25800
rect 26202 25744 26207 25800
rect 20529 25742 26207 25744
rect 20529 25739 20595 25742
rect 26141 25739 26207 25742
rect 12198 25604 12204 25668
rect 12268 25666 12274 25668
rect 17217 25666 17283 25669
rect 12268 25664 17283 25666
rect 12268 25608 17222 25664
rect 17278 25608 17283 25664
rect 12268 25606 17283 25608
rect 12268 25604 12274 25606
rect 17217 25603 17283 25606
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 13905 25530 13971 25533
rect 10734 25528 13971 25530
rect 10734 25472 13910 25528
rect 13966 25472 13971 25528
rect 10734 25470 13971 25472
rect 0 25394 480 25424
rect 2773 25394 2839 25397
rect 0 25392 2839 25394
rect 0 25336 2778 25392
rect 2834 25336 2839 25392
rect 0 25334 2839 25336
rect 0 25304 480 25334
rect 2773 25331 2839 25334
rect 9213 25394 9279 25397
rect 10734 25394 10794 25470
rect 13905 25467 13971 25470
rect 14457 25530 14523 25533
rect 19374 25530 19380 25532
rect 14457 25528 19380 25530
rect 14457 25472 14462 25528
rect 14518 25472 19380 25528
rect 14457 25470 19380 25472
rect 14457 25467 14523 25470
rect 19374 25468 19380 25470
rect 19444 25468 19450 25532
rect 20253 25530 20319 25533
rect 25814 25530 25820 25532
rect 20253 25528 25820 25530
rect 20253 25472 20258 25528
rect 20314 25472 25820 25528
rect 20253 25470 25820 25472
rect 20253 25467 20319 25470
rect 25814 25468 25820 25470
rect 25884 25468 25890 25532
rect 19324 25394 19390 25397
rect 9213 25392 10794 25394
rect 9213 25336 9218 25392
rect 9274 25336 10794 25392
rect 9213 25334 10794 25336
rect 14460 25392 19390 25394
rect 14460 25336 19329 25392
rect 19385 25336 19390 25392
rect 14460 25334 19390 25336
rect 9213 25331 9279 25334
rect 9622 25196 9628 25260
rect 9692 25258 9698 25260
rect 14460 25258 14520 25334
rect 19324 25331 19390 25334
rect 20345 25394 20411 25397
rect 21214 25394 21220 25396
rect 20345 25392 21220 25394
rect 20345 25336 20350 25392
rect 20406 25336 21220 25392
rect 20345 25334 21220 25336
rect 20345 25331 20411 25334
rect 21214 25332 21220 25334
rect 21284 25332 21290 25396
rect 24761 25394 24827 25397
rect 27520 25394 28000 25424
rect 24761 25392 28000 25394
rect 24761 25336 24766 25392
rect 24822 25336 28000 25392
rect 24761 25334 28000 25336
rect 24761 25331 24827 25334
rect 27520 25304 28000 25334
rect 17217 25258 17283 25261
rect 23105 25258 23171 25261
rect 9692 25198 14520 25258
rect 14782 25198 15394 25258
rect 9692 25196 9698 25198
rect 7741 25122 7807 25125
rect 14641 25122 14707 25125
rect 7741 25120 14707 25122
rect 7741 25064 7746 25120
rect 7802 25064 14646 25120
rect 14702 25064 14707 25120
rect 7741 25062 14707 25064
rect 7741 25059 7807 25062
rect 14641 25059 14707 25062
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 9397 24986 9463 24989
rect 14782 24986 14842 25198
rect 15334 25122 15394 25198
rect 17217 25256 23171 25258
rect 17217 25200 17222 25256
rect 17278 25200 23110 25256
rect 23166 25200 23171 25256
rect 17217 25198 23171 25200
rect 17217 25195 17283 25198
rect 23105 25195 23171 25198
rect 23790 25122 23796 25124
rect 15334 25062 23796 25122
rect 23790 25060 23796 25062
rect 23860 25060 23866 25124
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 23422 24986 23428 24988
rect 9397 24984 14842 24986
rect 9397 24928 9402 24984
rect 9458 24928 14842 24984
rect 9397 24926 14842 24928
rect 15334 24926 23428 24986
rect 9397 24923 9463 24926
rect 0 24850 480 24880
rect 933 24850 999 24853
rect 0 24848 999 24850
rect 0 24792 938 24848
rect 994 24792 999 24848
rect 0 24790 999 24792
rect 0 24760 480 24790
rect 933 24787 999 24790
rect 3785 24850 3851 24853
rect 5165 24850 5231 24853
rect 3785 24848 5231 24850
rect 3785 24792 3790 24848
rect 3846 24792 5170 24848
rect 5226 24792 5231 24848
rect 3785 24790 5231 24792
rect 3785 24787 3851 24790
rect 5165 24787 5231 24790
rect 9489 24850 9555 24853
rect 11053 24850 11119 24853
rect 9489 24848 11119 24850
rect 9489 24792 9494 24848
rect 9550 24792 11058 24848
rect 11114 24792 11119 24848
rect 9489 24790 11119 24792
rect 9489 24787 9555 24790
rect 11053 24787 11119 24790
rect 11421 24850 11487 24853
rect 14273 24850 14339 24853
rect 14774 24850 14780 24852
rect 11421 24848 13738 24850
rect 11421 24792 11426 24848
rect 11482 24792 13738 24848
rect 11421 24790 13738 24792
rect 11421 24787 11487 24790
rect 1526 24652 1532 24716
rect 1596 24714 1602 24716
rect 2405 24714 2471 24717
rect 1596 24712 2471 24714
rect 1596 24656 2410 24712
rect 2466 24656 2471 24712
rect 1596 24654 2471 24656
rect 1596 24652 1602 24654
rect 2405 24651 2471 24654
rect 3233 24714 3299 24717
rect 4797 24714 4863 24717
rect 3233 24712 4863 24714
rect 3233 24656 3238 24712
rect 3294 24656 4802 24712
rect 4858 24656 4863 24712
rect 3233 24654 4863 24656
rect 3233 24651 3299 24654
rect 4797 24651 4863 24654
rect 10133 24714 10199 24717
rect 12985 24714 13051 24717
rect 10133 24712 13051 24714
rect 10133 24656 10138 24712
rect 10194 24656 12990 24712
rect 13046 24656 13051 24712
rect 10133 24654 13051 24656
rect 10133 24651 10199 24654
rect 12985 24651 13051 24654
rect 2129 24578 2195 24581
rect 8845 24578 8911 24581
rect 2129 24576 8911 24578
rect 2129 24520 2134 24576
rect 2190 24520 8850 24576
rect 8906 24520 8911 24576
rect 2129 24518 8911 24520
rect 2129 24515 2195 24518
rect 8845 24515 8911 24518
rect 11094 24516 11100 24580
rect 11164 24578 11170 24580
rect 11605 24578 11671 24581
rect 11164 24576 11671 24578
rect 11164 24520 11610 24576
rect 11666 24520 11671 24576
rect 11164 24518 11671 24520
rect 13678 24578 13738 24790
rect 14273 24848 14780 24850
rect 14273 24792 14278 24848
rect 14334 24792 14780 24848
rect 14273 24790 14780 24792
rect 14273 24787 14339 24790
rect 14774 24788 14780 24790
rect 14844 24788 14850 24852
rect 15101 24850 15167 24853
rect 15334 24850 15394 24926
rect 23422 24924 23428 24926
rect 23492 24924 23498 24988
rect 15101 24848 15394 24850
rect 15101 24792 15106 24848
rect 15162 24792 15394 24848
rect 15101 24790 15394 24792
rect 15101 24787 15167 24790
rect 16062 24788 16068 24852
rect 16132 24850 16138 24852
rect 20529 24850 20595 24853
rect 16132 24848 20595 24850
rect 16132 24792 20534 24848
rect 20590 24792 20595 24848
rect 16132 24790 20595 24792
rect 16132 24788 16138 24790
rect 20529 24787 20595 24790
rect 21817 24850 21883 24853
rect 23565 24850 23631 24853
rect 21817 24848 23631 24850
rect 21817 24792 21822 24848
rect 21878 24792 23570 24848
rect 23626 24792 23631 24848
rect 21817 24790 23631 24792
rect 21817 24787 21883 24790
rect 23565 24787 23631 24790
rect 25221 24850 25287 24853
rect 27520 24850 28000 24880
rect 25221 24848 28000 24850
rect 25221 24792 25226 24848
rect 25282 24792 28000 24848
rect 25221 24790 28000 24792
rect 25221 24787 25287 24790
rect 27520 24760 28000 24790
rect 14917 24714 14983 24717
rect 15285 24714 15351 24717
rect 21081 24714 21147 24717
rect 14917 24712 21147 24714
rect 14917 24656 14922 24712
rect 14978 24656 15290 24712
rect 15346 24656 21086 24712
rect 21142 24656 21147 24712
rect 14917 24654 21147 24656
rect 14917 24651 14983 24654
rect 15285 24651 15351 24654
rect 21081 24651 21147 24654
rect 24025 24714 24091 24717
rect 25865 24714 25931 24717
rect 24025 24712 25931 24714
rect 24025 24656 24030 24712
rect 24086 24656 25870 24712
rect 25926 24656 25931 24712
rect 24025 24654 25931 24656
rect 24025 24651 24091 24654
rect 25865 24651 25931 24654
rect 17125 24578 17191 24581
rect 13678 24576 17191 24578
rect 13678 24520 17130 24576
rect 17186 24520 17191 24576
rect 13678 24518 17191 24520
rect 11164 24516 11170 24518
rect 11605 24515 11671 24518
rect 17125 24515 17191 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 657 24442 723 24445
rect 9121 24442 9187 24445
rect 9489 24442 9555 24445
rect 657 24440 9555 24442
rect 657 24384 662 24440
rect 718 24384 9126 24440
rect 9182 24384 9494 24440
rect 9550 24384 9555 24440
rect 657 24382 9555 24384
rect 657 24379 723 24382
rect 9121 24379 9187 24382
rect 9489 24379 9555 24382
rect 12525 24442 12591 24445
rect 15377 24442 15443 24445
rect 17166 24442 17172 24444
rect 12525 24440 12634 24442
rect 12525 24384 12530 24440
rect 12586 24384 12634 24440
rect 12525 24379 12634 24384
rect 15377 24440 17172 24442
rect 15377 24384 15382 24440
rect 15438 24384 17172 24440
rect 15377 24382 17172 24384
rect 15377 24379 15443 24382
rect 17166 24380 17172 24382
rect 17236 24380 17242 24444
rect 24669 24442 24735 24445
rect 26509 24442 26575 24445
rect 24669 24440 26575 24442
rect 24669 24384 24674 24440
rect 24730 24384 26514 24440
rect 26570 24384 26575 24440
rect 24669 24382 26575 24384
rect 24669 24379 24735 24382
rect 26509 24379 26575 24382
rect 2221 24306 2287 24309
rect 6177 24306 6243 24309
rect 2221 24304 6243 24306
rect 2221 24248 2226 24304
rect 2282 24248 6182 24304
rect 6238 24248 6243 24304
rect 2221 24246 6243 24248
rect 2221 24243 2287 24246
rect 6177 24243 6243 24246
rect 6637 24306 6703 24309
rect 11421 24306 11487 24309
rect 6637 24304 11487 24306
rect 6637 24248 6642 24304
rect 6698 24248 11426 24304
rect 11482 24248 11487 24304
rect 6637 24246 11487 24248
rect 6637 24243 6703 24246
rect 11421 24243 11487 24246
rect 11605 24306 11671 24309
rect 12574 24306 12634 24379
rect 13353 24306 13419 24309
rect 11605 24304 13419 24306
rect 11605 24248 11610 24304
rect 11666 24248 13358 24304
rect 13414 24248 13419 24304
rect 11605 24246 13419 24248
rect 11605 24243 11671 24246
rect 13353 24243 13419 24246
rect 13905 24306 13971 24309
rect 19149 24306 19215 24309
rect 24393 24306 24459 24309
rect 13905 24304 15394 24306
rect 13905 24248 13910 24304
rect 13966 24248 15394 24304
rect 13905 24246 15394 24248
rect 13905 24243 13971 24246
rect 0 24170 480 24200
rect 1209 24170 1275 24173
rect 0 24168 1275 24170
rect 0 24112 1214 24168
rect 1270 24112 1275 24168
rect 0 24110 1275 24112
rect 0 24080 480 24110
rect 1209 24107 1275 24110
rect 9029 24170 9095 24173
rect 10685 24170 10751 24173
rect 14733 24170 14799 24173
rect 9029 24168 10751 24170
rect 9029 24112 9034 24168
rect 9090 24112 10690 24168
rect 10746 24112 10751 24168
rect 9029 24110 10751 24112
rect 9029 24107 9095 24110
rect 10685 24107 10751 24110
rect 11102 24168 14799 24170
rect 11102 24112 14738 24168
rect 14794 24112 14799 24168
rect 11102 24110 14799 24112
rect 8661 24034 8727 24037
rect 10961 24034 11027 24037
rect 8661 24032 11027 24034
rect 8661 23976 8666 24032
rect 8722 23976 10966 24032
rect 11022 23976 11027 24032
rect 8661 23974 11027 23976
rect 8661 23971 8727 23974
rect 10961 23971 11027 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 2814 23836 2820 23900
rect 2884 23898 2890 23900
rect 4245 23898 4311 23901
rect 2884 23896 4311 23898
rect 2884 23840 4250 23896
rect 4306 23840 4311 23896
rect 2884 23838 4311 23840
rect 2884 23836 2890 23838
rect 4245 23835 4311 23838
rect 6361 23898 6427 23901
rect 10777 23898 10843 23901
rect 6361 23896 10843 23898
rect 6361 23840 6366 23896
rect 6422 23840 10782 23896
rect 10838 23840 10843 23896
rect 6361 23838 10843 23840
rect 6361 23835 6427 23838
rect 10777 23835 10843 23838
rect 1945 23764 2011 23765
rect 1894 23700 1900 23764
rect 1964 23762 2011 23764
rect 3877 23762 3943 23765
rect 6821 23762 6887 23765
rect 1964 23760 2056 23762
rect 2006 23704 2056 23760
rect 1964 23702 2056 23704
rect 3877 23760 6887 23762
rect 3877 23704 3882 23760
rect 3938 23704 6826 23760
rect 6882 23704 6887 23760
rect 3877 23702 6887 23704
rect 1964 23700 2011 23702
rect 1945 23699 2011 23700
rect 3877 23699 3943 23702
rect 6821 23699 6887 23702
rect 7281 23762 7347 23765
rect 11102 23762 11162 24110
rect 14733 24107 14799 24110
rect 12433 24034 12499 24037
rect 14365 24034 14431 24037
rect 12433 24032 14431 24034
rect 12433 23976 12438 24032
rect 12494 23976 14370 24032
rect 14426 23976 14431 24032
rect 12433 23974 14431 23976
rect 15334 24034 15394 24246
rect 19149 24304 24459 24306
rect 19149 24248 19154 24304
rect 19210 24248 24398 24304
rect 24454 24248 24459 24304
rect 19149 24246 24459 24248
rect 19149 24243 19215 24246
rect 24393 24243 24459 24246
rect 16941 24170 17007 24173
rect 23013 24170 23079 24173
rect 27520 24170 28000 24200
rect 16941 24168 28000 24170
rect 16941 24112 16946 24168
rect 17002 24112 23018 24168
rect 23074 24112 28000 24168
rect 16941 24110 28000 24112
rect 16941 24107 17007 24110
rect 23013 24107 23079 24110
rect 27520 24080 28000 24110
rect 21398 24034 21404 24036
rect 15334 23974 21404 24034
rect 12433 23971 12499 23974
rect 14365 23971 14431 23974
rect 21398 23972 21404 23974
rect 21468 23972 21474 24036
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 17033 23898 17099 23901
rect 20069 23898 20135 23901
rect 17033 23896 20135 23898
rect 17033 23840 17038 23896
rect 17094 23840 20074 23896
rect 20130 23840 20135 23896
rect 17033 23838 20135 23840
rect 17033 23835 17099 23838
rect 20069 23835 20135 23838
rect 24761 23898 24827 23901
rect 27613 23898 27679 23901
rect 24761 23896 27679 23898
rect 24761 23840 24766 23896
rect 24822 23840 27618 23896
rect 27674 23840 27679 23896
rect 24761 23838 27679 23840
rect 24761 23835 24827 23838
rect 27613 23835 27679 23838
rect 11329 23762 11395 23765
rect 7281 23760 11395 23762
rect 7281 23704 7286 23760
rect 7342 23704 11334 23760
rect 11390 23704 11395 23760
rect 7281 23702 11395 23704
rect 7281 23699 7347 23702
rect 11329 23699 11395 23702
rect 13353 23762 13419 23765
rect 17493 23762 17559 23765
rect 22553 23762 22619 23765
rect 23657 23762 23723 23765
rect 13353 23760 16314 23762
rect 13353 23704 13358 23760
rect 13414 23704 16314 23760
rect 13353 23702 16314 23704
rect 13353 23699 13419 23702
rect 0 23626 480 23656
rect 3969 23626 4035 23629
rect 0 23624 4035 23626
rect 0 23568 3974 23624
rect 4030 23568 4035 23624
rect 0 23566 4035 23568
rect 0 23536 480 23566
rect 3969 23563 4035 23566
rect 4245 23626 4311 23629
rect 11605 23626 11671 23629
rect 4245 23624 11671 23626
rect 4245 23568 4250 23624
rect 4306 23568 11610 23624
rect 11666 23568 11671 23624
rect 4245 23566 11671 23568
rect 4245 23563 4311 23566
rect 11605 23563 11671 23566
rect 11881 23626 11947 23629
rect 16113 23626 16179 23629
rect 11881 23624 16179 23626
rect 11881 23568 11886 23624
rect 11942 23568 16118 23624
rect 16174 23568 16179 23624
rect 11881 23566 16179 23568
rect 16254 23626 16314 23702
rect 17493 23760 23723 23762
rect 17493 23704 17498 23760
rect 17554 23704 22558 23760
rect 22614 23704 23662 23760
rect 23718 23704 23723 23760
rect 17493 23702 23723 23704
rect 17493 23699 17559 23702
rect 22553 23699 22619 23702
rect 23657 23699 23723 23702
rect 23841 23762 23907 23765
rect 25313 23762 25379 23765
rect 23841 23760 25379 23762
rect 23841 23704 23846 23760
rect 23902 23704 25318 23760
rect 25374 23704 25379 23760
rect 23841 23702 25379 23704
rect 23841 23699 23907 23702
rect 25313 23699 25379 23702
rect 19977 23626 20043 23629
rect 27520 23626 28000 23656
rect 16254 23624 20043 23626
rect 16254 23568 19982 23624
rect 20038 23568 20043 23624
rect 16254 23566 20043 23568
rect 11881 23563 11947 23566
rect 16113 23563 16179 23566
rect 19977 23563 20043 23566
rect 24350 23566 28000 23626
rect 4061 23490 4127 23493
rect 7005 23490 7071 23493
rect 4061 23488 7071 23490
rect 4061 23432 4066 23488
rect 4122 23432 7010 23488
rect 7066 23432 7071 23488
rect 4061 23430 7071 23432
rect 4061 23427 4127 23430
rect 7005 23427 7071 23430
rect 12433 23490 12499 23493
rect 18229 23490 18295 23493
rect 18689 23490 18755 23493
rect 12433 23488 18755 23490
rect 12433 23432 12438 23488
rect 12494 23432 18234 23488
rect 18290 23432 18694 23488
rect 18750 23432 18755 23488
rect 12433 23430 18755 23432
rect 12433 23427 12499 23430
rect 18229 23427 18295 23430
rect 18689 23427 18755 23430
rect 21766 23428 21772 23492
rect 21836 23490 21842 23492
rect 22645 23490 22711 23493
rect 21836 23488 22711 23490
rect 21836 23432 22650 23488
rect 22706 23432 22711 23488
rect 21836 23430 22711 23432
rect 21836 23428 21842 23430
rect 22645 23427 22711 23430
rect 23657 23490 23723 23493
rect 24350 23490 24410 23566
rect 27520 23536 28000 23566
rect 23657 23488 24410 23490
rect 23657 23432 23662 23488
rect 23718 23432 24410 23488
rect 23657 23430 24410 23432
rect 24761 23490 24827 23493
rect 27061 23490 27127 23493
rect 24761 23488 27127 23490
rect 24761 23432 24766 23488
rect 24822 23432 27066 23488
rect 27122 23432 27127 23488
rect 24761 23430 27127 23432
rect 23657 23427 23723 23430
rect 24761 23427 24827 23430
rect 27061 23427 27127 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 7465 23354 7531 23357
rect 14273 23354 14339 23357
rect 17769 23354 17835 23357
rect 7465 23352 10058 23354
rect 7465 23296 7470 23352
rect 7526 23296 10058 23352
rect 7465 23294 10058 23296
rect 7465 23291 7531 23294
rect 9857 23218 9923 23221
rect 3374 23216 9923 23218
rect 3374 23160 9862 23216
rect 9918 23160 9923 23216
rect 3374 23158 9923 23160
rect 9998 23218 10058 23294
rect 14273 23352 17835 23354
rect 14273 23296 14278 23352
rect 14334 23296 17774 23352
rect 17830 23296 17835 23352
rect 14273 23294 17835 23296
rect 14273 23291 14339 23294
rect 17769 23291 17835 23294
rect 20989 23354 21055 23357
rect 25221 23354 25287 23357
rect 20989 23352 25287 23354
rect 20989 23296 20994 23352
rect 21050 23296 25226 23352
rect 25282 23296 25287 23352
rect 20989 23294 25287 23296
rect 20989 23291 21055 23294
rect 25221 23291 25287 23294
rect 11053 23218 11119 23221
rect 9998 23216 11119 23218
rect 9998 23160 11058 23216
rect 11114 23160 11119 23216
rect 9998 23158 11119 23160
rect 0 23082 480 23112
rect 3374 23082 3434 23158
rect 9857 23155 9923 23158
rect 11053 23155 11119 23158
rect 11421 23218 11487 23221
rect 16573 23218 16639 23221
rect 11421 23216 16639 23218
rect 11421 23160 11426 23216
rect 11482 23160 16578 23216
rect 16634 23160 16639 23216
rect 11421 23158 16639 23160
rect 11421 23155 11487 23158
rect 16573 23155 16639 23158
rect 17677 23218 17743 23221
rect 22277 23218 22343 23221
rect 17677 23216 22343 23218
rect 17677 23160 17682 23216
rect 17738 23160 22282 23216
rect 22338 23160 22343 23216
rect 17677 23158 22343 23160
rect 17677 23155 17743 23158
rect 22277 23155 22343 23158
rect 0 23022 3434 23082
rect 3509 23082 3575 23085
rect 8017 23082 8083 23085
rect 10777 23082 10843 23085
rect 3509 23080 8083 23082
rect 3509 23024 3514 23080
rect 3570 23024 8022 23080
rect 8078 23024 8083 23080
rect 3509 23022 8083 23024
rect 0 22992 480 23022
rect 3509 23019 3575 23022
rect 8017 23019 8083 23022
rect 9262 23080 10843 23082
rect 9262 23024 10782 23080
rect 10838 23024 10843 23080
rect 9262 23022 10843 23024
rect 4337 22946 4403 22949
rect 4294 22944 4403 22946
rect 4294 22888 4342 22944
rect 4398 22888 4403 22944
rect 4294 22883 4403 22888
rect 6361 22946 6427 22949
rect 8477 22946 8543 22949
rect 9262 22946 9322 23022
rect 10777 23019 10843 23022
rect 11237 23082 11303 23085
rect 17217 23082 17283 23085
rect 11237 23080 17283 23082
rect 11237 23024 11242 23080
rect 11298 23024 17222 23080
rect 17278 23024 17283 23080
rect 11237 23022 17283 23024
rect 11237 23019 11303 23022
rect 17217 23019 17283 23022
rect 18413 23082 18479 23085
rect 20437 23082 20503 23085
rect 20989 23082 21055 23085
rect 18413 23080 21055 23082
rect 18413 23024 18418 23080
rect 18474 23024 20442 23080
rect 20498 23024 20994 23080
rect 21050 23024 21055 23080
rect 18413 23022 21055 23024
rect 18413 23019 18479 23022
rect 20437 23019 20503 23022
rect 20989 23019 21055 23022
rect 21173 23082 21239 23085
rect 22829 23082 22895 23085
rect 21173 23080 22895 23082
rect 21173 23024 21178 23080
rect 21234 23024 22834 23080
rect 22890 23024 22895 23080
rect 21173 23022 22895 23024
rect 21173 23019 21239 23022
rect 22829 23019 22895 23022
rect 25405 23082 25471 23085
rect 27520 23082 28000 23112
rect 25405 23080 28000 23082
rect 25405 23024 25410 23080
rect 25466 23024 28000 23080
rect 25405 23022 28000 23024
rect 25405 23019 25471 23022
rect 27520 22992 28000 23022
rect 6361 22944 9322 22946
rect 6361 22888 6366 22944
rect 6422 22888 8482 22944
rect 8538 22888 9322 22944
rect 6361 22886 9322 22888
rect 9489 22946 9555 22949
rect 11145 22946 11211 22949
rect 12801 22946 12867 22949
rect 9489 22944 12867 22946
rect 9489 22888 9494 22944
rect 9550 22888 11150 22944
rect 11206 22888 12806 22944
rect 12862 22888 12867 22944
rect 9489 22886 12867 22888
rect 6361 22883 6427 22886
rect 8477 22883 8543 22886
rect 9489 22883 9555 22886
rect 11145 22883 11211 22886
rect 12801 22883 12867 22886
rect 17493 22946 17559 22949
rect 23657 22946 23723 22949
rect 17493 22944 23723 22946
rect 17493 22888 17498 22944
rect 17554 22888 23662 22944
rect 23718 22888 23723 22944
rect 17493 22886 23723 22888
rect 17493 22883 17559 22886
rect 23657 22883 23723 22886
rect 4294 22677 4354 22883
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 6177 22810 6243 22813
rect 11237 22810 11303 22813
rect 6177 22808 11303 22810
rect 6177 22752 6182 22808
rect 6238 22752 11242 22808
rect 11298 22752 11303 22808
rect 6177 22750 11303 22752
rect 6177 22747 6243 22750
rect 11237 22747 11303 22750
rect 12065 22810 12131 22813
rect 14733 22810 14799 22813
rect 12065 22808 14799 22810
rect 12065 22752 12070 22808
rect 12126 22752 14738 22808
rect 14794 22752 14799 22808
rect 12065 22750 14799 22752
rect 12065 22747 12131 22750
rect 14733 22747 14799 22750
rect 18505 22810 18571 22813
rect 18505 22808 20914 22810
rect 18505 22752 18510 22808
rect 18566 22752 20914 22808
rect 18505 22750 20914 22752
rect 18505 22747 18571 22750
rect 4294 22672 4403 22677
rect 4294 22616 4342 22672
rect 4398 22616 4403 22672
rect 4294 22614 4403 22616
rect 4337 22611 4403 22614
rect 10685 22674 10751 22677
rect 20713 22674 20779 22677
rect 10685 22672 20779 22674
rect 10685 22616 10690 22672
rect 10746 22616 20718 22672
rect 20774 22616 20779 22672
rect 10685 22614 20779 22616
rect 20854 22674 20914 22750
rect 23473 22674 23539 22677
rect 20854 22672 23539 22674
rect 20854 22616 23478 22672
rect 23534 22616 23539 22672
rect 20854 22614 23539 22616
rect 10685 22611 10751 22614
rect 20713 22611 20779 22614
rect 23473 22611 23539 22614
rect 0 22538 480 22568
rect 4061 22538 4127 22541
rect 0 22536 4127 22538
rect 0 22480 4066 22536
rect 4122 22480 4127 22536
rect 0 22478 4127 22480
rect 0 22448 480 22478
rect 4061 22475 4127 22478
rect 15561 22538 15627 22541
rect 19425 22538 19491 22541
rect 15561 22536 19491 22538
rect 15561 22480 15566 22536
rect 15622 22480 19430 22536
rect 19486 22480 19491 22536
rect 15561 22478 19491 22480
rect 15561 22475 15627 22478
rect 19425 22475 19491 22478
rect 19793 22538 19859 22541
rect 21173 22538 21239 22541
rect 19793 22536 21239 22538
rect 19793 22480 19798 22536
rect 19854 22480 21178 22536
rect 21234 22480 21239 22536
rect 19793 22478 21239 22480
rect 19793 22475 19859 22478
rect 21173 22475 21239 22478
rect 25129 22538 25195 22541
rect 27520 22538 28000 22568
rect 25129 22536 28000 22538
rect 25129 22480 25134 22536
rect 25190 22480 28000 22536
rect 25129 22478 28000 22480
rect 25129 22475 25195 22478
rect 27520 22448 28000 22478
rect 3325 22402 3391 22405
rect 5625 22402 5691 22405
rect 3325 22400 5691 22402
rect 3325 22344 3330 22400
rect 3386 22344 5630 22400
rect 5686 22344 5691 22400
rect 3325 22342 5691 22344
rect 3325 22339 3391 22342
rect 5625 22339 5691 22342
rect 17217 22402 17283 22405
rect 19241 22402 19307 22405
rect 17217 22400 19307 22402
rect 17217 22344 17222 22400
rect 17278 22344 19246 22400
rect 19302 22344 19307 22400
rect 17217 22342 19307 22344
rect 17217 22339 17283 22342
rect 19241 22339 19307 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 1894 22204 1900 22268
rect 1964 22204 1970 22268
rect 3182 22204 3188 22268
rect 3252 22266 3258 22268
rect 9438 22266 9444 22268
rect 3252 22206 9444 22266
rect 3252 22204 3258 22206
rect 9438 22204 9444 22206
rect 9508 22204 9514 22268
rect 12985 22266 13051 22269
rect 18229 22266 18295 22269
rect 12985 22264 18295 22266
rect 12985 22208 12990 22264
rect 13046 22208 18234 22264
rect 18290 22208 18295 22264
rect 12985 22206 18295 22208
rect 1902 22133 1962 22204
rect 12985 22203 13051 22206
rect 18229 22203 18295 22206
rect 18597 22266 18663 22269
rect 18965 22266 19031 22269
rect 18597 22264 19031 22266
rect 18597 22208 18602 22264
rect 18658 22208 18970 22264
rect 19026 22208 19031 22264
rect 18597 22206 19031 22208
rect 18597 22203 18663 22206
rect 18965 22203 19031 22206
rect 23749 22266 23815 22269
rect 23974 22266 23980 22268
rect 23749 22264 23980 22266
rect 23749 22208 23754 22264
rect 23810 22208 23980 22264
rect 23749 22206 23980 22208
rect 23749 22203 23815 22206
rect 23974 22204 23980 22206
rect 24044 22204 24050 22268
rect 1853 22128 1962 22133
rect 1853 22072 1858 22128
rect 1914 22072 1962 22128
rect 1853 22070 1962 22072
rect 4889 22130 4955 22133
rect 11697 22130 11763 22133
rect 4889 22128 11763 22130
rect 4889 22072 4894 22128
rect 4950 22072 11702 22128
rect 11758 22072 11763 22128
rect 4889 22070 11763 22072
rect 1853 22067 1919 22070
rect 4889 22067 4955 22070
rect 11697 22067 11763 22070
rect 11881 22130 11947 22133
rect 17033 22130 17099 22133
rect 11881 22128 17099 22130
rect 11881 22072 11886 22128
rect 11942 22072 17038 22128
rect 17094 22072 17099 22128
rect 11881 22070 17099 22072
rect 11881 22067 11947 22070
rect 17033 22067 17099 22070
rect 17309 22130 17375 22133
rect 24945 22130 25011 22133
rect 17309 22128 25011 22130
rect 17309 22072 17314 22128
rect 17370 22072 24950 22128
rect 25006 22072 25011 22128
rect 17309 22070 25011 22072
rect 17309 22067 17375 22070
rect 24945 22067 25011 22070
rect 5993 21994 6059 21997
rect 3926 21992 6059 21994
rect 3926 21936 5998 21992
rect 6054 21936 6059 21992
rect 3926 21934 6059 21936
rect 0 21858 480 21888
rect 3693 21858 3759 21861
rect 0 21856 3759 21858
rect 0 21800 3698 21856
rect 3754 21800 3759 21856
rect 0 21798 3759 21800
rect 0 21768 480 21798
rect 3693 21795 3759 21798
rect 3417 21722 3483 21725
rect 3926 21722 3986 21934
rect 5993 21931 6059 21934
rect 13997 21994 14063 21997
rect 15929 21994 15995 21997
rect 13997 21992 15995 21994
rect 13997 21936 14002 21992
rect 14058 21936 15934 21992
rect 15990 21936 15995 21992
rect 13997 21934 15995 21936
rect 13997 21931 14063 21934
rect 15929 21931 15995 21934
rect 23841 21994 23907 21997
rect 23974 21994 23980 21996
rect 23841 21992 23980 21994
rect 23841 21936 23846 21992
rect 23902 21936 23980 21992
rect 23841 21934 23980 21936
rect 23841 21931 23907 21934
rect 23974 21932 23980 21934
rect 24044 21932 24050 21996
rect 5993 21858 6059 21861
rect 13629 21858 13695 21861
rect 5993 21856 13695 21858
rect 5993 21800 5998 21856
rect 6054 21800 13634 21856
rect 13690 21800 13695 21856
rect 5993 21798 13695 21800
rect 5993 21795 6059 21798
rect 13629 21795 13695 21798
rect 17677 21858 17743 21861
rect 19793 21858 19859 21861
rect 17677 21856 19859 21858
rect 17677 21800 17682 21856
rect 17738 21800 19798 21856
rect 19854 21800 19859 21856
rect 17677 21798 19859 21800
rect 17677 21795 17743 21798
rect 19793 21795 19859 21798
rect 21541 21858 21607 21861
rect 24025 21858 24091 21861
rect 21541 21856 24091 21858
rect 21541 21800 21546 21856
rect 21602 21800 24030 21856
rect 24086 21800 24091 21856
rect 21541 21798 24091 21800
rect 21541 21795 21607 21798
rect 24025 21795 24091 21798
rect 25681 21858 25747 21861
rect 27520 21858 28000 21888
rect 25681 21856 28000 21858
rect 25681 21800 25686 21856
rect 25742 21800 28000 21856
rect 25681 21798 28000 21800
rect 25681 21795 25747 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 27520 21768 28000 21798
rect 24277 21727 24597 21728
rect 14181 21722 14247 21725
rect 3417 21720 3986 21722
rect 3417 21664 3422 21720
rect 3478 21664 3986 21720
rect 3417 21662 3986 21664
rect 6088 21720 14247 21722
rect 6088 21664 14186 21720
rect 14242 21664 14247 21720
rect 6088 21662 14247 21664
rect 3417 21659 3483 21662
rect 3233 21586 3299 21589
rect 6088 21586 6148 21662
rect 14181 21659 14247 21662
rect 16021 21722 16087 21725
rect 19701 21722 19767 21725
rect 16021 21720 19767 21722
rect 16021 21664 16026 21720
rect 16082 21664 19706 21720
rect 19762 21664 19767 21720
rect 16021 21662 19767 21664
rect 16021 21659 16087 21662
rect 19701 21659 19767 21662
rect 19885 21722 19951 21725
rect 22185 21722 22251 21725
rect 23933 21724 23999 21725
rect 23933 21722 23980 21724
rect 19885 21720 22251 21722
rect 19885 21664 19890 21720
rect 19946 21664 22190 21720
rect 22246 21664 22251 21720
rect 19885 21662 22251 21664
rect 23888 21720 23980 21722
rect 23888 21664 23938 21720
rect 23888 21662 23980 21664
rect 19885 21659 19951 21662
rect 22185 21659 22251 21662
rect 23933 21660 23980 21662
rect 24044 21660 24050 21724
rect 23933 21659 23999 21660
rect 3233 21584 6148 21586
rect 3233 21528 3238 21584
rect 3294 21528 6148 21584
rect 3233 21526 6148 21528
rect 8753 21586 8819 21589
rect 12249 21586 12315 21589
rect 8753 21584 12315 21586
rect 8753 21528 8758 21584
rect 8814 21528 12254 21584
rect 12310 21528 12315 21584
rect 8753 21526 12315 21528
rect 3233 21523 3299 21526
rect 8753 21523 8819 21526
rect 12249 21523 12315 21526
rect 20621 21586 20687 21589
rect 23933 21586 23999 21589
rect 20621 21584 23999 21586
rect 20621 21528 20626 21584
rect 20682 21528 23938 21584
rect 23994 21528 23999 21584
rect 20621 21526 23999 21528
rect 20621 21523 20687 21526
rect 23933 21523 23999 21526
rect 3417 21450 3483 21453
rect 5993 21450 6059 21453
rect 3417 21448 6059 21450
rect 3417 21392 3422 21448
rect 3478 21392 5998 21448
rect 6054 21392 6059 21448
rect 3417 21390 6059 21392
rect 3417 21387 3483 21390
rect 5993 21387 6059 21390
rect 19428 21390 20178 21450
rect 0 21314 480 21344
rect 2865 21314 2931 21317
rect 0 21312 2931 21314
rect 0 21256 2870 21312
rect 2926 21256 2931 21312
rect 0 21254 2931 21256
rect 0 21224 480 21254
rect 2865 21251 2931 21254
rect 15101 21314 15167 21317
rect 17033 21314 17099 21317
rect 15101 21312 17099 21314
rect 15101 21256 15106 21312
rect 15162 21256 17038 21312
rect 17094 21256 17099 21312
rect 15101 21254 17099 21256
rect 15101 21251 15167 21254
rect 17033 21251 17099 21254
rect 17166 21252 17172 21316
rect 17236 21314 17242 21316
rect 18229 21314 18295 21317
rect 19428 21314 19488 21390
rect 17236 21312 19488 21314
rect 17236 21256 18234 21312
rect 18290 21256 19488 21312
rect 17236 21254 19488 21256
rect 20118 21314 20178 21390
rect 20294 21388 20300 21452
rect 20364 21450 20370 21452
rect 20713 21450 20779 21453
rect 25262 21450 25268 21452
rect 20364 21448 25268 21450
rect 20364 21392 20718 21448
rect 20774 21392 25268 21448
rect 20364 21390 25268 21392
rect 20364 21388 20370 21390
rect 20713 21387 20779 21390
rect 25262 21388 25268 21390
rect 25332 21388 25338 21452
rect 24209 21314 24275 21317
rect 24577 21314 24643 21317
rect 20118 21312 24643 21314
rect 20118 21256 24214 21312
rect 24270 21256 24582 21312
rect 24638 21256 24643 21312
rect 20118 21254 24643 21256
rect 17236 21252 17242 21254
rect 18229 21251 18295 21254
rect 24209 21251 24275 21254
rect 24577 21251 24643 21254
rect 25221 21314 25287 21317
rect 27520 21314 28000 21344
rect 25221 21312 28000 21314
rect 25221 21256 25226 21312
rect 25282 21256 28000 21312
rect 25221 21254 28000 21256
rect 25221 21251 25287 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 27520 21224 28000 21254
rect 19610 21183 19930 21184
rect 1894 21116 1900 21180
rect 1964 21178 1970 21180
rect 5390 21178 5396 21180
rect 1964 21118 5396 21178
rect 1964 21116 1970 21118
rect 5390 21116 5396 21118
rect 5460 21116 5466 21180
rect 6729 21178 6795 21181
rect 8385 21178 8451 21181
rect 9213 21178 9279 21181
rect 6729 21176 8034 21178
rect 6729 21120 6734 21176
rect 6790 21120 8034 21176
rect 6729 21118 8034 21120
rect 6729 21115 6795 21118
rect 3233 21042 3299 21045
rect 7833 21042 7899 21045
rect 3233 21040 7899 21042
rect 3233 20984 3238 21040
rect 3294 20984 7838 21040
rect 7894 20984 7899 21040
rect 3233 20982 7899 20984
rect 7974 21042 8034 21118
rect 8385 21176 9279 21178
rect 8385 21120 8390 21176
rect 8446 21120 9218 21176
rect 9274 21120 9279 21176
rect 8385 21118 9279 21120
rect 8385 21115 8451 21118
rect 9213 21115 9279 21118
rect 13629 21178 13695 21181
rect 13905 21178 13971 21181
rect 16021 21178 16087 21181
rect 13629 21176 16087 21178
rect 13629 21120 13634 21176
rect 13690 21120 13910 21176
rect 13966 21120 16026 21176
rect 16082 21120 16087 21176
rect 13629 21118 16087 21120
rect 13629 21115 13695 21118
rect 13905 21115 13971 21118
rect 16021 21115 16087 21118
rect 16389 21178 16455 21181
rect 18137 21178 18203 21181
rect 16389 21176 18203 21178
rect 16389 21120 16394 21176
rect 16450 21120 18142 21176
rect 18198 21120 18203 21176
rect 16389 21118 18203 21120
rect 16389 21115 16455 21118
rect 18137 21115 18203 21118
rect 20713 21178 20779 21181
rect 21541 21178 21607 21181
rect 20713 21176 21607 21178
rect 20713 21120 20718 21176
rect 20774 21120 21546 21176
rect 21602 21120 21607 21176
rect 20713 21118 21607 21120
rect 20713 21115 20779 21118
rect 21541 21115 21607 21118
rect 10685 21042 10751 21045
rect 7974 21040 10751 21042
rect 7974 20984 10690 21040
rect 10746 20984 10751 21040
rect 7974 20982 10751 20984
rect 3233 20979 3299 20982
rect 7833 20979 7899 20982
rect 10685 20979 10751 20982
rect 11053 21042 11119 21045
rect 12709 21042 12775 21045
rect 11053 21040 12775 21042
rect 11053 20984 11058 21040
rect 11114 20984 12714 21040
rect 12770 20984 12775 21040
rect 11053 20982 12775 20984
rect 11053 20979 11119 20982
rect 12709 20979 12775 20982
rect 12985 21042 13051 21045
rect 22093 21042 22159 21045
rect 12985 21040 22159 21042
rect 12985 20984 12990 21040
rect 13046 20984 22098 21040
rect 22154 20984 22159 21040
rect 12985 20982 22159 20984
rect 12985 20979 13051 20982
rect 22093 20979 22159 20982
rect 9305 20906 9371 20909
rect 9806 20906 9812 20908
rect 9305 20904 9812 20906
rect 9305 20848 9310 20904
rect 9366 20848 9812 20904
rect 9305 20846 9812 20848
rect 9305 20843 9371 20846
rect 9806 20844 9812 20846
rect 9876 20906 9882 20908
rect 10133 20906 10199 20909
rect 9876 20904 10199 20906
rect 9876 20848 10138 20904
rect 10194 20848 10199 20904
rect 9876 20846 10199 20848
rect 9876 20844 9882 20846
rect 10133 20843 10199 20846
rect 12801 20906 12867 20909
rect 14825 20906 14891 20909
rect 17677 20906 17743 20909
rect 12801 20904 17743 20906
rect 12801 20848 12806 20904
rect 12862 20848 14830 20904
rect 14886 20848 17682 20904
rect 17738 20848 17743 20904
rect 12801 20846 17743 20848
rect 12801 20843 12867 20846
rect 14825 20843 14891 20846
rect 17677 20843 17743 20846
rect 0 20770 480 20800
rect 2405 20770 2471 20773
rect 0 20768 2471 20770
rect 0 20712 2410 20768
rect 2466 20712 2471 20768
rect 0 20710 2471 20712
rect 0 20680 480 20710
rect 2405 20707 2471 20710
rect 8201 20770 8267 20773
rect 10041 20770 10107 20773
rect 24025 20772 24091 20773
rect 8201 20768 10107 20770
rect 8201 20712 8206 20768
rect 8262 20712 10046 20768
rect 10102 20712 10107 20768
rect 8201 20710 10107 20712
rect 8201 20707 8267 20710
rect 10041 20707 10107 20710
rect 20110 20708 20116 20772
rect 20180 20770 20186 20772
rect 20846 20770 20852 20772
rect 20180 20710 20852 20770
rect 20180 20708 20186 20710
rect 20846 20708 20852 20710
rect 20916 20708 20922 20772
rect 23974 20708 23980 20772
rect 24044 20770 24091 20772
rect 27520 20770 28000 20800
rect 24044 20768 24136 20770
rect 24086 20712 24136 20768
rect 24044 20710 24136 20712
rect 25638 20710 28000 20770
rect 24044 20708 24091 20710
rect 24025 20707 24091 20708
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 9305 20634 9371 20637
rect 10777 20634 10843 20637
rect 9305 20632 10843 20634
rect 9305 20576 9310 20632
rect 9366 20576 10782 20632
rect 10838 20576 10843 20632
rect 9305 20574 10843 20576
rect 9305 20571 9371 20574
rect 10777 20571 10843 20574
rect 11237 20634 11303 20637
rect 13905 20634 13971 20637
rect 11237 20632 13971 20634
rect 11237 20576 11242 20632
rect 11298 20576 13910 20632
rect 13966 20576 13971 20632
rect 11237 20574 13971 20576
rect 11237 20571 11303 20574
rect 13905 20571 13971 20574
rect 15377 20634 15443 20637
rect 16481 20634 16547 20637
rect 20713 20634 20779 20637
rect 15377 20632 20779 20634
rect 15377 20576 15382 20632
rect 15438 20576 16486 20632
rect 16542 20576 20718 20632
rect 20774 20576 20779 20632
rect 15377 20574 20779 20576
rect 15377 20571 15443 20574
rect 16481 20571 16547 20574
rect 20713 20571 20779 20574
rect 25497 20634 25563 20637
rect 25638 20634 25698 20710
rect 27520 20680 28000 20710
rect 25497 20632 25698 20634
rect 25497 20576 25502 20632
rect 25558 20576 25698 20632
rect 25497 20574 25698 20576
rect 25497 20571 25563 20574
rect 3509 20498 3575 20501
rect 16389 20498 16455 20501
rect 19977 20498 20043 20501
rect 3509 20496 7114 20498
rect 3509 20440 3514 20496
rect 3570 20440 7114 20496
rect 3509 20438 7114 20440
rect 3509 20435 3575 20438
rect 2405 20362 2471 20365
rect 5809 20362 5875 20365
rect 2405 20360 5875 20362
rect 2405 20304 2410 20360
rect 2466 20304 5814 20360
rect 5870 20304 5875 20360
rect 2405 20302 5875 20304
rect 2405 20299 2471 20302
rect 5809 20299 5875 20302
rect 2865 20226 2931 20229
rect 6085 20226 6151 20229
rect 6913 20226 6979 20229
rect 2865 20224 6979 20226
rect 2865 20168 2870 20224
rect 2926 20168 6090 20224
rect 6146 20168 6918 20224
rect 6974 20168 6979 20224
rect 2865 20166 6979 20168
rect 7054 20226 7114 20438
rect 16389 20496 20043 20498
rect 16389 20440 16394 20496
rect 16450 20440 19982 20496
rect 20038 20440 20043 20496
rect 16389 20438 20043 20440
rect 16389 20435 16455 20438
rect 19977 20435 20043 20438
rect 7189 20362 7255 20365
rect 12065 20362 12131 20365
rect 7189 20360 12131 20362
rect 7189 20304 7194 20360
rect 7250 20304 12070 20360
rect 12126 20304 12131 20360
rect 7189 20302 12131 20304
rect 7189 20299 7255 20302
rect 12065 20299 12131 20302
rect 14273 20362 14339 20365
rect 16389 20362 16455 20365
rect 25957 20362 26023 20365
rect 14273 20360 26023 20362
rect 14273 20304 14278 20360
rect 14334 20304 16394 20360
rect 16450 20304 25962 20360
rect 26018 20304 26023 20360
rect 14273 20302 26023 20304
rect 14273 20299 14339 20302
rect 16389 20299 16455 20302
rect 25957 20299 26023 20302
rect 9673 20226 9739 20229
rect 10041 20228 10107 20229
rect 7054 20224 9739 20226
rect 7054 20168 9678 20224
rect 9734 20168 9739 20224
rect 7054 20166 9739 20168
rect 2865 20163 2931 20166
rect 6085 20163 6151 20166
rect 6913 20163 6979 20166
rect 9673 20163 9739 20166
rect 9990 20164 9996 20228
rect 10060 20226 10107 20228
rect 14825 20226 14891 20229
rect 15377 20226 15443 20229
rect 10060 20224 10152 20226
rect 10102 20168 10152 20224
rect 10060 20166 10152 20168
rect 14825 20224 15443 20226
rect 14825 20168 14830 20224
rect 14886 20168 15382 20224
rect 15438 20168 15443 20224
rect 14825 20166 15443 20168
rect 10060 20164 10107 20166
rect 10041 20163 10107 20164
rect 14825 20163 14891 20166
rect 15377 20163 15443 20166
rect 21214 20164 21220 20228
rect 21284 20226 21290 20228
rect 21633 20226 21699 20229
rect 21284 20224 21699 20226
rect 21284 20168 21638 20224
rect 21694 20168 21699 20224
rect 21284 20166 21699 20168
rect 21284 20164 21290 20166
rect 21633 20163 21699 20166
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 565 20090 631 20093
rect 0 20088 631 20090
rect 0 20032 570 20088
rect 626 20032 631 20088
rect 0 20030 631 20032
rect 0 20000 480 20030
rect 565 20027 631 20030
rect 6729 20090 6795 20093
rect 8293 20090 8359 20093
rect 12893 20092 12959 20093
rect 6729 20088 8359 20090
rect 6729 20032 6734 20088
rect 6790 20032 8298 20088
rect 8354 20032 8359 20088
rect 6729 20030 8359 20032
rect 6729 20027 6795 20030
rect 8293 20027 8359 20030
rect 10726 20028 10732 20092
rect 10796 20090 10802 20092
rect 12893 20090 12940 20092
rect 10796 20088 12940 20090
rect 10796 20032 12898 20088
rect 10796 20030 12940 20032
rect 10796 20028 10802 20030
rect 12893 20028 12940 20030
rect 13004 20028 13010 20092
rect 13445 20090 13511 20093
rect 15837 20090 15903 20093
rect 13445 20088 15903 20090
rect 13445 20032 13450 20088
rect 13506 20032 15842 20088
rect 15898 20032 15903 20088
rect 13445 20030 15903 20032
rect 12893 20027 12959 20028
rect 13445 20027 13511 20030
rect 15837 20027 15903 20030
rect 17033 20090 17099 20093
rect 18781 20090 18847 20093
rect 19149 20090 19215 20093
rect 22737 20092 22803 20093
rect 22686 20090 22692 20092
rect 17033 20088 19215 20090
rect 17033 20032 17038 20088
rect 17094 20032 18786 20088
rect 18842 20032 19154 20088
rect 19210 20032 19215 20088
rect 17033 20030 19215 20032
rect 22646 20030 22692 20090
rect 22756 20088 22803 20092
rect 22798 20032 22803 20088
rect 17033 20027 17099 20030
rect 18781 20027 18847 20030
rect 19149 20027 19215 20030
rect 22686 20028 22692 20030
rect 22756 20028 22803 20032
rect 22737 20027 22803 20028
rect 25405 20090 25471 20093
rect 27520 20090 28000 20120
rect 25405 20088 28000 20090
rect 25405 20032 25410 20088
rect 25466 20032 28000 20088
rect 25405 20030 28000 20032
rect 25405 20027 25471 20030
rect 27520 20000 28000 20030
rect 9622 19892 9628 19956
rect 9692 19954 9698 19956
rect 19382 19954 19580 19988
rect 24894 19954 24900 19956
rect 9692 19928 24900 19954
rect 9692 19894 19442 19928
rect 19520 19894 24900 19928
rect 9692 19892 9698 19894
rect 24894 19892 24900 19894
rect 24964 19892 24970 19956
rect 7925 19818 7991 19821
rect 11697 19818 11763 19821
rect 19324 19818 19390 19821
rect 7925 19816 11763 19818
rect 7925 19760 7930 19816
rect 7986 19760 11702 19816
rect 11758 19760 11763 19816
rect 7925 19758 11763 19760
rect 7925 19755 7991 19758
rect 11697 19755 11763 19758
rect 14460 19816 19390 19818
rect 14460 19760 19329 19816
rect 19385 19760 19390 19816
rect 14460 19758 19390 19760
rect 6177 19682 6243 19685
rect 14460 19682 14520 19758
rect 19324 19755 19390 19758
rect 22318 19756 22324 19820
rect 22388 19818 22394 19820
rect 25129 19818 25195 19821
rect 22388 19816 25195 19818
rect 22388 19760 25134 19816
rect 25190 19760 25195 19816
rect 22388 19758 25195 19760
rect 22388 19756 22394 19758
rect 25129 19755 25195 19758
rect 6177 19680 14520 19682
rect 6177 19624 6182 19680
rect 6238 19624 14520 19680
rect 6177 19622 14520 19624
rect 15837 19682 15903 19685
rect 23381 19682 23447 19685
rect 15837 19680 23447 19682
rect 15837 19624 15842 19680
rect 15898 19624 23386 19680
rect 23442 19624 23447 19680
rect 15837 19622 23447 19624
rect 6177 19619 6243 19622
rect 15837 19619 15903 19622
rect 23381 19619 23447 19622
rect 5610 19616 5930 19617
rect 0 19546 480 19576
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 16205 19546 16271 19549
rect 0 19486 5458 19546
rect 0 19456 480 19486
rect 5398 19410 5458 19486
rect 15702 19544 16271 19546
rect 15702 19488 16210 19544
rect 16266 19488 16271 19544
rect 15702 19486 16271 19488
rect 9489 19410 9555 19413
rect 15702 19410 15762 19486
rect 16205 19483 16271 19486
rect 16573 19546 16639 19549
rect 20253 19546 20319 19549
rect 16573 19544 20319 19546
rect 16573 19488 16578 19544
rect 16634 19488 20258 19544
rect 20314 19488 20319 19544
rect 16573 19486 20319 19488
rect 16573 19483 16639 19486
rect 20253 19483 20319 19486
rect 20529 19546 20595 19549
rect 21766 19546 21772 19548
rect 20529 19544 21772 19546
rect 20529 19488 20534 19544
rect 20590 19488 21772 19544
rect 20529 19486 21772 19488
rect 20529 19483 20595 19486
rect 21766 19484 21772 19486
rect 21836 19484 21842 19548
rect 25773 19546 25839 19549
rect 27520 19546 28000 19576
rect 25773 19544 28000 19546
rect 25773 19488 25778 19544
rect 25834 19488 28000 19544
rect 25773 19486 28000 19488
rect 25773 19483 25839 19486
rect 27520 19456 28000 19486
rect 5398 19408 9555 19410
rect 5398 19352 9494 19408
rect 9550 19352 9555 19408
rect 5398 19350 9555 19352
rect 9489 19347 9555 19350
rect 9630 19350 15762 19410
rect 15837 19410 15903 19413
rect 21541 19410 21607 19413
rect 15837 19408 21607 19410
rect 15837 19352 15842 19408
rect 15898 19352 21546 19408
rect 21602 19352 21607 19408
rect 15837 19350 21607 19352
rect 4470 19212 4476 19276
rect 4540 19274 4546 19276
rect 9630 19274 9690 19350
rect 15837 19347 15903 19350
rect 21541 19347 21607 19350
rect 22737 19410 22803 19413
rect 24485 19410 24551 19413
rect 22737 19408 24551 19410
rect 22737 19352 22742 19408
rect 22798 19352 24490 19408
rect 24546 19352 24551 19408
rect 22737 19350 24551 19352
rect 22737 19347 22803 19350
rect 24485 19347 24551 19350
rect 4540 19214 9690 19274
rect 16941 19274 17007 19277
rect 21725 19274 21791 19277
rect 16941 19272 21791 19274
rect 16941 19216 16946 19272
rect 17002 19216 21730 19272
rect 21786 19216 21791 19272
rect 16941 19214 21791 19216
rect 4540 19212 4546 19214
rect 16941 19211 17007 19214
rect 21725 19211 21791 19214
rect 14733 19138 14799 19141
rect 17769 19138 17835 19141
rect 14733 19136 17835 19138
rect 14733 19080 14738 19136
rect 14794 19080 17774 19136
rect 17830 19080 17835 19136
rect 14733 19078 17835 19080
rect 14733 19075 14799 19078
rect 17769 19075 17835 19078
rect 20069 19138 20135 19141
rect 22369 19138 22435 19141
rect 20069 19136 22435 19138
rect 20069 19080 20074 19136
rect 20130 19080 22374 19136
rect 22430 19080 22435 19136
rect 20069 19078 22435 19080
rect 20069 19075 20135 19078
rect 22369 19075 22435 19078
rect 10277 19072 10597 19073
rect 0 19002 480 19032
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 1393 19002 1459 19005
rect 0 19000 1459 19002
rect 0 18944 1398 19000
rect 1454 18944 1459 19000
rect 0 18942 1459 18944
rect 0 18912 480 18942
rect 1393 18939 1459 18942
rect 2773 19004 2839 19005
rect 2773 19000 2820 19004
rect 2884 19002 2890 19004
rect 2773 18944 2778 19000
rect 2773 18940 2820 18944
rect 2884 18942 2930 19002
rect 2884 18940 2890 18942
rect 14774 18940 14780 19004
rect 14844 19002 14850 19004
rect 25681 19002 25747 19005
rect 27520 19002 28000 19032
rect 14844 18942 19488 19002
rect 14844 18940 14850 18942
rect 2773 18939 2839 18940
rect 4153 18866 4219 18869
rect 5390 18866 5396 18868
rect 4153 18864 5396 18866
rect 4153 18808 4158 18864
rect 4214 18808 5396 18864
rect 4153 18806 5396 18808
rect 4153 18803 4219 18806
rect 5390 18804 5396 18806
rect 5460 18804 5466 18868
rect 7373 18866 7439 18869
rect 9673 18866 9739 18869
rect 7373 18864 9739 18866
rect 7373 18808 7378 18864
rect 7434 18808 9678 18864
rect 9734 18808 9739 18864
rect 7373 18806 9739 18808
rect 7373 18803 7439 18806
rect 9673 18803 9739 18806
rect 10685 18866 10751 18869
rect 11462 18866 11468 18868
rect 10685 18864 11468 18866
rect 10685 18808 10690 18864
rect 10746 18808 11468 18864
rect 10685 18806 11468 18808
rect 10685 18803 10751 18806
rect 11462 18804 11468 18806
rect 11532 18804 11538 18868
rect 18505 18866 18571 18869
rect 15748 18864 18571 18866
rect 15748 18808 18510 18864
rect 18566 18808 18571 18864
rect 15748 18806 18571 18808
rect 19428 18866 19488 18942
rect 25681 19000 28000 19002
rect 25681 18944 25686 19000
rect 25742 18944 28000 19000
rect 25681 18942 28000 18944
rect 25681 18939 25747 18942
rect 27520 18912 28000 18942
rect 20897 18866 20963 18869
rect 19428 18864 20963 18866
rect 19428 18808 20902 18864
rect 20958 18808 20963 18864
rect 19428 18806 20963 18808
rect 5993 18730 6059 18733
rect 7782 18730 7788 18732
rect 5993 18728 7788 18730
rect 5993 18672 5998 18728
rect 6054 18672 7788 18728
rect 5993 18670 7788 18672
rect 5993 18667 6059 18670
rect 7782 18668 7788 18670
rect 7852 18668 7858 18732
rect 15748 18730 15808 18806
rect 18505 18803 18571 18806
rect 20897 18803 20963 18806
rect 21081 18866 21147 18869
rect 23565 18866 23631 18869
rect 21081 18864 23631 18866
rect 21081 18808 21086 18864
rect 21142 18808 23570 18864
rect 23626 18808 23631 18864
rect 21081 18806 23631 18808
rect 21081 18803 21147 18806
rect 23565 18803 23631 18806
rect 7928 18670 15808 18730
rect 7373 18594 7439 18597
rect 7928 18594 7988 18670
rect 15878 18668 15884 18732
rect 15948 18730 15954 18732
rect 16205 18730 16271 18733
rect 15948 18728 16271 18730
rect 15948 18672 16210 18728
rect 16266 18672 16271 18728
rect 15948 18670 16271 18672
rect 15948 18668 15954 18670
rect 16205 18667 16271 18670
rect 17125 18730 17191 18733
rect 22461 18730 22527 18733
rect 17125 18728 22527 18730
rect 17125 18672 17130 18728
rect 17186 18672 22466 18728
rect 22522 18672 22527 18728
rect 17125 18670 22527 18672
rect 17125 18667 17191 18670
rect 22461 18667 22527 18670
rect 22870 18668 22876 18732
rect 22940 18730 22946 18732
rect 23013 18730 23079 18733
rect 22940 18728 23079 18730
rect 22940 18672 23018 18728
rect 23074 18672 23079 18728
rect 22940 18670 23079 18672
rect 22940 18668 22946 18670
rect 23013 18667 23079 18670
rect 23565 18730 23631 18733
rect 23974 18730 23980 18732
rect 23565 18728 23980 18730
rect 23565 18672 23570 18728
rect 23626 18672 23980 18728
rect 23565 18670 23980 18672
rect 23565 18667 23631 18670
rect 23974 18668 23980 18670
rect 24044 18668 24050 18732
rect 24485 18730 24551 18733
rect 24485 18728 25146 18730
rect 24485 18672 24490 18728
rect 24546 18672 25146 18728
rect 24485 18670 25146 18672
rect 24485 18667 24551 18670
rect 7373 18592 7988 18594
rect 7373 18536 7378 18592
rect 7434 18536 7988 18592
rect 7373 18534 7988 18536
rect 15653 18594 15719 18597
rect 20069 18594 20135 18597
rect 15653 18592 20135 18594
rect 15653 18536 15658 18592
rect 15714 18536 20074 18592
rect 20130 18536 20135 18592
rect 15653 18534 20135 18536
rect 7373 18531 7439 18534
rect 15653 18531 15719 18534
rect 20069 18531 20135 18534
rect 20294 18532 20300 18596
rect 20364 18594 20370 18596
rect 20437 18594 20503 18597
rect 20364 18592 20503 18594
rect 20364 18536 20442 18592
rect 20498 18536 20503 18592
rect 20364 18534 20503 18536
rect 20364 18532 20370 18534
rect 20437 18531 20503 18534
rect 21449 18594 21515 18597
rect 23657 18594 23723 18597
rect 24025 18594 24091 18597
rect 21449 18592 24091 18594
rect 21449 18536 21454 18592
rect 21510 18536 23662 18592
rect 23718 18536 24030 18592
rect 24086 18536 24091 18592
rect 21449 18534 24091 18536
rect 21449 18531 21515 18534
rect 23657 18531 23723 18534
rect 24025 18531 24091 18534
rect 5610 18528 5930 18529
rect 0 18458 480 18488
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 7465 18458 7531 18461
rect 8937 18458 9003 18461
rect 0 18398 4906 18458
rect 0 18368 480 18398
rect 1577 18322 1643 18325
rect 4061 18322 4127 18325
rect 4337 18322 4403 18325
rect 1577 18320 4403 18322
rect 1577 18264 1582 18320
rect 1638 18264 4066 18320
rect 4122 18264 4342 18320
rect 4398 18264 4403 18320
rect 1577 18262 4403 18264
rect 4846 18322 4906 18398
rect 7465 18456 9003 18458
rect 7465 18400 7470 18456
rect 7526 18400 8942 18456
rect 8998 18400 9003 18456
rect 7465 18398 9003 18400
rect 7465 18395 7531 18398
rect 8937 18395 9003 18398
rect 19057 18458 19123 18461
rect 21633 18458 21699 18461
rect 19057 18456 21699 18458
rect 19057 18400 19062 18456
rect 19118 18400 21638 18456
rect 21694 18400 21699 18456
rect 19057 18398 21699 18400
rect 19057 18395 19123 18398
rect 21633 18395 21699 18398
rect 8661 18322 8727 18325
rect 4846 18320 8727 18322
rect 4846 18264 8666 18320
rect 8722 18264 8727 18320
rect 4846 18262 8727 18264
rect 1577 18259 1643 18262
rect 4061 18259 4127 18262
rect 4337 18259 4403 18262
rect 8661 18259 8727 18262
rect 18321 18322 18387 18325
rect 24945 18322 25011 18325
rect 18321 18320 25011 18322
rect 18321 18264 18326 18320
rect 18382 18264 24950 18320
rect 25006 18264 25011 18320
rect 18321 18262 25011 18264
rect 25086 18322 25146 18670
rect 25221 18458 25287 18461
rect 27520 18458 28000 18488
rect 25221 18456 28000 18458
rect 25221 18400 25226 18456
rect 25282 18400 28000 18456
rect 25221 18398 28000 18400
rect 25221 18395 25287 18398
rect 27520 18368 28000 18398
rect 25497 18322 25563 18325
rect 25086 18320 25563 18322
rect 25086 18264 25502 18320
rect 25558 18264 25563 18320
rect 25086 18262 25563 18264
rect 18321 18259 18387 18262
rect 24945 18259 25011 18262
rect 25497 18259 25563 18262
rect 14365 18186 14431 18189
rect 10136 18184 14431 18186
rect 10136 18128 14370 18184
rect 14426 18128 14431 18184
rect 10136 18126 14431 18128
rect 6913 18050 6979 18053
rect 4708 18048 6979 18050
rect 4708 17992 6918 18048
rect 6974 17992 6979 18048
rect 4708 17990 6979 17992
rect 0 17778 480 17808
rect 4708 17778 4768 17990
rect 6913 17987 6979 17990
rect 7046 17988 7052 18052
rect 7116 18050 7122 18052
rect 7465 18050 7531 18053
rect 7116 18048 7531 18050
rect 7116 17992 7470 18048
rect 7526 17992 7531 18048
rect 7116 17990 7531 17992
rect 7116 17988 7122 17990
rect 7465 17987 7531 17990
rect 7833 18050 7899 18053
rect 10136 18050 10196 18126
rect 14365 18123 14431 18126
rect 15101 18186 15167 18189
rect 18597 18186 18663 18189
rect 24025 18186 24091 18189
rect 24761 18186 24827 18189
rect 15101 18184 18663 18186
rect 15101 18128 15106 18184
rect 15162 18128 18602 18184
rect 18658 18128 18663 18184
rect 15101 18126 18663 18128
rect 15101 18123 15167 18126
rect 18597 18123 18663 18126
rect 18830 18184 24827 18186
rect 18830 18128 24030 18184
rect 24086 18128 24766 18184
rect 24822 18128 24827 18184
rect 18830 18126 24827 18128
rect 7833 18048 10196 18050
rect 7833 17992 7838 18048
rect 7894 17992 10196 18048
rect 7833 17990 10196 17992
rect 11053 18050 11119 18053
rect 12157 18050 12223 18053
rect 12433 18050 12499 18053
rect 11053 18048 12499 18050
rect 11053 17992 11058 18048
rect 11114 17992 12162 18048
rect 12218 17992 12438 18048
rect 12494 17992 12499 18048
rect 11053 17990 12499 17992
rect 7833 17987 7899 17990
rect 11053 17987 11119 17990
rect 12157 17987 12223 17990
rect 12433 17987 12499 17990
rect 16481 18050 16547 18053
rect 18830 18050 18890 18126
rect 24025 18123 24091 18126
rect 24761 18123 24827 18126
rect 16481 18048 18890 18050
rect 16481 17992 16486 18048
rect 16542 17992 18890 18048
rect 16481 17990 18890 17992
rect 22185 18050 22251 18053
rect 22318 18050 22324 18052
rect 22185 18048 22324 18050
rect 22185 17992 22190 18048
rect 22246 17992 22324 18048
rect 22185 17990 22324 17992
rect 16481 17987 16547 17990
rect 22185 17987 22251 17990
rect 22318 17988 22324 17990
rect 22388 17988 22394 18052
rect 23606 17988 23612 18052
rect 23676 18050 23682 18052
rect 24710 18050 24716 18052
rect 23676 17990 24716 18050
rect 23676 17988 23682 17990
rect 24710 17988 24716 17990
rect 24780 17988 24786 18052
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 5165 17916 5231 17917
rect 5165 17914 5212 17916
rect 5120 17912 5212 17914
rect 5120 17856 5170 17912
rect 5120 17854 5212 17856
rect 5165 17852 5212 17854
rect 5276 17852 5282 17916
rect 9673 17914 9739 17917
rect 5398 17912 9739 17914
rect 5398 17856 9678 17912
rect 9734 17856 9739 17912
rect 5398 17854 9739 17856
rect 5165 17851 5231 17852
rect 0 17718 4768 17778
rect 5073 17778 5139 17781
rect 5398 17778 5458 17854
rect 9673 17851 9739 17854
rect 10869 17914 10935 17917
rect 11237 17914 11303 17917
rect 16113 17914 16179 17917
rect 18229 17914 18295 17917
rect 10869 17912 18295 17914
rect 10869 17856 10874 17912
rect 10930 17856 11242 17912
rect 11298 17856 16118 17912
rect 16174 17856 18234 17912
rect 18290 17856 18295 17912
rect 10869 17854 18295 17856
rect 10869 17851 10935 17854
rect 11237 17851 11303 17854
rect 16113 17851 16179 17854
rect 18229 17851 18295 17854
rect 21541 17914 21607 17917
rect 25129 17914 25195 17917
rect 21541 17912 25195 17914
rect 21541 17856 21546 17912
rect 21602 17856 25134 17912
rect 25190 17856 25195 17912
rect 21541 17854 25195 17856
rect 21541 17851 21607 17854
rect 25129 17851 25195 17854
rect 5073 17776 5458 17778
rect 5073 17720 5078 17776
rect 5134 17720 5458 17776
rect 5073 17718 5458 17720
rect 5625 17778 5691 17781
rect 14181 17778 14247 17781
rect 5625 17776 14247 17778
rect 5625 17720 5630 17776
rect 5686 17720 14186 17776
rect 14242 17720 14247 17776
rect 5625 17718 14247 17720
rect 0 17688 480 17718
rect 5073 17715 5139 17718
rect 5625 17715 5691 17718
rect 14181 17715 14247 17718
rect 18873 17778 18939 17781
rect 21909 17778 21975 17781
rect 18873 17776 21975 17778
rect 18873 17720 18878 17776
rect 18934 17720 21914 17776
rect 21970 17720 21975 17776
rect 18873 17718 21975 17720
rect 18873 17715 18939 17718
rect 21909 17715 21975 17718
rect 24761 17778 24827 17781
rect 27520 17778 28000 17808
rect 24761 17776 28000 17778
rect 24761 17720 24766 17776
rect 24822 17720 28000 17776
rect 24761 17718 28000 17720
rect 24761 17715 24827 17718
rect 27520 17688 28000 17718
rect 3693 17642 3759 17645
rect 6453 17642 6519 17645
rect 8937 17642 9003 17645
rect 17953 17642 18019 17645
rect 3693 17640 8770 17642
rect 3693 17584 3698 17640
rect 3754 17584 6458 17640
rect 6514 17584 8770 17640
rect 3693 17582 8770 17584
rect 3693 17579 3759 17582
rect 6453 17579 6519 17582
rect 2497 17506 2563 17509
rect 4153 17506 4219 17509
rect 2497 17504 4219 17506
rect 2497 17448 2502 17504
rect 2558 17448 4158 17504
rect 4214 17448 4219 17504
rect 2497 17446 4219 17448
rect 8710 17506 8770 17582
rect 8937 17640 18019 17642
rect 8937 17584 8942 17640
rect 8998 17584 17958 17640
rect 18014 17584 18019 17640
rect 8937 17582 18019 17584
rect 8937 17579 9003 17582
rect 17953 17579 18019 17582
rect 18137 17642 18203 17645
rect 23657 17642 23723 17645
rect 18137 17640 23723 17642
rect 18137 17584 18142 17640
rect 18198 17584 23662 17640
rect 23718 17584 23723 17640
rect 18137 17582 23723 17584
rect 18137 17579 18203 17582
rect 23657 17579 23723 17582
rect 14549 17506 14615 17509
rect 8710 17504 14615 17506
rect 8710 17448 14554 17504
rect 14610 17448 14615 17504
rect 8710 17446 14615 17448
rect 2497 17443 2563 17446
rect 4153 17443 4219 17446
rect 14549 17443 14615 17446
rect 18689 17506 18755 17509
rect 20345 17506 20411 17509
rect 21173 17506 21239 17509
rect 18689 17504 21239 17506
rect 18689 17448 18694 17504
rect 18750 17448 20350 17504
rect 20406 17448 21178 17504
rect 21234 17448 21239 17504
rect 18689 17446 21239 17448
rect 18689 17443 18755 17446
rect 20345 17443 20411 17446
rect 21173 17443 21239 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 2129 17370 2195 17373
rect 2814 17370 2820 17372
rect 2129 17368 2820 17370
rect 2129 17312 2134 17368
rect 2190 17312 2820 17368
rect 2129 17310 2820 17312
rect 2129 17307 2195 17310
rect 2814 17308 2820 17310
rect 2884 17308 2890 17372
rect 8569 17370 8635 17373
rect 11237 17370 11303 17373
rect 13077 17372 13143 17373
rect 13077 17370 13124 17372
rect 8569 17368 11303 17370
rect 8569 17312 8574 17368
rect 8630 17312 11242 17368
rect 11298 17312 11303 17368
rect 8569 17310 11303 17312
rect 13032 17368 13124 17370
rect 13032 17312 13082 17368
rect 13032 17310 13124 17312
rect 8569 17307 8635 17310
rect 11237 17307 11303 17310
rect 13077 17308 13124 17310
rect 13188 17308 13194 17372
rect 15837 17370 15903 17373
rect 16665 17370 16731 17373
rect 23473 17370 23539 17373
rect 15837 17368 23539 17370
rect 15837 17312 15842 17368
rect 15898 17312 16670 17368
rect 16726 17312 23478 17368
rect 23534 17312 23539 17368
rect 15837 17310 23539 17312
rect 13077 17307 13143 17308
rect 15837 17307 15903 17310
rect 16665 17307 16731 17310
rect 23473 17307 23539 17310
rect 0 17234 480 17264
rect 2957 17234 3023 17237
rect 0 17232 3023 17234
rect 0 17176 2962 17232
rect 3018 17176 3023 17232
rect 0 17174 3023 17176
rect 0 17144 480 17174
rect 2957 17171 3023 17174
rect 7649 17234 7715 17237
rect 9397 17234 9463 17237
rect 7649 17232 9463 17234
rect 7649 17176 7654 17232
rect 7710 17176 9402 17232
rect 9458 17176 9463 17232
rect 7649 17174 9463 17176
rect 7649 17171 7715 17174
rect 9397 17171 9463 17174
rect 12433 17234 12499 17237
rect 16481 17234 16547 17237
rect 21357 17234 21423 17237
rect 12433 17232 14612 17234
rect 12433 17176 12438 17232
rect 12494 17176 14612 17232
rect 12433 17174 14612 17176
rect 12433 17171 12499 17174
rect 1945 17098 2011 17101
rect 8017 17098 8083 17101
rect 14365 17098 14431 17101
rect 1945 17096 8083 17098
rect 1945 17040 1950 17096
rect 2006 17040 8022 17096
rect 8078 17040 8083 17096
rect 1945 17038 8083 17040
rect 1945 17035 2011 17038
rect 8017 17035 8083 17038
rect 8158 17096 14431 17098
rect 8158 17040 14370 17096
rect 14426 17040 14431 17096
rect 8158 17038 14431 17040
rect 14552 17098 14612 17174
rect 16481 17232 21423 17234
rect 16481 17176 16486 17232
rect 16542 17176 21362 17232
rect 21418 17176 21423 17232
rect 16481 17174 21423 17176
rect 16481 17171 16547 17174
rect 21357 17171 21423 17174
rect 23054 17172 23060 17236
rect 23124 17234 23130 17236
rect 24853 17234 24919 17237
rect 23124 17232 24919 17234
rect 23124 17176 24858 17232
rect 24914 17176 24919 17232
rect 23124 17174 24919 17176
rect 23124 17172 23130 17174
rect 24853 17171 24919 17174
rect 25957 17234 26023 17237
rect 27520 17234 28000 17264
rect 25957 17232 28000 17234
rect 25957 17176 25962 17232
rect 26018 17176 28000 17232
rect 25957 17174 28000 17176
rect 25957 17171 26023 17174
rect 27520 17144 28000 17174
rect 19190 17098 19196 17100
rect 14552 17038 19196 17098
rect 2773 16962 2839 16965
rect 5206 16962 5212 16964
rect 2773 16960 5212 16962
rect 2773 16904 2778 16960
rect 2834 16904 5212 16960
rect 2773 16902 5212 16904
rect 2773 16899 2839 16902
rect 5206 16900 5212 16902
rect 5276 16900 5282 16964
rect 6913 16962 6979 16965
rect 7189 16962 7255 16965
rect 8158 16962 8218 17038
rect 14365 17035 14431 17038
rect 19190 17036 19196 17038
rect 19260 17036 19266 17100
rect 19977 17098 20043 17101
rect 22185 17098 22251 17101
rect 19977 17096 22251 17098
rect 19977 17040 19982 17096
rect 20038 17040 22190 17096
rect 22246 17040 22251 17096
rect 19977 17038 22251 17040
rect 19977 17035 20043 17038
rect 22185 17035 22251 17038
rect 6913 16960 8218 16962
rect 6913 16904 6918 16960
rect 6974 16904 7194 16960
rect 7250 16904 8218 16960
rect 6913 16902 8218 16904
rect 17769 16962 17835 16965
rect 19425 16962 19491 16965
rect 17769 16960 19491 16962
rect 17769 16904 17774 16960
rect 17830 16904 19430 16960
rect 19486 16904 19491 16960
rect 17769 16902 19491 16904
rect 6913 16899 6979 16902
rect 7189 16899 7255 16902
rect 17769 16899 17835 16902
rect 19425 16899 19491 16902
rect 22093 16962 22159 16965
rect 23013 16962 23079 16965
rect 22093 16960 23079 16962
rect 22093 16904 22098 16960
rect 22154 16904 23018 16960
rect 23074 16904 23079 16960
rect 22093 16902 23079 16904
rect 22093 16899 22159 16902
rect 23013 16899 23079 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 4245 16826 4311 16829
rect 1350 16824 4311 16826
rect 1350 16768 4250 16824
rect 4306 16768 4311 16824
rect 1350 16766 4311 16768
rect 0 16690 480 16720
rect 1350 16690 1410 16766
rect 4245 16763 4311 16766
rect 4838 16764 4844 16828
rect 4908 16826 4914 16828
rect 4981 16826 5047 16829
rect 4908 16824 5047 16826
rect 4908 16768 4986 16824
rect 5042 16768 5047 16824
rect 4908 16766 5047 16768
rect 4908 16764 4914 16766
rect 4981 16763 5047 16766
rect 5441 16826 5507 16829
rect 14917 16826 14983 16829
rect 19241 16826 19307 16829
rect 5441 16824 7298 16826
rect 5441 16768 5446 16824
rect 5502 16768 7298 16824
rect 5441 16766 7298 16768
rect 5441 16763 5507 16766
rect 0 16630 1410 16690
rect 2405 16690 2471 16693
rect 3049 16690 3115 16693
rect 2405 16688 3115 16690
rect 2405 16632 2410 16688
rect 2466 16632 3054 16688
rect 3110 16632 3115 16688
rect 2405 16630 3115 16632
rect 0 16600 480 16630
rect 2405 16627 2471 16630
rect 3049 16627 3115 16630
rect 4061 16690 4127 16693
rect 7005 16690 7071 16693
rect 4061 16688 7071 16690
rect 4061 16632 4066 16688
rect 4122 16632 7010 16688
rect 7066 16632 7071 16688
rect 4061 16630 7071 16632
rect 4061 16627 4127 16630
rect 7005 16627 7071 16630
rect 2037 16554 2103 16557
rect 3141 16554 3207 16557
rect 2037 16552 3207 16554
rect 2037 16496 2042 16552
rect 2098 16496 3146 16552
rect 3202 16496 3207 16552
rect 2037 16494 3207 16496
rect 7238 16554 7298 16766
rect 14917 16824 19307 16826
rect 14917 16768 14922 16824
rect 14978 16768 19246 16824
rect 19302 16768 19307 16824
rect 14917 16766 19307 16768
rect 14917 16763 14983 16766
rect 19241 16763 19307 16766
rect 21265 16826 21331 16829
rect 25037 16826 25103 16829
rect 21265 16824 25103 16826
rect 21265 16768 21270 16824
rect 21326 16768 25042 16824
rect 25098 16768 25103 16824
rect 21265 16766 25103 16768
rect 21265 16763 21331 16766
rect 25037 16763 25103 16766
rect 13905 16692 13971 16693
rect 13854 16690 13860 16692
rect 13814 16630 13860 16690
rect 13924 16688 13971 16692
rect 13966 16632 13971 16688
rect 13854 16628 13860 16630
rect 13924 16628 13971 16632
rect 13905 16627 13971 16628
rect 14825 16690 14891 16693
rect 15101 16690 15167 16693
rect 19609 16690 19675 16693
rect 14825 16688 15026 16690
rect 14825 16632 14830 16688
rect 14886 16632 15026 16688
rect 14825 16630 15026 16632
rect 14825 16627 14891 16630
rect 11237 16554 11303 16557
rect 7238 16552 11303 16554
rect 7238 16496 11242 16552
rect 11298 16496 11303 16552
rect 7238 16494 11303 16496
rect 2037 16491 2103 16494
rect 3141 16491 3207 16494
rect 11237 16491 11303 16494
rect 11881 16554 11947 16557
rect 13169 16554 13235 16557
rect 11881 16552 13235 16554
rect 11881 16496 11886 16552
rect 11942 16496 13174 16552
rect 13230 16496 13235 16552
rect 11881 16494 13235 16496
rect 14966 16554 15026 16630
rect 15101 16688 19675 16690
rect 15101 16632 15106 16688
rect 15162 16632 19614 16688
rect 19670 16632 19675 16688
rect 15101 16630 19675 16632
rect 15101 16627 15167 16630
rect 19609 16627 19675 16630
rect 22645 16690 22711 16693
rect 27520 16690 28000 16720
rect 22645 16688 28000 16690
rect 22645 16632 22650 16688
rect 22706 16632 28000 16688
rect 22645 16630 28000 16632
rect 22645 16627 22711 16630
rect 27520 16600 28000 16630
rect 21766 16554 21772 16556
rect 14966 16494 21772 16554
rect 11881 16491 11947 16494
rect 13169 16491 13235 16494
rect 21766 16492 21772 16494
rect 21836 16492 21842 16556
rect 2405 16418 2471 16421
rect 5349 16418 5415 16421
rect 2405 16416 5415 16418
rect 2405 16360 2410 16416
rect 2466 16360 5354 16416
rect 5410 16360 5415 16416
rect 2405 16358 5415 16360
rect 2405 16355 2471 16358
rect 5349 16355 5415 16358
rect 9949 16418 10015 16421
rect 13537 16418 13603 16421
rect 9949 16416 13603 16418
rect 9949 16360 9954 16416
rect 10010 16360 13542 16416
rect 13598 16360 13603 16416
rect 9949 16358 13603 16360
rect 9949 16355 10015 16358
rect 13537 16355 13603 16358
rect 18137 16418 18203 16421
rect 18965 16418 19031 16421
rect 20897 16418 20963 16421
rect 18137 16416 20963 16418
rect 18137 16360 18142 16416
rect 18198 16360 18970 16416
rect 19026 16360 20902 16416
rect 20958 16360 20963 16416
rect 18137 16358 20963 16360
rect 18137 16355 18203 16358
rect 18965 16355 19031 16358
rect 20897 16355 20963 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 8477 16282 8543 16285
rect 12341 16282 12407 16285
rect 14774 16282 14780 16284
rect 8477 16280 12407 16282
rect 8477 16224 8482 16280
rect 8538 16224 12346 16280
rect 12402 16224 12407 16280
rect 8477 16222 12407 16224
rect 8477 16219 8543 16222
rect 12341 16219 12407 16222
rect 12758 16222 14780 16282
rect 1526 16084 1532 16148
rect 1596 16146 1602 16148
rect 1761 16146 1827 16149
rect 1596 16144 1827 16146
rect 1596 16088 1766 16144
rect 1822 16088 1827 16144
rect 1596 16086 1827 16088
rect 1596 16084 1602 16086
rect 1761 16083 1827 16086
rect 3785 16146 3851 16149
rect 8017 16146 8083 16149
rect 3785 16144 8083 16146
rect 3785 16088 3790 16144
rect 3846 16088 8022 16144
rect 8078 16088 8083 16144
rect 3785 16086 8083 16088
rect 3785 16083 3851 16086
rect 8017 16083 8083 16086
rect 8385 16146 8451 16149
rect 11094 16146 11100 16148
rect 8385 16144 11100 16146
rect 8385 16088 8390 16144
rect 8446 16088 11100 16144
rect 8385 16086 11100 16088
rect 8385 16083 8451 16086
rect 11094 16084 11100 16086
rect 11164 16084 11170 16148
rect 12014 16084 12020 16148
rect 12084 16146 12090 16148
rect 12758 16146 12818 16222
rect 14774 16220 14780 16222
rect 14844 16220 14850 16284
rect 22645 16282 22711 16285
rect 15334 16280 22711 16282
rect 15334 16224 22650 16280
rect 22706 16224 22711 16280
rect 15334 16222 22711 16224
rect 12084 16086 12818 16146
rect 12893 16146 12959 16149
rect 14365 16146 14431 16149
rect 15334 16146 15394 16222
rect 22645 16219 22711 16222
rect 12893 16144 15394 16146
rect 12893 16088 12898 16144
rect 12954 16088 14370 16144
rect 14426 16088 15394 16144
rect 12893 16086 15394 16088
rect 17861 16146 17927 16149
rect 21449 16146 21515 16149
rect 22001 16148 22067 16149
rect 21950 16146 21956 16148
rect 17861 16144 21515 16146
rect 17861 16088 17866 16144
rect 17922 16088 21454 16144
rect 21510 16088 21515 16144
rect 17861 16086 21515 16088
rect 21910 16086 21956 16146
rect 22020 16144 22067 16148
rect 22062 16088 22067 16144
rect 12084 16084 12090 16086
rect 12893 16083 12959 16086
rect 14365 16083 14431 16086
rect 17861 16083 17927 16086
rect 21449 16083 21515 16086
rect 21950 16084 21956 16086
rect 22020 16084 22067 16088
rect 22001 16083 22067 16084
rect 0 16010 480 16040
rect 4061 16010 4127 16013
rect 0 16008 4127 16010
rect 0 15952 4066 16008
rect 4122 15952 4127 16008
rect 0 15950 4127 15952
rect 0 15920 480 15950
rect 4061 15947 4127 15950
rect 5165 16010 5231 16013
rect 14273 16010 14339 16013
rect 5165 16008 14339 16010
rect 5165 15952 5170 16008
rect 5226 15952 14278 16008
rect 14334 15952 14339 16008
rect 5165 15950 14339 15952
rect 5165 15947 5231 15950
rect 14273 15947 14339 15950
rect 14917 16010 14983 16013
rect 26233 16010 26299 16013
rect 27520 16010 28000 16040
rect 14917 16008 26299 16010
rect 14917 15952 14922 16008
rect 14978 15952 26238 16008
rect 26294 15952 26299 16008
rect 14917 15950 26299 15952
rect 14917 15947 14983 15950
rect 26233 15947 26299 15950
rect 26558 15950 28000 16010
rect 3141 15874 3207 15877
rect 9857 15874 9923 15877
rect 3141 15872 9923 15874
rect 3141 15816 3146 15872
rect 3202 15816 9862 15872
rect 9918 15816 9923 15872
rect 3141 15814 9923 15816
rect 3141 15811 3207 15814
rect 9857 15811 9923 15814
rect 13445 15874 13511 15877
rect 19425 15874 19491 15877
rect 13445 15872 19491 15874
rect 13445 15816 13450 15872
rect 13506 15816 19430 15872
rect 19486 15816 19491 15872
rect 13445 15814 19491 15816
rect 13445 15811 13511 15814
rect 19425 15811 19491 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 5441 15738 5507 15741
rect 7557 15738 7623 15741
rect 8569 15738 8635 15741
rect 5441 15736 8635 15738
rect 5441 15680 5446 15736
rect 5502 15680 7562 15736
rect 7618 15680 8574 15736
rect 8630 15680 8635 15736
rect 5441 15678 8635 15680
rect 5441 15675 5507 15678
rect 7557 15675 7623 15678
rect 8569 15675 8635 15678
rect 8753 15738 8819 15741
rect 12157 15738 12223 15741
rect 13813 15738 13879 15741
rect 22001 15738 22067 15741
rect 24025 15738 24091 15741
rect 8753 15736 9644 15738
rect 8753 15680 8758 15736
rect 8814 15680 9644 15736
rect 8753 15678 9644 15680
rect 8753 15675 8819 15678
rect 5390 15540 5396 15604
rect 5460 15602 5466 15604
rect 6269 15602 6335 15605
rect 5460 15600 6335 15602
rect 5460 15544 6274 15600
rect 6330 15544 6335 15600
rect 5460 15542 6335 15544
rect 9584 15602 9644 15678
rect 12157 15736 13879 15738
rect 12157 15680 12162 15736
rect 12218 15680 13818 15736
rect 13874 15680 13879 15736
rect 12157 15678 13879 15680
rect 12157 15675 12223 15678
rect 13813 15675 13879 15678
rect 14000 15678 16636 15738
rect 11789 15602 11855 15605
rect 9584 15600 11855 15602
rect 9584 15544 11794 15600
rect 11850 15544 11855 15600
rect 9584 15542 11855 15544
rect 5460 15540 5466 15542
rect 6269 15539 6335 15542
rect 11789 15539 11855 15542
rect 13445 15602 13511 15605
rect 14000 15602 14060 15678
rect 13445 15600 14060 15602
rect 13445 15544 13450 15600
rect 13506 15544 14060 15600
rect 13445 15542 14060 15544
rect 16576 15602 16636 15678
rect 22001 15736 24091 15738
rect 22001 15680 22006 15736
rect 22062 15680 24030 15736
rect 24086 15680 24091 15736
rect 22001 15678 24091 15680
rect 22001 15675 22067 15678
rect 24025 15675 24091 15678
rect 25405 15738 25471 15741
rect 26558 15738 26618 15950
rect 27520 15920 28000 15950
rect 25405 15736 26618 15738
rect 25405 15680 25410 15736
rect 25466 15680 26618 15736
rect 25405 15678 26618 15680
rect 25405 15675 25471 15678
rect 25497 15602 25563 15605
rect 16576 15600 25563 15602
rect 16576 15544 25502 15600
rect 25558 15544 25563 15600
rect 16576 15542 25563 15544
rect 13445 15539 13511 15542
rect 25497 15539 25563 15542
rect 0 15466 480 15496
rect 3969 15466 4035 15469
rect 7741 15466 7807 15469
rect 0 15464 4035 15466
rect 0 15408 3974 15464
rect 4030 15408 4035 15464
rect 0 15406 4035 15408
rect 0 15376 480 15406
rect 3969 15403 4035 15406
rect 5214 15464 7807 15466
rect 5214 15408 7746 15464
rect 7802 15408 7807 15464
rect 5214 15406 7807 15408
rect 1669 15330 1735 15333
rect 5214 15330 5274 15406
rect 7741 15403 7807 15406
rect 8017 15466 8083 15469
rect 11513 15466 11579 15469
rect 13537 15466 13603 15469
rect 8017 15464 11579 15466
rect 8017 15408 8022 15464
rect 8078 15408 11518 15464
rect 11574 15408 11579 15464
rect 8017 15406 11579 15408
rect 8017 15403 8083 15406
rect 11513 15403 11579 15406
rect 11654 15464 13603 15466
rect 11654 15408 13542 15464
rect 13598 15408 13603 15464
rect 11654 15406 13603 15408
rect 1669 15328 5274 15330
rect 1669 15272 1674 15328
rect 1730 15272 5274 15328
rect 1669 15270 5274 15272
rect 7005 15330 7071 15333
rect 8661 15330 8727 15333
rect 7005 15328 8727 15330
rect 7005 15272 7010 15328
rect 7066 15272 8666 15328
rect 8722 15272 8727 15328
rect 7005 15270 8727 15272
rect 1669 15267 1735 15270
rect 7005 15267 7071 15270
rect 8661 15267 8727 15270
rect 8845 15330 8911 15333
rect 11654 15330 11714 15406
rect 13537 15403 13603 15406
rect 13721 15466 13787 15469
rect 14641 15466 14707 15469
rect 14917 15466 14983 15469
rect 13721 15464 14983 15466
rect 13721 15408 13726 15464
rect 13782 15408 14646 15464
rect 14702 15408 14922 15464
rect 14978 15408 14983 15464
rect 13721 15406 14983 15408
rect 13721 15403 13787 15406
rect 14641 15403 14707 15406
rect 14917 15403 14983 15406
rect 15101 15466 15167 15469
rect 16021 15466 16087 15469
rect 18229 15466 18295 15469
rect 15101 15464 18295 15466
rect 15101 15408 15106 15464
rect 15162 15408 16026 15464
rect 16082 15408 18234 15464
rect 18290 15408 18295 15464
rect 15101 15406 18295 15408
rect 15101 15403 15167 15406
rect 16021 15403 16087 15406
rect 18229 15403 18295 15406
rect 22093 15468 22159 15469
rect 22093 15464 22140 15468
rect 22204 15466 22210 15468
rect 25313 15466 25379 15469
rect 27520 15466 28000 15496
rect 22093 15408 22098 15464
rect 22093 15404 22140 15408
rect 22204 15406 22250 15466
rect 25313 15464 28000 15466
rect 25313 15408 25318 15464
rect 25374 15408 28000 15464
rect 25313 15406 28000 15408
rect 22204 15404 22210 15406
rect 22093 15403 22159 15404
rect 25313 15403 25379 15406
rect 27520 15376 28000 15406
rect 8845 15328 11714 15330
rect 8845 15272 8850 15328
rect 8906 15272 11714 15328
rect 8845 15270 11714 15272
rect 11789 15330 11855 15333
rect 14181 15330 14247 15333
rect 11789 15328 14247 15330
rect 11789 15272 11794 15328
rect 11850 15272 14186 15328
rect 14242 15272 14247 15328
rect 11789 15270 14247 15272
rect 8845 15267 8911 15270
rect 11789 15267 11855 15270
rect 14181 15267 14247 15270
rect 15653 15330 15719 15333
rect 18505 15330 18571 15333
rect 15653 15328 18571 15330
rect 15653 15272 15658 15328
rect 15714 15272 18510 15328
rect 18566 15272 18571 15328
rect 15653 15270 18571 15272
rect 15653 15267 15719 15270
rect 18505 15267 18571 15270
rect 19057 15330 19123 15333
rect 19057 15328 21834 15330
rect 19057 15272 19062 15328
rect 19118 15272 21834 15328
rect 19057 15270 21834 15272
rect 19057 15267 19123 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 2405 15194 2471 15197
rect 3785 15194 3851 15197
rect 7741 15196 7807 15197
rect 7741 15194 7788 15196
rect 2405 15192 3851 15194
rect 2405 15136 2410 15192
rect 2466 15136 3790 15192
rect 3846 15136 3851 15192
rect 2405 15134 3851 15136
rect 7696 15192 7788 15194
rect 7696 15136 7746 15192
rect 7696 15134 7788 15136
rect 2405 15131 2471 15134
rect 3785 15131 3851 15134
rect 7741 15132 7788 15134
rect 7852 15132 7858 15196
rect 9397 15194 9463 15197
rect 11329 15194 11395 15197
rect 13629 15194 13695 15197
rect 14273 15194 14339 15197
rect 9397 15192 11162 15194
rect 9397 15136 9402 15192
rect 9458 15136 11162 15192
rect 9397 15134 11162 15136
rect 7741 15131 7807 15132
rect 9397 15131 9463 15134
rect 1577 15058 1643 15061
rect 6729 15058 6795 15061
rect 10869 15058 10935 15061
rect 1577 15056 10935 15058
rect 1577 15000 1582 15056
rect 1638 15000 6734 15056
rect 6790 15000 10874 15056
rect 10930 15000 10935 15056
rect 1577 14998 10935 15000
rect 11102 15058 11162 15134
rect 11329 15192 14339 15194
rect 11329 15136 11334 15192
rect 11390 15136 13634 15192
rect 13690 15136 14278 15192
rect 14334 15136 14339 15192
rect 11329 15134 14339 15136
rect 11329 15131 11395 15134
rect 13629 15131 13695 15134
rect 14273 15131 14339 15134
rect 19374 15132 19380 15196
rect 19444 15194 19450 15196
rect 19517 15194 19583 15197
rect 19444 15192 19583 15194
rect 19444 15136 19522 15192
rect 19578 15136 19583 15192
rect 19444 15134 19583 15136
rect 21774 15194 21834 15270
rect 21950 15268 21956 15332
rect 22020 15330 22026 15332
rect 22093 15330 22159 15333
rect 23933 15330 23999 15333
rect 22020 15328 22159 15330
rect 22020 15272 22098 15328
rect 22154 15272 22159 15328
rect 22020 15270 22159 15272
rect 22020 15268 22026 15270
rect 22093 15267 22159 15270
rect 22326 15328 23999 15330
rect 22326 15272 23938 15328
rect 23994 15272 23999 15328
rect 22326 15270 23999 15272
rect 22326 15194 22386 15270
rect 23933 15267 23999 15270
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 21774 15134 22386 15194
rect 19444 15132 19450 15134
rect 19517 15131 19583 15134
rect 13670 15058 13676 15060
rect 11102 14998 13676 15058
rect 1577 14995 1643 14998
rect 6729 14995 6795 14998
rect 10869 14995 10935 14998
rect 13670 14996 13676 14998
rect 13740 14996 13746 15060
rect 14917 15058 14983 15061
rect 26233 15058 26299 15061
rect 14917 15056 26299 15058
rect 14917 15000 14922 15056
rect 14978 15000 26238 15056
rect 26294 15000 26299 15056
rect 14917 14998 26299 15000
rect 14917 14995 14983 14998
rect 26233 14995 26299 14998
rect 0 14922 480 14952
rect 1577 14922 1643 14925
rect 0 14920 1643 14922
rect 0 14864 1582 14920
rect 1638 14864 1643 14920
rect 0 14862 1643 14864
rect 0 14832 480 14862
rect 1577 14859 1643 14862
rect 4245 14922 4311 14925
rect 12617 14922 12683 14925
rect 13353 14922 13419 14925
rect 4245 14920 13419 14922
rect 4245 14864 4250 14920
rect 4306 14864 12622 14920
rect 12678 14864 13358 14920
rect 13414 14864 13419 14920
rect 4245 14862 13419 14864
rect 4245 14859 4311 14862
rect 12617 14859 12683 14862
rect 13353 14859 13419 14862
rect 16849 14922 16915 14925
rect 20253 14922 20319 14925
rect 23473 14922 23539 14925
rect 16849 14920 20178 14922
rect 16849 14864 16854 14920
rect 16910 14864 20178 14920
rect 16849 14862 20178 14864
rect 16849 14859 16915 14862
rect 6361 14788 6427 14789
rect 6310 14786 6316 14788
rect 6270 14726 6316 14786
rect 6380 14784 6427 14788
rect 6422 14728 6427 14784
rect 6310 14724 6316 14726
rect 6380 14724 6427 14728
rect 20118 14786 20178 14862
rect 20253 14920 23539 14922
rect 20253 14864 20258 14920
rect 20314 14864 23478 14920
rect 23534 14864 23539 14920
rect 20253 14862 23539 14864
rect 20253 14859 20319 14862
rect 23473 14859 23539 14862
rect 24761 14922 24827 14925
rect 27520 14922 28000 14952
rect 24761 14920 28000 14922
rect 24761 14864 24766 14920
rect 24822 14864 28000 14920
rect 24761 14862 28000 14864
rect 24761 14859 24827 14862
rect 27520 14832 28000 14862
rect 21173 14786 21239 14789
rect 20118 14784 21239 14786
rect 20118 14728 21178 14784
rect 21234 14728 21239 14784
rect 20118 14726 21239 14728
rect 6361 14723 6427 14724
rect 21173 14723 21239 14726
rect 23054 14724 23060 14788
rect 23124 14786 23130 14788
rect 25630 14786 25636 14788
rect 23124 14726 25636 14786
rect 23124 14724 23130 14726
rect 25630 14724 25636 14726
rect 25700 14724 25706 14788
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 2405 14650 2471 14653
rect 6177 14650 6243 14653
rect 2405 14648 6243 14650
rect 2405 14592 2410 14648
rect 2466 14592 6182 14648
rect 6238 14592 6243 14648
rect 2405 14590 6243 14592
rect 2405 14587 2471 14590
rect 6177 14587 6243 14590
rect 6361 14650 6427 14653
rect 8569 14650 8635 14653
rect 6361 14648 8635 14650
rect 6361 14592 6366 14648
rect 6422 14592 8574 14648
rect 8630 14592 8635 14648
rect 6361 14590 8635 14592
rect 6361 14587 6427 14590
rect 8569 14587 8635 14590
rect 10961 14650 11027 14653
rect 12014 14650 12020 14652
rect 10961 14648 12020 14650
rect 10961 14592 10966 14648
rect 11022 14592 12020 14648
rect 10961 14590 12020 14592
rect 10961 14587 11027 14590
rect 12014 14588 12020 14590
rect 12084 14588 12090 14652
rect 13813 14650 13879 14653
rect 18689 14650 18755 14653
rect 13813 14648 18755 14650
rect 13813 14592 13818 14648
rect 13874 14592 18694 14648
rect 18750 14592 18755 14648
rect 13813 14590 18755 14592
rect 13813 14587 13879 14590
rect 18689 14587 18755 14590
rect 20294 14588 20300 14652
rect 20364 14650 20370 14652
rect 22185 14650 22251 14653
rect 20364 14648 22251 14650
rect 20364 14592 22190 14648
rect 22246 14592 22251 14648
rect 20364 14590 22251 14592
rect 20364 14588 20370 14590
rect 22185 14587 22251 14590
rect 23381 14650 23447 14653
rect 23606 14650 23612 14652
rect 23381 14648 23612 14650
rect 23381 14592 23386 14648
rect 23442 14592 23612 14648
rect 23381 14590 23612 14592
rect 23381 14587 23447 14590
rect 23606 14588 23612 14590
rect 23676 14588 23682 14652
rect 4797 14514 4863 14517
rect 10593 14514 10659 14517
rect 12893 14514 12959 14517
rect 18597 14514 18663 14517
rect 20897 14514 20963 14517
rect 4797 14512 7114 14514
rect 4797 14456 4802 14512
rect 4858 14456 7114 14512
rect 4797 14454 7114 14456
rect 4797 14451 4863 14454
rect 0 14378 480 14408
rect 6913 14378 6979 14381
rect 0 14376 6979 14378
rect 0 14320 6918 14376
rect 6974 14320 6979 14376
rect 0 14318 6979 14320
rect 0 14288 480 14318
rect 6913 14315 6979 14318
rect 7054 14242 7114 14454
rect 10593 14512 15762 14514
rect 10593 14456 10598 14512
rect 10654 14456 12898 14512
rect 12954 14456 15762 14512
rect 10593 14454 15762 14456
rect 10593 14451 10659 14454
rect 12893 14451 12959 14454
rect 8017 14378 8083 14381
rect 11237 14378 11303 14381
rect 12985 14378 13051 14381
rect 8017 14376 11303 14378
rect 8017 14320 8022 14376
rect 8078 14320 11242 14376
rect 11298 14320 11303 14376
rect 8017 14318 11303 14320
rect 8017 14315 8083 14318
rect 11237 14315 11303 14318
rect 11470 14376 13051 14378
rect 11470 14320 12990 14376
rect 13046 14320 13051 14376
rect 11470 14318 13051 14320
rect 11329 14242 11395 14245
rect 7054 14240 11395 14242
rect 7054 14184 11334 14240
rect 11390 14184 11395 14240
rect 7054 14182 11395 14184
rect 11329 14179 11395 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 8201 14106 8267 14109
rect 11470 14106 11530 14318
rect 12985 14315 13051 14318
rect 13169 14378 13235 14381
rect 15285 14378 15351 14381
rect 13169 14376 15351 14378
rect 13169 14320 13174 14376
rect 13230 14320 15290 14376
rect 15346 14320 15351 14376
rect 13169 14318 15351 14320
rect 15702 14378 15762 14454
rect 18597 14512 20963 14514
rect 18597 14456 18602 14512
rect 18658 14456 20902 14512
rect 20958 14456 20963 14512
rect 18597 14454 20963 14456
rect 18597 14451 18663 14454
rect 20897 14451 20963 14454
rect 22645 14514 22711 14517
rect 22645 14512 26434 14514
rect 22645 14456 22650 14512
rect 22706 14456 26434 14512
rect 22645 14454 26434 14456
rect 22645 14451 22711 14454
rect 26233 14378 26299 14381
rect 15702 14376 26299 14378
rect 15702 14320 26238 14376
rect 26294 14320 26299 14376
rect 15702 14318 26299 14320
rect 26374 14378 26434 14454
rect 27520 14378 28000 14408
rect 26374 14318 28000 14378
rect 13169 14315 13235 14318
rect 15285 14315 15351 14318
rect 26233 14315 26299 14318
rect 27520 14288 28000 14318
rect 11973 14242 12039 14245
rect 14365 14242 14431 14245
rect 11973 14240 14431 14242
rect 11973 14184 11978 14240
rect 12034 14184 14370 14240
rect 14426 14184 14431 14240
rect 11973 14182 14431 14184
rect 11973 14179 12039 14182
rect 14365 14179 14431 14182
rect 17401 14242 17467 14245
rect 20805 14242 20871 14245
rect 17401 14240 20871 14242
rect 17401 14184 17406 14240
rect 17462 14184 20810 14240
rect 20866 14184 20871 14240
rect 17401 14182 20871 14184
rect 17401 14179 17467 14182
rect 20805 14179 20871 14182
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 8201 14104 11530 14106
rect 8201 14048 8206 14104
rect 8262 14048 11530 14104
rect 8201 14046 11530 14048
rect 17953 14106 18019 14109
rect 20621 14106 20687 14109
rect 17953 14104 20687 14106
rect 17953 14048 17958 14104
rect 18014 14048 20626 14104
rect 20682 14048 20687 14104
rect 17953 14046 20687 14048
rect 8201 14043 8267 14046
rect 17953 14043 18019 14046
rect 20621 14043 20687 14046
rect 4981 13970 5047 13973
rect 9029 13970 9095 13973
rect 9305 13972 9371 13973
rect 9254 13970 9260 13972
rect 4981 13968 9095 13970
rect 4981 13912 4986 13968
rect 5042 13912 9034 13968
rect 9090 13912 9095 13968
rect 4981 13910 9095 13912
rect 9214 13910 9260 13970
rect 9324 13970 9371 13972
rect 14406 13970 14412 13972
rect 9324 13968 14412 13970
rect 9366 13912 14412 13968
rect 4981 13907 5047 13910
rect 9029 13907 9095 13910
rect 9254 13908 9260 13910
rect 9324 13910 14412 13912
rect 9324 13908 9371 13910
rect 14406 13908 14412 13910
rect 14476 13908 14482 13972
rect 25773 13970 25839 13973
rect 15150 13968 25839 13970
rect 15150 13912 25778 13968
rect 25834 13912 25839 13968
rect 15150 13910 25839 13912
rect 9305 13907 9371 13908
rect 5349 13834 5415 13837
rect 8385 13834 8451 13837
rect 5349 13832 8451 13834
rect 5349 13776 5354 13832
rect 5410 13776 8390 13832
rect 8446 13776 8451 13832
rect 5349 13774 8451 13776
rect 5349 13771 5415 13774
rect 8385 13771 8451 13774
rect 9121 13834 9187 13837
rect 9673 13834 9739 13837
rect 10961 13834 11027 13837
rect 9121 13832 11027 13834
rect 9121 13776 9126 13832
rect 9182 13776 9678 13832
rect 9734 13776 10966 13832
rect 11022 13776 11027 13832
rect 9121 13774 11027 13776
rect 9121 13771 9187 13774
rect 9673 13771 9739 13774
rect 10961 13771 11027 13774
rect 11237 13834 11303 13837
rect 14457 13834 14523 13837
rect 15150 13834 15210 13910
rect 25773 13907 25839 13910
rect 11237 13832 15210 13834
rect 11237 13776 11242 13832
rect 11298 13776 14462 13832
rect 14518 13776 15210 13832
rect 11237 13774 15210 13776
rect 11237 13771 11303 13774
rect 14457 13771 14523 13774
rect 15326 13772 15332 13836
rect 15396 13834 15402 13836
rect 20478 13834 20484 13836
rect 15396 13774 20484 13834
rect 15396 13772 15402 13774
rect 20478 13772 20484 13774
rect 20548 13772 20554 13836
rect 20621 13834 20687 13837
rect 22001 13834 22067 13837
rect 20621 13832 22067 13834
rect 20621 13776 20626 13832
rect 20682 13776 22006 13832
rect 22062 13776 22067 13832
rect 20621 13774 22067 13776
rect 20621 13771 20687 13774
rect 22001 13771 22067 13774
rect 22369 13834 22435 13837
rect 25221 13834 25287 13837
rect 22369 13832 25287 13834
rect 22369 13776 22374 13832
rect 22430 13776 25226 13832
rect 25282 13776 25287 13832
rect 22369 13774 25287 13776
rect 22369 13771 22435 13774
rect 25221 13771 25287 13774
rect 0 13698 480 13728
rect 4245 13698 4311 13701
rect 0 13696 4311 13698
rect 0 13640 4250 13696
rect 4306 13640 4311 13696
rect 0 13638 4311 13640
rect 0 13608 480 13638
rect 4245 13635 4311 13638
rect 5993 13698 6059 13701
rect 9121 13698 9187 13701
rect 5993 13696 9187 13698
rect 5993 13640 5998 13696
rect 6054 13640 9126 13696
rect 9182 13640 9187 13696
rect 5993 13638 9187 13640
rect 5993 13635 6059 13638
rect 9121 13635 9187 13638
rect 10910 13636 10916 13700
rect 10980 13698 10986 13700
rect 14365 13698 14431 13701
rect 10980 13696 14431 13698
rect 10980 13640 14370 13696
rect 14426 13640 14431 13696
rect 10980 13638 14431 13640
rect 10980 13636 10986 13638
rect 14365 13635 14431 13638
rect 14590 13636 14596 13700
rect 14660 13698 14666 13700
rect 18505 13698 18571 13701
rect 14660 13696 18571 13698
rect 14660 13640 18510 13696
rect 18566 13640 18571 13696
rect 14660 13638 18571 13640
rect 14660 13636 14666 13638
rect 18505 13635 18571 13638
rect 20069 13698 20135 13701
rect 20713 13698 20779 13701
rect 26233 13698 26299 13701
rect 27520 13698 28000 13728
rect 20069 13696 20178 13698
rect 20069 13640 20074 13696
rect 20130 13640 20178 13696
rect 20069 13635 20178 13640
rect 20713 13696 26299 13698
rect 20713 13640 20718 13696
rect 20774 13640 26238 13696
rect 26294 13640 26299 13696
rect 20713 13638 26299 13640
rect 20713 13635 20779 13638
rect 26233 13635 26299 13638
rect 26374 13638 28000 13698
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 3785 13562 3851 13565
rect 8937 13562 9003 13565
rect 3785 13560 9003 13562
rect 3785 13504 3790 13560
rect 3846 13504 8942 13560
rect 8998 13504 9003 13560
rect 3785 13502 9003 13504
rect 3785 13499 3851 13502
rect 8937 13499 9003 13502
rect 10869 13562 10935 13565
rect 13813 13562 13879 13565
rect 10869 13560 13879 13562
rect 10869 13504 10874 13560
rect 10930 13504 13818 13560
rect 13874 13504 13879 13560
rect 10869 13502 13879 13504
rect 10869 13499 10935 13502
rect 13813 13499 13879 13502
rect 13997 13562 14063 13565
rect 20118 13562 20178 13635
rect 23381 13562 23447 13565
rect 13997 13560 17602 13562
rect 13997 13504 14002 13560
rect 14058 13504 17602 13560
rect 13997 13502 17602 13504
rect 20118 13560 23447 13562
rect 20118 13504 23386 13560
rect 23442 13504 23447 13560
rect 20118 13502 23447 13504
rect 13997 13499 14063 13502
rect 3785 13426 3851 13429
rect 6729 13426 6795 13429
rect 3785 13424 6795 13426
rect 3785 13368 3790 13424
rect 3846 13368 6734 13424
rect 6790 13368 6795 13424
rect 3785 13366 6795 13368
rect 3785 13363 3851 13366
rect 6729 13363 6795 13366
rect 9949 13426 10015 13429
rect 10225 13426 10291 13429
rect 17309 13426 17375 13429
rect 9949 13424 17375 13426
rect 9949 13368 9954 13424
rect 10010 13368 10230 13424
rect 10286 13368 17314 13424
rect 17370 13368 17375 13424
rect 9949 13366 17375 13368
rect 17542 13426 17602 13502
rect 23381 13499 23447 13502
rect 24669 13562 24735 13565
rect 26374 13562 26434 13638
rect 27520 13608 28000 13638
rect 24669 13560 26434 13562
rect 24669 13504 24674 13560
rect 24730 13504 26434 13560
rect 24669 13502 26434 13504
rect 24669 13499 24735 13502
rect 25773 13426 25839 13429
rect 17542 13424 25839 13426
rect 17542 13368 25778 13424
rect 25834 13368 25839 13424
rect 17542 13366 25839 13368
rect 9949 13363 10015 13366
rect 10225 13363 10291 13366
rect 17309 13363 17375 13366
rect 25773 13363 25839 13366
rect 5441 13290 5507 13293
rect 11697 13290 11763 13293
rect 14917 13290 14983 13293
rect 5441 13288 11763 13290
rect 5441 13232 5446 13288
rect 5502 13232 11702 13288
rect 11758 13232 11763 13288
rect 5441 13230 11763 13232
rect 5441 13227 5507 13230
rect 11697 13227 11763 13230
rect 11838 13288 14983 13290
rect 11838 13232 14922 13288
rect 14978 13232 14983 13288
rect 11838 13230 14983 13232
rect 0 13154 480 13184
rect 2037 13154 2103 13157
rect 5165 13154 5231 13157
rect 0 13094 1410 13154
rect 0 13064 480 13094
rect 1350 13018 1410 13094
rect 2037 13152 5231 13154
rect 2037 13096 2042 13152
rect 2098 13096 5170 13152
rect 5226 13096 5231 13152
rect 2037 13094 5231 13096
rect 2037 13091 2103 13094
rect 5165 13091 5231 13094
rect 6729 13154 6795 13157
rect 11838 13154 11898 13230
rect 14917 13227 14983 13230
rect 17493 13290 17559 13293
rect 20621 13290 20687 13293
rect 17493 13288 20687 13290
rect 17493 13232 17498 13288
rect 17554 13232 20626 13288
rect 20682 13232 20687 13288
rect 17493 13230 20687 13232
rect 17493 13227 17559 13230
rect 20621 13227 20687 13230
rect 23054 13228 23060 13292
rect 23124 13290 23130 13292
rect 24209 13290 24275 13293
rect 23124 13288 24275 13290
rect 23124 13232 24214 13288
rect 24270 13232 24275 13288
rect 23124 13230 24275 13232
rect 23124 13228 23130 13230
rect 24209 13227 24275 13230
rect 24710 13228 24716 13292
rect 24780 13290 24786 13292
rect 24853 13290 24919 13293
rect 24780 13288 24919 13290
rect 24780 13232 24858 13288
rect 24914 13232 24919 13288
rect 24780 13230 24919 13232
rect 24780 13228 24786 13230
rect 24853 13227 24919 13230
rect 25262 13228 25268 13292
rect 25332 13290 25338 13292
rect 25865 13290 25931 13293
rect 25332 13288 25931 13290
rect 25332 13232 25870 13288
rect 25926 13232 25931 13288
rect 25332 13230 25931 13232
rect 25332 13228 25338 13230
rect 25865 13227 25931 13230
rect 6729 13152 11898 13154
rect 6729 13096 6734 13152
rect 6790 13096 11898 13152
rect 6729 13094 11898 13096
rect 12065 13154 12131 13157
rect 13169 13154 13235 13157
rect 12065 13152 13235 13154
rect 12065 13096 12070 13152
rect 12126 13096 13174 13152
rect 13230 13096 13235 13152
rect 12065 13094 13235 13096
rect 6729 13091 6795 13094
rect 12065 13091 12131 13094
rect 13169 13091 13235 13094
rect 13353 13154 13419 13157
rect 13486 13154 13492 13156
rect 13353 13152 13492 13154
rect 13353 13096 13358 13152
rect 13414 13096 13492 13152
rect 13353 13094 13492 13096
rect 13353 13091 13419 13094
rect 13486 13092 13492 13094
rect 13556 13092 13562 13156
rect 15929 13154 15995 13157
rect 20805 13154 20871 13157
rect 15929 13152 20871 13154
rect 15929 13096 15934 13152
rect 15990 13096 20810 13152
rect 20866 13096 20871 13152
rect 15929 13094 20871 13096
rect 15929 13091 15995 13094
rect 20805 13091 20871 13094
rect 20989 13154 21055 13157
rect 22277 13154 22343 13157
rect 20989 13152 22343 13154
rect 20989 13096 20994 13152
rect 21050 13096 22282 13152
rect 22338 13096 22343 13152
rect 20989 13094 22343 13096
rect 20989 13091 21055 13094
rect 22277 13091 22343 13094
rect 25405 13154 25471 13157
rect 27520 13154 28000 13184
rect 25405 13152 28000 13154
rect 25405 13096 25410 13152
rect 25466 13096 28000 13152
rect 25405 13094 28000 13096
rect 25405 13091 25471 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 27520 13064 28000 13094
rect 24277 13023 24597 13024
rect 3969 13018 4035 13021
rect 1350 13016 4035 13018
rect 1350 12960 3974 13016
rect 4030 12960 4035 13016
rect 1350 12958 4035 12960
rect 3969 12955 4035 12958
rect 9990 12956 9996 13020
rect 10060 13018 10066 13020
rect 10910 13018 10916 13020
rect 10060 12958 10916 13018
rect 10060 12956 10066 12958
rect 10910 12956 10916 12958
rect 10980 12956 10986 13020
rect 11145 13018 11211 13021
rect 13537 13018 13603 13021
rect 16113 13020 16179 13021
rect 11145 13016 13603 13018
rect 11145 12960 11150 13016
rect 11206 12960 13542 13016
rect 13598 12960 13603 13016
rect 11145 12958 13603 12960
rect 11145 12955 11211 12958
rect 13537 12955 13603 12958
rect 16062 12956 16068 13020
rect 16132 13018 16179 13020
rect 18781 13018 18847 13021
rect 22737 13018 22803 13021
rect 16132 13016 16224 13018
rect 16174 12960 16224 13016
rect 16132 12958 16224 12960
rect 18781 13016 22803 13018
rect 18781 12960 18786 13016
rect 18842 12960 22742 13016
rect 22798 12960 22803 13016
rect 18781 12958 22803 12960
rect 16132 12956 16179 12958
rect 16113 12955 16179 12956
rect 18781 12955 18847 12958
rect 22737 12955 22803 12958
rect 4061 12882 4127 12885
rect 6545 12882 6611 12885
rect 8385 12882 8451 12885
rect 10041 12882 10107 12885
rect 17493 12882 17559 12885
rect 4061 12880 6611 12882
rect 4061 12824 4066 12880
rect 4122 12824 6550 12880
rect 6606 12824 6611 12880
rect 4061 12822 6611 12824
rect 4061 12819 4127 12822
rect 6545 12819 6611 12822
rect 7790 12880 9920 12882
rect 7790 12824 8390 12880
rect 8446 12824 9920 12880
rect 7790 12822 9920 12824
rect 4061 12746 4127 12749
rect 7790 12746 7850 12822
rect 8385 12819 8451 12822
rect 4061 12744 7850 12746
rect 4061 12688 4066 12744
rect 4122 12688 7850 12744
rect 4061 12686 7850 12688
rect 9860 12746 9920 12822
rect 10041 12880 17559 12882
rect 10041 12824 10046 12880
rect 10102 12824 17498 12880
rect 17554 12824 17559 12880
rect 10041 12822 17559 12824
rect 10041 12819 10107 12822
rect 17493 12819 17559 12822
rect 18505 12882 18571 12885
rect 22369 12882 22435 12885
rect 18505 12880 22435 12882
rect 18505 12824 18510 12880
rect 18566 12824 22374 12880
rect 22430 12824 22435 12880
rect 18505 12822 22435 12824
rect 18505 12819 18571 12822
rect 22369 12819 22435 12822
rect 22686 12820 22692 12884
rect 22756 12882 22762 12884
rect 25262 12882 25268 12884
rect 22756 12822 25268 12882
rect 22756 12820 22762 12822
rect 25262 12820 25268 12822
rect 25332 12820 25338 12884
rect 11145 12746 11211 12749
rect 9860 12744 11211 12746
rect 9860 12688 11150 12744
rect 11206 12688 11211 12744
rect 9860 12686 11211 12688
rect 4061 12683 4127 12686
rect 11145 12683 11211 12686
rect 11462 12684 11468 12748
rect 11532 12746 11538 12748
rect 11605 12746 11671 12749
rect 11532 12744 11671 12746
rect 11532 12688 11610 12744
rect 11666 12688 11671 12744
rect 11532 12686 11671 12688
rect 11532 12684 11538 12686
rect 11605 12683 11671 12686
rect 13169 12746 13235 12749
rect 16205 12746 16271 12749
rect 21725 12746 21791 12749
rect 13169 12744 15026 12746
rect 13169 12688 13174 12744
rect 13230 12688 15026 12744
rect 13169 12686 15026 12688
rect 13169 12683 13235 12686
rect 0 12610 480 12640
rect 3693 12610 3759 12613
rect 0 12608 3759 12610
rect 0 12552 3698 12608
rect 3754 12552 3759 12608
rect 0 12550 3759 12552
rect 0 12520 480 12550
rect 3693 12547 3759 12550
rect 5165 12610 5231 12613
rect 6361 12610 6427 12613
rect 6729 12610 6795 12613
rect 5165 12608 5964 12610
rect 5165 12552 5170 12608
rect 5226 12552 5964 12608
rect 5165 12550 5964 12552
rect 5165 12547 5231 12550
rect 2405 12474 2471 12477
rect 3601 12474 3667 12477
rect 2405 12472 3667 12474
rect 2405 12416 2410 12472
rect 2466 12416 3606 12472
rect 3662 12416 3667 12472
rect 2405 12414 3667 12416
rect 2405 12411 2471 12414
rect 3601 12411 3667 12414
rect 3785 12474 3851 12477
rect 5717 12474 5783 12477
rect 3785 12472 5783 12474
rect 3785 12416 3790 12472
rect 3846 12416 5722 12472
rect 5778 12416 5783 12472
rect 3785 12414 5783 12416
rect 5904 12474 5964 12550
rect 6361 12608 6795 12610
rect 6361 12552 6366 12608
rect 6422 12552 6734 12608
rect 6790 12552 6795 12608
rect 6361 12550 6795 12552
rect 6361 12547 6427 12550
rect 6729 12547 6795 12550
rect 10777 12610 10843 12613
rect 10910 12610 10916 12612
rect 10777 12608 10916 12610
rect 10777 12552 10782 12608
rect 10838 12552 10916 12608
rect 10777 12550 10916 12552
rect 10777 12547 10843 12550
rect 10910 12548 10916 12550
rect 10980 12548 10986 12612
rect 12065 12610 12131 12613
rect 11654 12608 12131 12610
rect 11654 12552 12070 12608
rect 12126 12552 12131 12608
rect 11654 12550 12131 12552
rect 14966 12610 15026 12686
rect 16205 12744 21791 12746
rect 16205 12688 16210 12744
rect 16266 12688 21730 12744
rect 21786 12688 21791 12744
rect 16205 12686 21791 12688
rect 16205 12683 16271 12686
rect 21725 12683 21791 12686
rect 22645 12746 22711 12749
rect 25497 12746 25563 12749
rect 22645 12744 25563 12746
rect 22645 12688 22650 12744
rect 22706 12688 25502 12744
rect 25558 12688 25563 12744
rect 22645 12686 25563 12688
rect 22645 12683 22711 12686
rect 25497 12683 25563 12686
rect 18873 12610 18939 12613
rect 14966 12608 18939 12610
rect 14966 12552 18878 12608
rect 18934 12552 18939 12608
rect 14966 12550 18939 12552
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 11513 12474 11579 12477
rect 5904 12414 10058 12474
rect 3785 12411 3851 12414
rect 5717 12411 5783 12414
rect 13 12338 79 12341
rect 1761 12338 1827 12341
rect 13 12336 1827 12338
rect 13 12280 18 12336
rect 74 12280 1766 12336
rect 1822 12280 1827 12336
rect 13 12278 1827 12280
rect 13 12275 79 12278
rect 1761 12275 1827 12278
rect 2681 12338 2747 12341
rect 5441 12338 5507 12341
rect 8293 12338 8359 12341
rect 8661 12338 8727 12341
rect 2681 12336 6930 12338
rect 2681 12280 2686 12336
rect 2742 12280 5446 12336
rect 5502 12280 6930 12336
rect 2681 12278 6930 12280
rect 2681 12275 2747 12278
rect 5441 12275 5507 12278
rect 2405 12204 2471 12205
rect 2405 12202 2452 12204
rect 2360 12200 2452 12202
rect 2360 12144 2410 12200
rect 2360 12142 2452 12144
rect 2405 12140 2452 12142
rect 2516 12140 2522 12204
rect 3969 12202 4035 12205
rect 5533 12202 5599 12205
rect 3969 12200 5599 12202
rect 3969 12144 3974 12200
rect 4030 12144 5538 12200
rect 5594 12144 5599 12200
rect 3969 12142 5599 12144
rect 2405 12139 2471 12140
rect 3969 12139 4035 12142
rect 5533 12139 5599 12142
rect 6453 12204 6519 12205
rect 6453 12200 6500 12204
rect 6564 12202 6570 12204
rect 6870 12202 6930 12278
rect 8293 12336 8727 12338
rect 8293 12280 8298 12336
rect 8354 12280 8666 12336
rect 8722 12280 8727 12336
rect 8293 12278 8727 12280
rect 9998 12338 10058 12414
rect 10734 12472 11579 12474
rect 10734 12416 11518 12472
rect 11574 12416 11579 12472
rect 10734 12414 11579 12416
rect 10734 12338 10794 12414
rect 11513 12411 11579 12414
rect 11654 12341 11714 12550
rect 12065 12547 12131 12550
rect 18873 12547 18939 12550
rect 20253 12610 20319 12613
rect 20989 12610 21055 12613
rect 20253 12608 21055 12610
rect 20253 12552 20258 12608
rect 20314 12552 20994 12608
rect 21050 12552 21055 12608
rect 20253 12550 21055 12552
rect 20253 12547 20319 12550
rect 20989 12547 21055 12550
rect 21541 12610 21607 12613
rect 21817 12610 21883 12613
rect 21541 12608 21883 12610
rect 21541 12552 21546 12608
rect 21602 12552 21822 12608
rect 21878 12552 21883 12608
rect 21541 12550 21883 12552
rect 21541 12547 21607 12550
rect 21817 12547 21883 12550
rect 23105 12610 23171 12613
rect 23565 12610 23631 12613
rect 23105 12608 23631 12610
rect 23105 12552 23110 12608
rect 23166 12552 23570 12608
rect 23626 12552 23631 12608
rect 23105 12550 23631 12552
rect 23105 12547 23171 12550
rect 23565 12547 23631 12550
rect 24209 12610 24275 12613
rect 27520 12610 28000 12640
rect 24209 12608 28000 12610
rect 24209 12552 24214 12608
rect 24270 12552 28000 12608
rect 24209 12550 28000 12552
rect 24209 12547 24275 12550
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 27520 12520 28000 12550
rect 19610 12479 19930 12480
rect 12065 12474 12131 12477
rect 14549 12474 14615 12477
rect 16430 12474 16436 12476
rect 12065 12472 14615 12474
rect 12065 12416 12070 12472
rect 12126 12416 14554 12472
rect 14610 12416 14615 12472
rect 12065 12414 14615 12416
rect 12065 12411 12131 12414
rect 14549 12411 14615 12414
rect 14736 12414 16436 12474
rect 9998 12278 10794 12338
rect 10869 12338 10935 12341
rect 10869 12336 11162 12338
rect 10869 12280 10874 12336
rect 10930 12280 11162 12336
rect 10869 12278 11162 12280
rect 11654 12336 11763 12341
rect 11654 12280 11702 12336
rect 11758 12280 11763 12336
rect 11654 12278 11763 12280
rect 8293 12275 8359 12278
rect 8661 12275 8727 12278
rect 10869 12275 10935 12278
rect 10869 12202 10935 12205
rect 6453 12144 6458 12200
rect 6453 12140 6500 12144
rect 6564 12142 6610 12202
rect 6870 12200 10935 12202
rect 6870 12144 10874 12200
rect 10930 12144 10935 12200
rect 6870 12142 10935 12144
rect 11102 12202 11162 12278
rect 11697 12275 11763 12278
rect 11881 12338 11947 12341
rect 12014 12338 12020 12340
rect 11881 12336 12020 12338
rect 11881 12280 11886 12336
rect 11942 12280 12020 12336
rect 11881 12278 12020 12280
rect 11881 12275 11947 12278
rect 12014 12276 12020 12278
rect 12084 12276 12090 12340
rect 14549 12338 14615 12341
rect 14736 12338 14796 12414
rect 16430 12412 16436 12414
rect 16500 12412 16506 12476
rect 18229 12474 18295 12477
rect 19057 12474 19123 12477
rect 18229 12472 19123 12474
rect 18229 12416 18234 12472
rect 18290 12416 19062 12472
rect 19118 12416 19123 12472
rect 18229 12414 19123 12416
rect 18229 12411 18295 12414
rect 19057 12411 19123 12414
rect 19190 12412 19196 12476
rect 19260 12474 19266 12476
rect 19333 12474 19399 12477
rect 19260 12472 19399 12474
rect 19260 12416 19338 12472
rect 19394 12416 19399 12472
rect 19260 12414 19399 12416
rect 19260 12412 19266 12414
rect 19333 12411 19399 12414
rect 20713 12474 20779 12477
rect 21449 12474 21515 12477
rect 20713 12472 21515 12474
rect 20713 12416 20718 12472
rect 20774 12416 21454 12472
rect 21510 12416 21515 12472
rect 20713 12414 21515 12416
rect 20713 12411 20779 12414
rect 21449 12411 21515 12414
rect 23381 12474 23447 12477
rect 24945 12474 25011 12477
rect 23381 12472 25011 12474
rect 23381 12416 23386 12472
rect 23442 12416 24950 12472
rect 25006 12416 25011 12472
rect 23381 12414 25011 12416
rect 23381 12411 23447 12414
rect 24945 12411 25011 12414
rect 14549 12336 14796 12338
rect 14549 12280 14554 12336
rect 14610 12280 14796 12336
rect 14549 12278 14796 12280
rect 16113 12338 16179 12341
rect 16573 12338 16639 12341
rect 24853 12338 24919 12341
rect 16113 12336 24919 12338
rect 16113 12280 16118 12336
rect 16174 12280 16578 12336
rect 16634 12280 24858 12336
rect 24914 12280 24919 12336
rect 16113 12278 24919 12280
rect 14549 12275 14615 12278
rect 16113 12275 16179 12278
rect 16573 12275 16639 12278
rect 24853 12275 24919 12278
rect 25589 12338 25655 12341
rect 25814 12338 25820 12340
rect 25589 12336 25820 12338
rect 25589 12280 25594 12336
rect 25650 12280 25820 12336
rect 25589 12278 25820 12280
rect 25589 12275 25655 12278
rect 25814 12276 25820 12278
rect 25884 12276 25890 12340
rect 13905 12202 13971 12205
rect 11102 12200 13971 12202
rect 11102 12144 13910 12200
rect 13966 12144 13971 12200
rect 11102 12142 13971 12144
rect 6564 12140 6570 12142
rect 6453 12139 6519 12140
rect 10869 12139 10935 12142
rect 13905 12139 13971 12142
rect 15377 12202 15443 12205
rect 16665 12202 16731 12205
rect 23565 12202 23631 12205
rect 15377 12200 23631 12202
rect 15377 12144 15382 12200
rect 15438 12144 16670 12200
rect 16726 12144 23570 12200
rect 23626 12144 23631 12200
rect 15377 12142 23631 12144
rect 15377 12139 15443 12142
rect 16665 12139 16731 12142
rect 23565 12139 23631 12142
rect 1945 12066 2011 12069
rect 4613 12066 4679 12069
rect 1945 12064 4679 12066
rect 1945 12008 1950 12064
rect 2006 12008 4618 12064
rect 4674 12008 4679 12064
rect 1945 12006 4679 12008
rect 1945 12003 2011 12006
rect 4613 12003 4679 12006
rect 6085 12066 6151 12069
rect 8293 12066 8359 12069
rect 6085 12064 8359 12066
rect 6085 12008 6090 12064
rect 6146 12008 8298 12064
rect 8354 12008 8359 12064
rect 6085 12006 8359 12008
rect 6085 12003 6151 12006
rect 8293 12003 8359 12006
rect 9254 12004 9260 12068
rect 9324 12066 9330 12068
rect 9949 12066 10015 12069
rect 9324 12064 10015 12066
rect 9324 12008 9954 12064
rect 10010 12008 10015 12064
rect 9324 12006 10015 12008
rect 9324 12004 9330 12006
rect 9949 12003 10015 12006
rect 15469 12066 15535 12069
rect 19977 12066 20043 12069
rect 20345 12066 20411 12069
rect 21725 12066 21791 12069
rect 15469 12064 20411 12066
rect 15469 12008 15474 12064
rect 15530 12008 19982 12064
rect 20038 12008 20350 12064
rect 20406 12008 20411 12064
rect 15469 12006 20411 12008
rect 15469 12003 15535 12006
rect 19977 12003 20043 12006
rect 20345 12003 20411 12006
rect 21222 12064 21791 12066
rect 21222 12008 21730 12064
rect 21786 12008 21791 12064
rect 21222 12006 21791 12008
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 21222 11933 21282 12006
rect 21725 12003 21791 12006
rect 23606 12004 23612 12068
rect 23676 12066 23682 12068
rect 23933 12066 23999 12069
rect 23676 12064 23999 12066
rect 23676 12008 23938 12064
rect 23994 12008 23999 12064
rect 23676 12006 23999 12008
rect 23676 12004 23682 12006
rect 23933 12003 23999 12006
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 3969 11930 4035 11933
rect 0 11928 4035 11930
rect 0 11872 3974 11928
rect 4030 11872 4035 11928
rect 0 11870 4035 11872
rect 0 11840 480 11870
rect 3969 11867 4035 11870
rect 6085 11930 6151 11933
rect 11421 11930 11487 11933
rect 6085 11928 11487 11930
rect 6085 11872 6090 11928
rect 6146 11872 11426 11928
rect 11482 11872 11487 11928
rect 6085 11870 11487 11872
rect 6085 11867 6151 11870
rect 11421 11867 11487 11870
rect 16389 11930 16455 11933
rect 21222 11930 21331 11933
rect 21449 11932 21515 11933
rect 16389 11928 21331 11930
rect 16389 11872 16394 11928
rect 16450 11872 21270 11928
rect 21326 11872 21331 11928
rect 16389 11870 21331 11872
rect 16389 11867 16455 11870
rect 21265 11867 21331 11870
rect 21398 11868 21404 11932
rect 21468 11930 21515 11932
rect 21468 11928 21560 11930
rect 21510 11872 21560 11928
rect 21468 11870 21560 11872
rect 21468 11868 21515 11870
rect 22134 11868 22140 11932
rect 22204 11930 22210 11932
rect 22369 11930 22435 11933
rect 22204 11928 22435 11930
rect 22204 11872 22374 11928
rect 22430 11872 22435 11928
rect 22204 11870 22435 11872
rect 22204 11868 22210 11870
rect 21449 11867 21515 11868
rect 22369 11867 22435 11870
rect 24761 11930 24827 11933
rect 27520 11930 28000 11960
rect 24761 11928 28000 11930
rect 24761 11872 24766 11928
rect 24822 11872 28000 11928
rect 24761 11870 28000 11872
rect 24761 11867 24827 11870
rect 27520 11840 28000 11870
rect 2221 11794 2287 11797
rect 8017 11794 8083 11797
rect 2221 11792 8083 11794
rect 2221 11736 2226 11792
rect 2282 11736 8022 11792
rect 8078 11736 8083 11792
rect 2221 11734 8083 11736
rect 2221 11731 2287 11734
rect 8017 11731 8083 11734
rect 8201 11794 8267 11797
rect 8845 11794 8911 11797
rect 12709 11794 12775 11797
rect 8201 11792 12775 11794
rect 8201 11736 8206 11792
rect 8262 11736 8850 11792
rect 8906 11736 12714 11792
rect 12770 11736 12775 11792
rect 8201 11734 12775 11736
rect 8201 11731 8267 11734
rect 8845 11731 8911 11734
rect 12709 11731 12775 11734
rect 16205 11794 16271 11797
rect 20713 11794 20779 11797
rect 26233 11794 26299 11797
rect 16205 11792 26299 11794
rect 16205 11736 16210 11792
rect 16266 11736 20718 11792
rect 20774 11736 26238 11792
rect 26294 11736 26299 11792
rect 16205 11734 26299 11736
rect 16205 11731 16271 11734
rect 20713 11731 20779 11734
rect 26233 11731 26299 11734
rect 1853 11658 1919 11661
rect 3601 11658 3667 11661
rect 4797 11658 4863 11661
rect 1853 11656 4863 11658
rect 1853 11600 1858 11656
rect 1914 11600 3606 11656
rect 3662 11600 4802 11656
rect 4858 11600 4863 11656
rect 1853 11598 4863 11600
rect 1853 11595 1919 11598
rect 3601 11595 3667 11598
rect 4797 11595 4863 11598
rect 6310 11596 6316 11660
rect 6380 11658 6386 11660
rect 6729 11658 6795 11661
rect 6380 11656 6795 11658
rect 6380 11600 6734 11656
rect 6790 11600 6795 11656
rect 6380 11598 6795 11600
rect 6380 11596 6386 11598
rect 6729 11595 6795 11598
rect 8201 11658 8267 11661
rect 10869 11658 10935 11661
rect 14181 11658 14247 11661
rect 8201 11656 10748 11658
rect 8201 11600 8206 11656
rect 8262 11600 10748 11656
rect 8201 11598 10748 11600
rect 8201 11595 8267 11598
rect 2865 11524 2931 11525
rect 2814 11460 2820 11524
rect 2884 11522 2931 11524
rect 6821 11522 6887 11525
rect 9673 11522 9739 11525
rect 2884 11520 6746 11522
rect 2926 11464 6746 11520
rect 2884 11462 6746 11464
rect 2884 11460 2931 11462
rect 2865 11459 2931 11460
rect 0 11386 480 11416
rect 3918 11386 3924 11388
rect 0 11326 3924 11386
rect 0 11296 480 11326
rect 3918 11324 3924 11326
rect 3988 11324 3994 11388
rect 6686 11386 6746 11462
rect 6821 11520 9739 11522
rect 6821 11464 6826 11520
rect 6882 11464 9678 11520
rect 9734 11464 9739 11520
rect 6821 11462 9739 11464
rect 10688 11522 10748 11598
rect 10869 11656 14247 11658
rect 10869 11600 10874 11656
rect 10930 11600 14186 11656
rect 14242 11600 14247 11656
rect 10869 11598 14247 11600
rect 10869 11595 10935 11598
rect 14181 11595 14247 11598
rect 18045 11658 18111 11661
rect 21265 11658 21331 11661
rect 18045 11656 21331 11658
rect 18045 11600 18050 11656
rect 18106 11600 21270 11656
rect 21326 11600 21331 11656
rect 18045 11598 21331 11600
rect 18045 11595 18111 11598
rect 21265 11595 21331 11598
rect 22318 11596 22324 11660
rect 22388 11658 22394 11660
rect 24669 11658 24735 11661
rect 22388 11656 24735 11658
rect 22388 11600 24674 11656
rect 24730 11600 24735 11656
rect 22388 11598 24735 11600
rect 22388 11596 22394 11598
rect 24669 11595 24735 11598
rect 13077 11522 13143 11525
rect 15469 11522 15535 11525
rect 10688 11520 15535 11522
rect 10688 11464 13082 11520
rect 13138 11464 15474 11520
rect 15530 11464 15535 11520
rect 10688 11462 15535 11464
rect 6821 11459 6887 11462
rect 9673 11459 9739 11462
rect 13077 11459 13143 11462
rect 15469 11459 15535 11462
rect 16798 11460 16804 11524
rect 16868 11522 16874 11524
rect 18781 11522 18847 11525
rect 19241 11524 19307 11525
rect 16868 11520 18847 11522
rect 16868 11464 18786 11520
rect 18842 11464 18847 11520
rect 16868 11462 18847 11464
rect 16868 11460 16874 11462
rect 18781 11459 18847 11462
rect 19190 11460 19196 11524
rect 19260 11522 19307 11524
rect 20897 11522 20963 11525
rect 24025 11522 24091 11525
rect 19260 11520 19352 11522
rect 19302 11464 19352 11520
rect 19260 11462 19352 11464
rect 20897 11520 24091 11522
rect 20897 11464 20902 11520
rect 20958 11464 24030 11520
rect 24086 11464 24091 11520
rect 20897 11462 24091 11464
rect 19260 11460 19307 11462
rect 19241 11459 19307 11460
rect 20897 11459 20963 11462
rect 24025 11459 24091 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 9581 11386 9647 11389
rect 6686 11384 9647 11386
rect 6686 11328 9586 11384
rect 9642 11328 9647 11384
rect 6686 11326 9647 11328
rect 9581 11323 9647 11326
rect 10777 11386 10843 11389
rect 13445 11386 13511 11389
rect 14273 11386 14339 11389
rect 10777 11384 14339 11386
rect 10777 11328 10782 11384
rect 10838 11328 13450 11384
rect 13506 11328 14278 11384
rect 14334 11328 14339 11384
rect 10777 11326 14339 11328
rect 10777 11323 10843 11326
rect 13445 11323 13511 11326
rect 14273 11323 14339 11326
rect 14590 11324 14596 11388
rect 14660 11386 14666 11388
rect 14825 11386 14891 11389
rect 14660 11384 14891 11386
rect 14660 11328 14830 11384
rect 14886 11328 14891 11384
rect 14660 11326 14891 11328
rect 14660 11324 14666 11326
rect 14825 11323 14891 11326
rect 15285 11386 15351 11389
rect 15510 11386 15516 11388
rect 15285 11384 15516 11386
rect 15285 11328 15290 11384
rect 15346 11328 15516 11384
rect 15285 11326 15516 11328
rect 15285 11323 15351 11326
rect 15510 11324 15516 11326
rect 15580 11324 15586 11388
rect 16757 11386 16823 11389
rect 20713 11386 20779 11389
rect 21950 11386 21956 11388
rect 16757 11384 18154 11386
rect 16757 11328 16762 11384
rect 16818 11328 18154 11384
rect 16757 11326 18154 11328
rect 16757 11323 16823 11326
rect 2037 11250 2103 11253
rect 7741 11250 7807 11253
rect 2037 11248 7807 11250
rect 2037 11192 2042 11248
rect 2098 11192 7746 11248
rect 7802 11192 7807 11248
rect 2037 11190 7807 11192
rect 2037 11187 2103 11190
rect 7741 11187 7807 11190
rect 8293 11250 8359 11253
rect 10133 11250 10199 11253
rect 8293 11248 10199 11250
rect 8293 11192 8298 11248
rect 8354 11192 10138 11248
rect 10194 11192 10199 11248
rect 8293 11190 10199 11192
rect 8293 11187 8359 11190
rect 10133 11187 10199 11190
rect 10777 11250 10843 11253
rect 11278 11250 11284 11252
rect 10777 11248 11284 11250
rect 10777 11192 10782 11248
rect 10838 11192 11284 11248
rect 10777 11190 11284 11192
rect 10777 11187 10843 11190
rect 11278 11188 11284 11190
rect 11348 11188 11354 11252
rect 11421 11250 11487 11253
rect 12985 11250 13051 11253
rect 11421 11248 13051 11250
rect 11421 11192 11426 11248
rect 11482 11192 12990 11248
rect 13046 11192 13051 11248
rect 11421 11190 13051 11192
rect 11421 11187 11487 11190
rect 12985 11187 13051 11190
rect 13629 11250 13695 11253
rect 17953 11250 18019 11253
rect 13629 11248 18019 11250
rect 13629 11192 13634 11248
rect 13690 11192 17958 11248
rect 18014 11192 18019 11248
rect 13629 11190 18019 11192
rect 18094 11250 18154 11326
rect 20713 11384 21956 11386
rect 20713 11328 20718 11384
rect 20774 11328 21956 11384
rect 20713 11326 21956 11328
rect 20713 11323 20779 11326
rect 21950 11324 21956 11326
rect 22020 11324 22026 11388
rect 22185 11386 22251 11389
rect 27520 11386 28000 11416
rect 22185 11384 28000 11386
rect 22185 11328 22190 11384
rect 22246 11328 28000 11384
rect 22185 11326 28000 11328
rect 22185 11323 22251 11326
rect 27520 11296 28000 11326
rect 18321 11250 18387 11253
rect 21817 11250 21883 11253
rect 18094 11248 21883 11250
rect 18094 11192 18326 11248
rect 18382 11192 21822 11248
rect 21878 11192 21883 11248
rect 18094 11190 21883 11192
rect 13629 11187 13695 11190
rect 17953 11187 18019 11190
rect 18321 11187 18387 11190
rect 21817 11187 21883 11190
rect 3918 11052 3924 11116
rect 3988 11114 3994 11116
rect 10961 11114 11027 11117
rect 14733 11114 14799 11117
rect 3988 11054 9690 11114
rect 3988 11052 3994 11054
rect 1485 10978 1551 10981
rect 3509 10978 3575 10981
rect 1485 10976 3575 10978
rect 1485 10920 1490 10976
rect 1546 10920 3514 10976
rect 3570 10920 3575 10976
rect 1485 10918 3575 10920
rect 9630 10978 9690 11054
rect 10961 11112 14799 11114
rect 10961 11056 10966 11112
rect 11022 11056 14738 11112
rect 14794 11056 14799 11112
rect 10961 11054 14799 11056
rect 10961 11051 11027 11054
rect 14733 11051 14799 11054
rect 16982 11052 16988 11116
rect 17052 11114 17058 11116
rect 17125 11114 17191 11117
rect 17052 11112 17191 11114
rect 17052 11056 17130 11112
rect 17186 11056 17191 11112
rect 17052 11054 17191 11056
rect 17052 11052 17058 11054
rect 17125 11051 17191 11054
rect 19374 11052 19380 11116
rect 19444 11114 19450 11116
rect 19517 11114 19583 11117
rect 21357 11114 21423 11117
rect 23473 11114 23539 11117
rect 19444 11112 19583 11114
rect 19444 11056 19522 11112
rect 19578 11056 19583 11112
rect 19444 11054 19583 11056
rect 19444 11052 19450 11054
rect 19517 11051 19583 11054
rect 20118 11054 21282 11114
rect 12525 10978 12591 10981
rect 13629 10978 13695 10981
rect 9630 10976 13695 10978
rect 9630 10920 12530 10976
rect 12586 10920 13634 10976
rect 13690 10920 13695 10976
rect 9630 10918 13695 10920
rect 1485 10915 1551 10918
rect 3509 10915 3575 10918
rect 12525 10915 12591 10918
rect 13629 10915 13695 10918
rect 15653 10978 15719 10981
rect 19793 10978 19859 10981
rect 15653 10976 19859 10978
rect 15653 10920 15658 10976
rect 15714 10920 19798 10976
rect 19854 10920 19859 10976
rect 15653 10918 19859 10920
rect 15653 10915 15719 10918
rect 19793 10915 19859 10918
rect 5610 10912 5930 10913
rect 0 10842 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 7281 10842 7347 10845
rect 11881 10842 11947 10845
rect 0 10782 4906 10842
rect 0 10752 480 10782
rect 2037 10572 2103 10573
rect 2037 10570 2084 10572
rect 1992 10568 2084 10570
rect 1992 10512 2042 10568
rect 1992 10510 2084 10512
rect 2037 10508 2084 10510
rect 2148 10508 2154 10572
rect 4846 10570 4906 10782
rect 7281 10840 11947 10842
rect 7281 10784 7286 10840
rect 7342 10784 11886 10840
rect 11942 10784 11947 10840
rect 7281 10782 11947 10784
rect 7281 10779 7347 10782
rect 11881 10779 11947 10782
rect 12525 10842 12591 10845
rect 14457 10842 14523 10845
rect 12525 10840 14523 10842
rect 12525 10784 12530 10840
rect 12586 10784 14462 10840
rect 14518 10784 14523 10840
rect 12525 10782 14523 10784
rect 12525 10779 12591 10782
rect 14457 10779 14523 10782
rect 16021 10842 16087 10845
rect 18965 10842 19031 10845
rect 20118 10842 20178 11054
rect 21222 10978 21282 11054
rect 21357 11112 23539 11114
rect 21357 11056 21362 11112
rect 21418 11056 23478 11112
rect 23534 11056 23539 11112
rect 21357 11054 23539 11056
rect 21357 11051 21423 11054
rect 23473 11051 23539 11054
rect 25037 10980 25103 10981
rect 21222 10918 24042 10978
rect 16021 10840 20178 10842
rect 16021 10784 16026 10840
rect 16082 10784 18970 10840
rect 19026 10784 20178 10840
rect 16021 10782 20178 10784
rect 20345 10842 20411 10845
rect 20478 10842 20484 10844
rect 20345 10840 20484 10842
rect 20345 10784 20350 10840
rect 20406 10784 20484 10840
rect 20345 10782 20484 10784
rect 16021 10779 16087 10782
rect 18965 10779 19031 10782
rect 20345 10779 20411 10782
rect 20478 10780 20484 10782
rect 20548 10780 20554 10844
rect 5165 10706 5231 10709
rect 7649 10706 7715 10709
rect 5165 10704 7715 10706
rect 5165 10648 5170 10704
rect 5226 10648 7654 10704
rect 7710 10648 7715 10704
rect 5165 10646 7715 10648
rect 5165 10643 5231 10646
rect 7649 10643 7715 10646
rect 7925 10706 7991 10709
rect 11053 10706 11119 10709
rect 12709 10706 12775 10709
rect 7925 10704 12775 10706
rect 7925 10648 7930 10704
rect 7986 10648 11058 10704
rect 11114 10648 12714 10704
rect 12770 10648 12775 10704
rect 7925 10646 12775 10648
rect 7925 10643 7991 10646
rect 11053 10643 11119 10646
rect 12709 10643 12775 10646
rect 13537 10706 13603 10709
rect 15745 10706 15811 10709
rect 21817 10706 21883 10709
rect 13537 10704 21883 10706
rect 13537 10648 13542 10704
rect 13598 10648 15750 10704
rect 15806 10648 21822 10704
rect 21878 10648 21883 10704
rect 13537 10646 21883 10648
rect 13537 10643 13603 10646
rect 15745 10643 15811 10646
rect 21817 10643 21883 10646
rect 22277 10706 22343 10709
rect 23565 10706 23631 10709
rect 22277 10704 23631 10706
rect 22277 10648 22282 10704
rect 22338 10648 23570 10704
rect 23626 10648 23631 10704
rect 22277 10646 23631 10648
rect 23982 10706 24042 10918
rect 25037 10976 25084 10980
rect 25148 10978 25154 10980
rect 25589 10978 25655 10981
rect 26366 10978 26372 10980
rect 25037 10920 25042 10976
rect 25037 10916 25084 10920
rect 25148 10918 25194 10978
rect 25589 10976 26372 10978
rect 25589 10920 25594 10976
rect 25650 10920 26372 10976
rect 25589 10918 26372 10920
rect 25148 10916 25154 10918
rect 25037 10915 25103 10916
rect 25589 10915 25655 10918
rect 26366 10916 26372 10918
rect 26436 10916 26442 10980
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 27520 10842 28000 10872
rect 24718 10782 28000 10842
rect 24718 10706 24778 10782
rect 27520 10752 28000 10782
rect 23982 10646 24778 10706
rect 22277 10643 22343 10646
rect 23565 10643 23631 10646
rect 16205 10570 16271 10573
rect 4846 10568 16271 10570
rect 4846 10512 16210 10568
rect 16266 10512 16271 10568
rect 4846 10510 16271 10512
rect 2037 10507 2103 10508
rect 16205 10507 16271 10510
rect 16757 10570 16823 10573
rect 22461 10570 22527 10573
rect 16757 10568 22527 10570
rect 16757 10512 16762 10568
rect 16818 10512 22466 10568
rect 22522 10512 22527 10568
rect 16757 10510 22527 10512
rect 16757 10507 16823 10510
rect 22461 10507 22527 10510
rect 23749 10570 23815 10573
rect 25957 10570 26023 10573
rect 23749 10568 26023 10570
rect 23749 10512 23754 10568
rect 23810 10512 25962 10568
rect 26018 10512 26023 10568
rect 23749 10510 26023 10512
rect 23749 10507 23815 10510
rect 25957 10507 26023 10510
rect 3509 10434 3575 10437
rect 5901 10434 5967 10437
rect 3509 10432 5967 10434
rect 3509 10376 3514 10432
rect 3570 10376 5906 10432
rect 5962 10376 5967 10432
rect 3509 10374 5967 10376
rect 3509 10371 3575 10374
rect 5901 10371 5967 10374
rect 10869 10434 10935 10437
rect 13813 10434 13879 10437
rect 10869 10432 13879 10434
rect 10869 10376 10874 10432
rect 10930 10376 13818 10432
rect 13874 10376 13879 10432
rect 10869 10374 13879 10376
rect 10869 10371 10935 10374
rect 13813 10371 13879 10374
rect 14457 10434 14523 10437
rect 15653 10434 15719 10437
rect 14457 10432 15719 10434
rect 14457 10376 14462 10432
rect 14518 10376 15658 10432
rect 15714 10376 15719 10432
rect 14457 10374 15719 10376
rect 14457 10371 14523 10374
rect 15653 10371 15719 10374
rect 16205 10434 16271 10437
rect 17861 10434 17927 10437
rect 16205 10432 17927 10434
rect 16205 10376 16210 10432
rect 16266 10376 17866 10432
rect 17922 10376 17927 10432
rect 16205 10374 17927 10376
rect 16205 10371 16271 10374
rect 17861 10371 17927 10374
rect 21725 10434 21791 10437
rect 25773 10434 25839 10437
rect 21725 10432 25839 10434
rect 21725 10376 21730 10432
rect 21786 10376 25778 10432
rect 25834 10376 25839 10432
rect 21725 10374 25839 10376
rect 21725 10371 21791 10374
rect 25773 10371 25839 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 2313 10298 2379 10301
rect 6453 10298 6519 10301
rect 2313 10296 6519 10298
rect 2313 10240 2318 10296
rect 2374 10240 6458 10296
rect 6514 10240 6519 10296
rect 2313 10238 6519 10240
rect 2313 10235 2379 10238
rect 6453 10235 6519 10238
rect 10910 10236 10916 10300
rect 10980 10298 10986 10300
rect 11053 10298 11119 10301
rect 10980 10296 11119 10298
rect 10980 10240 11058 10296
rect 11114 10240 11119 10296
rect 10980 10238 11119 10240
rect 10980 10236 10986 10238
rect 11053 10235 11119 10238
rect 11605 10298 11671 10301
rect 15285 10298 15351 10301
rect 11605 10296 15351 10298
rect 11605 10240 11610 10296
rect 11666 10240 15290 10296
rect 15346 10240 15351 10296
rect 11605 10238 15351 10240
rect 11605 10235 11671 10238
rect 15285 10235 15351 10238
rect 15653 10298 15719 10301
rect 16021 10298 16087 10301
rect 15653 10296 16087 10298
rect 15653 10240 15658 10296
rect 15714 10240 16026 10296
rect 16082 10240 16087 10296
rect 15653 10238 16087 10240
rect 15653 10235 15719 10238
rect 16021 10235 16087 10238
rect 16941 10298 17007 10301
rect 19425 10298 19491 10301
rect 16941 10296 19491 10298
rect 16941 10240 16946 10296
rect 17002 10240 19430 10296
rect 19486 10240 19491 10296
rect 16941 10238 19491 10240
rect 16941 10235 17007 10238
rect 19425 10235 19491 10238
rect 20294 10236 20300 10300
rect 20364 10298 20370 10300
rect 20437 10298 20503 10301
rect 20364 10296 20503 10298
rect 20364 10240 20442 10296
rect 20498 10240 20503 10296
rect 20364 10238 20503 10240
rect 20364 10236 20370 10238
rect 20437 10235 20503 10238
rect 0 10162 480 10192
rect 5533 10162 5599 10165
rect 0 10160 5599 10162
rect 0 10104 5538 10160
rect 5594 10104 5599 10160
rect 0 10102 5599 10104
rect 0 10072 480 10102
rect 5533 10099 5599 10102
rect 5809 10162 5875 10165
rect 12157 10162 12223 10165
rect 5809 10160 12223 10162
rect 5809 10104 5814 10160
rect 5870 10104 12162 10160
rect 12218 10104 12223 10160
rect 5809 10102 12223 10104
rect 5809 10099 5875 10102
rect 12157 10099 12223 10102
rect 14181 10162 14247 10165
rect 16021 10162 16087 10165
rect 18873 10162 18939 10165
rect 14181 10160 18939 10162
rect 14181 10104 14186 10160
rect 14242 10104 16026 10160
rect 16082 10104 18878 10160
rect 18934 10104 18939 10160
rect 14181 10102 18939 10104
rect 14181 10099 14247 10102
rect 16021 10099 16087 10102
rect 18873 10099 18939 10102
rect 19057 10162 19123 10165
rect 21541 10162 21607 10165
rect 19057 10160 21607 10162
rect 19057 10104 19062 10160
rect 19118 10104 21546 10160
rect 21602 10104 21607 10160
rect 19057 10102 21607 10104
rect 19057 10099 19123 10102
rect 21541 10099 21607 10102
rect 21817 10162 21883 10165
rect 22921 10162 22987 10165
rect 21817 10160 22987 10162
rect 21817 10104 21822 10160
rect 21878 10104 22926 10160
rect 22982 10104 22987 10160
rect 21817 10102 22987 10104
rect 21817 10099 21883 10102
rect 22921 10099 22987 10102
rect 23473 10162 23539 10165
rect 27520 10162 28000 10192
rect 23473 10160 28000 10162
rect 23473 10104 23478 10160
rect 23534 10104 28000 10160
rect 23473 10102 28000 10104
rect 23473 10099 23539 10102
rect 27520 10072 28000 10102
rect 1393 10026 1459 10029
rect 7649 10026 7715 10029
rect 11329 10026 11395 10029
rect 15326 10026 15332 10028
rect 1393 10024 7528 10026
rect 1393 9968 1398 10024
rect 1454 9968 7528 10024
rect 1393 9966 7528 9968
rect 1393 9963 1459 9966
rect 5349 9892 5415 9893
rect 5349 9890 5396 9892
rect 5304 9888 5396 9890
rect 5304 9832 5354 9888
rect 5304 9830 5396 9832
rect 5349 9828 5396 9830
rect 5460 9828 5466 9892
rect 6361 9890 6427 9893
rect 6678 9890 6684 9892
rect 6361 9888 6684 9890
rect 6361 9832 6366 9888
rect 6422 9832 6684 9888
rect 6361 9830 6684 9832
rect 5349 9827 5415 9828
rect 6361 9827 6427 9830
rect 6678 9828 6684 9830
rect 6748 9828 6754 9892
rect 7468 9890 7528 9966
rect 7649 10024 11395 10026
rect 7649 9968 7654 10024
rect 7710 9968 11334 10024
rect 11390 9968 11395 10024
rect 7649 9966 11395 9968
rect 7649 9963 7715 9966
rect 11329 9963 11395 9966
rect 14230 9966 15332 10026
rect 10133 9890 10199 9893
rect 10593 9890 10659 9893
rect 7468 9888 10659 9890
rect 7468 9832 10138 9888
rect 10194 9832 10598 9888
rect 10654 9832 10659 9888
rect 7468 9830 10659 9832
rect 10133 9827 10199 9830
rect 10593 9827 10659 9830
rect 10961 9890 11027 9893
rect 12893 9890 12959 9893
rect 10961 9888 12959 9890
rect 10961 9832 10966 9888
rect 11022 9832 12898 9888
rect 12954 9832 12959 9888
rect 10961 9830 12959 9832
rect 10961 9827 11027 9830
rect 12893 9827 12959 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 3233 9754 3299 9757
rect 4521 9754 4587 9757
rect 3233 9752 4587 9754
rect 3233 9696 3238 9752
rect 3294 9696 4526 9752
rect 4582 9696 4587 9752
rect 3233 9694 4587 9696
rect 3233 9691 3299 9694
rect 4521 9691 4587 9694
rect 7557 9754 7623 9757
rect 7782 9754 7788 9756
rect 7557 9752 7788 9754
rect 7557 9696 7562 9752
rect 7618 9696 7788 9752
rect 7557 9694 7788 9696
rect 7557 9691 7623 9694
rect 7782 9692 7788 9694
rect 7852 9692 7858 9756
rect 10593 9754 10659 9757
rect 14230 9754 14290 9966
rect 15326 9964 15332 9966
rect 15396 9964 15402 10028
rect 16389 10026 16455 10029
rect 18045 10026 18111 10029
rect 23289 10026 23355 10029
rect 16389 10024 23355 10026
rect 16389 9968 16394 10024
rect 16450 9968 18050 10024
rect 18106 9968 23294 10024
rect 23350 9968 23355 10024
rect 16389 9966 23355 9968
rect 16389 9963 16455 9966
rect 18045 9963 18111 9966
rect 23289 9963 23355 9966
rect 23565 10026 23631 10029
rect 25313 10026 25379 10029
rect 23565 10024 25379 10026
rect 23565 9968 23570 10024
rect 23626 9968 25318 10024
rect 25374 9968 25379 10024
rect 23565 9966 25379 9968
rect 23565 9963 23631 9966
rect 25313 9963 25379 9966
rect 16849 9890 16915 9893
rect 23289 9890 23355 9893
rect 16849 9888 23355 9890
rect 16849 9832 16854 9888
rect 16910 9832 23294 9888
rect 23350 9832 23355 9888
rect 16849 9830 23355 9832
rect 16849 9827 16915 9830
rect 23289 9827 23355 9830
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 10593 9752 14290 9754
rect 10593 9696 10598 9752
rect 10654 9696 14290 9752
rect 10593 9694 14290 9696
rect 18413 9754 18479 9757
rect 20713 9754 20779 9757
rect 18413 9752 20779 9754
rect 18413 9696 18418 9752
rect 18474 9696 20718 9752
rect 20774 9696 20779 9752
rect 18413 9694 20779 9696
rect 10593 9691 10659 9694
rect 18413 9691 18479 9694
rect 20713 9691 20779 9694
rect 21633 9754 21699 9757
rect 24025 9754 24091 9757
rect 21633 9752 24091 9754
rect 21633 9696 21638 9752
rect 21694 9696 24030 9752
rect 24086 9696 24091 9752
rect 21633 9694 24091 9696
rect 21633 9691 21699 9694
rect 24025 9691 24091 9694
rect 0 9618 480 9648
rect 1393 9618 1459 9621
rect 1761 9620 1827 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 480 9558
rect 1393 9555 1459 9558
rect 1710 9556 1716 9620
rect 1780 9618 1827 9620
rect 3693 9618 3759 9621
rect 4153 9618 4219 9621
rect 1780 9616 1872 9618
rect 1822 9560 1872 9616
rect 1780 9558 1872 9560
rect 3693 9616 4219 9618
rect 3693 9560 3698 9616
rect 3754 9560 4158 9616
rect 4214 9560 4219 9616
rect 3693 9558 4219 9560
rect 1780 9556 1827 9558
rect 1761 9555 1827 9556
rect 3693 9555 3759 9558
rect 4153 9555 4219 9558
rect 4705 9618 4771 9621
rect 8017 9618 8083 9621
rect 4705 9616 8083 9618
rect 4705 9560 4710 9616
rect 4766 9560 8022 9616
rect 8078 9560 8083 9616
rect 4705 9558 8083 9560
rect 4705 9555 4771 9558
rect 8017 9555 8083 9558
rect 9489 9618 9555 9621
rect 21449 9618 21515 9621
rect 9489 9616 21515 9618
rect 9489 9560 9494 9616
rect 9550 9560 21454 9616
rect 21510 9560 21515 9616
rect 9489 9558 21515 9560
rect 9489 9555 9555 9558
rect 21449 9555 21515 9558
rect 21817 9618 21883 9621
rect 22921 9618 22987 9621
rect 21817 9616 22987 9618
rect 21817 9560 21822 9616
rect 21878 9560 22926 9616
rect 22982 9560 22987 9616
rect 21817 9558 22987 9560
rect 21817 9555 21883 9558
rect 22921 9555 22987 9558
rect 23422 9556 23428 9620
rect 23492 9618 23498 9620
rect 23657 9618 23723 9621
rect 23492 9616 23723 9618
rect 23492 9560 23662 9616
rect 23718 9560 23723 9616
rect 23492 9558 23723 9560
rect 23492 9556 23498 9558
rect 23657 9555 23723 9558
rect 24894 9556 24900 9620
rect 24964 9618 24970 9620
rect 25037 9618 25103 9621
rect 24964 9616 25103 9618
rect 24964 9560 25042 9616
rect 25098 9560 25103 9616
rect 24964 9558 25103 9560
rect 24964 9556 24970 9558
rect 25037 9555 25103 9558
rect 25405 9620 25471 9621
rect 25957 9620 26023 9621
rect 25405 9616 25452 9620
rect 25516 9618 25522 9620
rect 25405 9560 25410 9616
rect 25405 9556 25452 9560
rect 25516 9558 25562 9618
rect 25957 9616 26004 9620
rect 26068 9618 26074 9620
rect 27520 9618 28000 9648
rect 25957 9560 25962 9616
rect 25516 9556 25522 9558
rect 25957 9556 26004 9560
rect 26068 9558 26114 9618
rect 26190 9558 28000 9618
rect 26068 9556 26074 9558
rect 25405 9555 25471 9556
rect 25957 9555 26023 9556
rect 2129 9482 2195 9485
rect 6177 9482 6243 9485
rect 2129 9480 6243 9482
rect 2129 9424 2134 9480
rect 2190 9424 6182 9480
rect 6238 9424 6243 9480
rect 9673 9480 9739 9485
rect 9673 9448 9678 9480
rect 2129 9422 6243 9424
rect 2129 9419 2195 9422
rect 6177 9419 6243 9422
rect 9492 9424 9678 9448
rect 9734 9424 9739 9480
rect 9492 9419 9739 9424
rect 10593 9482 10659 9485
rect 11094 9482 11100 9484
rect 10593 9480 11100 9482
rect 10593 9424 10598 9480
rect 10654 9424 11100 9480
rect 10593 9422 11100 9424
rect 10593 9419 10659 9422
rect 11094 9420 11100 9422
rect 11164 9420 11170 9484
rect 13997 9482 14063 9485
rect 19149 9482 19215 9485
rect 13997 9480 19215 9482
rect 13997 9424 14002 9480
rect 14058 9424 19154 9480
rect 19210 9424 19215 9480
rect 13997 9422 19215 9424
rect 13997 9419 14063 9422
rect 19149 9419 19215 9422
rect 23565 9482 23631 9485
rect 23565 9480 25146 9482
rect 23565 9424 23570 9480
rect 23626 9424 25146 9480
rect 23565 9422 25146 9424
rect 23565 9419 23631 9422
rect 9492 9388 9736 9419
rect 2037 9346 2103 9349
rect 9492 9346 9552 9388
rect 2037 9344 9552 9346
rect 2037 9288 2042 9344
rect 2098 9288 9552 9344
rect 2037 9286 9552 9288
rect 14273 9346 14339 9349
rect 14406 9346 14412 9348
rect 14273 9344 14412 9346
rect 14273 9288 14278 9344
rect 14334 9288 14412 9344
rect 14273 9286 14412 9288
rect 2037 9283 2103 9286
rect 14273 9283 14339 9286
rect 14406 9284 14412 9286
rect 14476 9284 14482 9348
rect 14917 9346 14983 9349
rect 19425 9346 19491 9349
rect 14917 9344 19491 9346
rect 14917 9288 14922 9344
rect 14978 9288 19430 9344
rect 19486 9288 19491 9344
rect 14917 9286 19491 9288
rect 14917 9283 14983 9286
rect 19425 9283 19491 9286
rect 20529 9346 20595 9349
rect 23473 9346 23539 9349
rect 20529 9344 23539 9346
rect 20529 9288 20534 9344
rect 20590 9288 23478 9344
rect 23534 9288 23539 9344
rect 20529 9286 23539 9288
rect 25086 9346 25146 9422
rect 25262 9420 25268 9484
rect 25332 9482 25338 9484
rect 25773 9482 25839 9485
rect 25332 9480 25839 9482
rect 25332 9424 25778 9480
rect 25834 9424 25839 9480
rect 25332 9422 25839 9424
rect 25332 9420 25338 9422
rect 25773 9419 25839 9422
rect 26190 9346 26250 9558
rect 27520 9528 28000 9558
rect 25086 9286 26250 9346
rect 20529 9283 20595 9286
rect 23473 9283 23539 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 2405 9210 2471 9213
rect 2998 9210 3004 9212
rect 2405 9208 3004 9210
rect 2405 9152 2410 9208
rect 2466 9152 3004 9208
rect 2405 9150 3004 9152
rect 2405 9147 2471 9150
rect 2998 9148 3004 9150
rect 3068 9148 3074 9212
rect 3417 9210 3483 9213
rect 5901 9210 5967 9213
rect 3417 9208 5967 9210
rect 3417 9152 3422 9208
rect 3478 9152 5906 9208
rect 5962 9152 5967 9208
rect 3417 9150 5967 9152
rect 3417 9147 3483 9150
rect 5901 9147 5967 9150
rect 6177 9210 6243 9213
rect 9622 9210 9628 9212
rect 6177 9208 9628 9210
rect 6177 9152 6182 9208
rect 6238 9152 9628 9208
rect 6177 9150 9628 9152
rect 6177 9147 6243 9150
rect 9622 9148 9628 9150
rect 9692 9148 9698 9212
rect 10910 9148 10916 9212
rect 10980 9210 10986 9212
rect 11053 9210 11119 9213
rect 10980 9208 11119 9210
rect 10980 9152 11058 9208
rect 11114 9152 11119 9208
rect 10980 9150 11119 9152
rect 10980 9148 10986 9150
rect 11053 9147 11119 9150
rect 12433 9210 12499 9213
rect 18781 9210 18847 9213
rect 12433 9208 18847 9210
rect 12433 9152 12438 9208
rect 12494 9152 18786 9208
rect 18842 9152 18847 9208
rect 12433 9150 18847 9152
rect 12433 9147 12499 9150
rect 18781 9147 18847 9150
rect 20662 9148 20668 9212
rect 20732 9210 20738 9212
rect 21265 9210 21331 9213
rect 20732 9208 21331 9210
rect 20732 9152 21270 9208
rect 21326 9152 21331 9208
rect 20732 9150 21331 9152
rect 20732 9148 20738 9150
rect 21265 9147 21331 9150
rect 26233 9210 26299 9213
rect 26734 9210 26740 9212
rect 26233 9208 26740 9210
rect 26233 9152 26238 9208
rect 26294 9152 26740 9208
rect 26233 9150 26740 9152
rect 26233 9147 26299 9150
rect 26734 9148 26740 9150
rect 26804 9148 26810 9212
rect 0 9074 480 9104
rect 2129 9074 2195 9077
rect 5809 9074 5875 9077
rect 0 9014 2008 9074
rect 0 8984 480 9014
rect 1948 8938 2008 9014
rect 2129 9072 5875 9074
rect 2129 9016 2134 9072
rect 2190 9016 5814 9072
rect 5870 9016 5875 9072
rect 2129 9014 5875 9016
rect 2129 9011 2195 9014
rect 5809 9011 5875 9014
rect 7649 9074 7715 9077
rect 13169 9074 13235 9077
rect 7649 9072 13235 9074
rect 7649 9016 7654 9072
rect 7710 9016 13174 9072
rect 13230 9016 13235 9072
rect 7649 9014 13235 9016
rect 7649 9011 7715 9014
rect 13169 9011 13235 9014
rect 13721 9074 13787 9077
rect 15745 9074 15811 9077
rect 13721 9072 15811 9074
rect 13721 9016 13726 9072
rect 13782 9016 15750 9072
rect 15806 9016 15811 9072
rect 13721 9014 15811 9016
rect 13721 9011 13787 9014
rect 15745 9011 15811 9014
rect 16297 9074 16363 9077
rect 21173 9074 21239 9077
rect 16297 9072 21239 9074
rect 16297 9016 16302 9072
rect 16358 9016 21178 9072
rect 21234 9016 21239 9072
rect 16297 9014 21239 9016
rect 16297 9011 16363 9014
rect 21173 9011 21239 9014
rect 21357 9074 21423 9077
rect 23473 9074 23539 9077
rect 21357 9072 23539 9074
rect 21357 9016 21362 9072
rect 21418 9016 23478 9072
rect 23534 9016 23539 9072
rect 21357 9014 23539 9016
rect 21357 9011 21423 9014
rect 23473 9011 23539 9014
rect 23749 9074 23815 9077
rect 27520 9074 28000 9104
rect 23749 9072 28000 9074
rect 23749 9016 23754 9072
rect 23810 9016 28000 9072
rect 23749 9014 28000 9016
rect 23749 9011 23815 9014
rect 27520 8984 28000 9014
rect 2865 8938 2931 8941
rect 1948 8936 2931 8938
rect 1948 8880 2870 8936
rect 2926 8880 2931 8936
rect 1948 8878 2931 8880
rect 2865 8875 2931 8878
rect 3785 8938 3851 8941
rect 4061 8938 4127 8941
rect 6177 8938 6243 8941
rect 14089 8938 14155 8941
rect 19425 8938 19491 8941
rect 3785 8936 6056 8938
rect 3785 8880 3790 8936
rect 3846 8880 4066 8936
rect 4122 8880 6056 8936
rect 3785 8878 6056 8880
rect 3785 8875 3851 8878
rect 4061 8875 4127 8878
rect 1945 8802 2011 8805
rect 4838 8802 4844 8804
rect 1945 8800 4844 8802
rect 1945 8744 1950 8800
rect 2006 8744 4844 8800
rect 1945 8742 4844 8744
rect 1945 8739 2011 8742
rect 4838 8740 4844 8742
rect 4908 8740 4914 8804
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 3325 8666 3391 8669
rect 4705 8666 4771 8669
rect 3325 8664 4771 8666
rect 3325 8608 3330 8664
rect 3386 8608 4710 8664
rect 4766 8608 4771 8664
rect 3325 8606 4771 8608
rect 5996 8666 6056 8878
rect 6177 8936 14155 8938
rect 6177 8880 6182 8936
rect 6238 8880 14094 8936
rect 14150 8880 14155 8936
rect 6177 8878 14155 8880
rect 6177 8875 6243 8878
rect 14089 8875 14155 8878
rect 14782 8936 19491 8938
rect 14782 8880 19430 8936
rect 19486 8880 19491 8936
rect 14782 8878 19491 8880
rect 9397 8802 9463 8805
rect 14782 8802 14842 8878
rect 19425 8875 19491 8878
rect 19609 8938 19675 8941
rect 20110 8938 20116 8940
rect 19609 8936 20116 8938
rect 19609 8880 19614 8936
rect 19670 8880 20116 8936
rect 19609 8878 20116 8880
rect 19609 8875 19675 8878
rect 20110 8876 20116 8878
rect 20180 8876 20186 8940
rect 20897 8938 20963 8941
rect 26417 8938 26483 8941
rect 20897 8936 26483 8938
rect 20897 8880 20902 8936
rect 20958 8880 26422 8936
rect 26478 8880 26483 8936
rect 20897 8878 26483 8880
rect 20897 8875 20963 8878
rect 26417 8875 26483 8878
rect 17493 8802 17559 8805
rect 9397 8800 14842 8802
rect 9397 8744 9402 8800
rect 9458 8744 14842 8800
rect 9397 8742 14842 8744
rect 15334 8800 17559 8802
rect 15334 8744 17498 8800
rect 17554 8744 17559 8800
rect 15334 8742 17559 8744
rect 9397 8739 9463 8742
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 5996 8606 14842 8666
rect 3325 8603 3391 8606
rect 4705 8603 4771 8606
rect 0 8530 480 8560
rect 1853 8530 1919 8533
rect 3141 8532 3207 8533
rect 3141 8530 3188 8532
rect 0 8470 1778 8530
rect 0 8440 480 8470
rect 1718 8394 1778 8470
rect 1853 8528 3188 8530
rect 1853 8472 1858 8528
rect 1914 8472 3146 8528
rect 1853 8470 3188 8472
rect 1853 8467 1919 8470
rect 3141 8468 3188 8470
rect 3252 8468 3258 8532
rect 3325 8530 3391 8533
rect 4470 8530 4476 8532
rect 3325 8528 4476 8530
rect 3325 8472 3330 8528
rect 3386 8472 4476 8528
rect 3325 8470 4476 8472
rect 3141 8467 3207 8468
rect 3325 8467 3391 8470
rect 4470 8468 4476 8470
rect 4540 8468 4546 8532
rect 5073 8530 5139 8533
rect 5206 8530 5212 8532
rect 5073 8528 5212 8530
rect 5073 8472 5078 8528
rect 5134 8472 5212 8528
rect 5073 8470 5212 8472
rect 5073 8467 5139 8470
rect 5206 8468 5212 8470
rect 5276 8468 5282 8532
rect 5625 8530 5691 8533
rect 11053 8530 11119 8533
rect 12065 8532 12131 8533
rect 5625 8528 11119 8530
rect 5625 8472 5630 8528
rect 5686 8472 11058 8528
rect 11114 8472 11119 8528
rect 5625 8470 11119 8472
rect 5625 8467 5691 8470
rect 11053 8467 11119 8470
rect 12014 8468 12020 8532
rect 12084 8530 12131 8532
rect 12893 8530 12959 8533
rect 13721 8530 13787 8533
rect 12084 8528 12176 8530
rect 12126 8472 12176 8528
rect 12084 8470 12176 8472
rect 12893 8528 13787 8530
rect 12893 8472 12898 8528
rect 12954 8472 13726 8528
rect 13782 8472 13787 8528
rect 12893 8470 13787 8472
rect 14782 8530 14842 8606
rect 15334 8530 15394 8742
rect 17493 8739 17559 8742
rect 18781 8802 18847 8805
rect 19190 8802 19196 8804
rect 18781 8800 19196 8802
rect 18781 8744 18786 8800
rect 18842 8744 19196 8800
rect 18781 8742 19196 8744
rect 18781 8739 18847 8742
rect 19190 8740 19196 8742
rect 19260 8740 19266 8804
rect 20161 8802 20227 8805
rect 23657 8802 23723 8805
rect 23841 8804 23907 8805
rect 20161 8800 23723 8802
rect 20161 8744 20166 8800
rect 20222 8744 23662 8800
rect 23718 8744 23723 8800
rect 20161 8742 23723 8744
rect 20161 8739 20227 8742
rect 23657 8739 23723 8742
rect 23790 8740 23796 8804
rect 23860 8802 23907 8804
rect 23860 8800 23952 8802
rect 23902 8744 23952 8800
rect 23860 8742 23952 8744
rect 23860 8740 23907 8742
rect 23841 8739 23907 8740
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 15745 8666 15811 8669
rect 17309 8666 17375 8669
rect 15745 8664 17375 8666
rect 15745 8608 15750 8664
rect 15806 8608 17314 8664
rect 17370 8608 17375 8664
rect 15745 8606 17375 8608
rect 15745 8603 15811 8606
rect 17309 8603 17375 8606
rect 18321 8666 18387 8669
rect 20989 8666 21055 8669
rect 18321 8664 21055 8666
rect 18321 8608 18326 8664
rect 18382 8608 20994 8664
rect 21050 8608 21055 8664
rect 18321 8606 21055 8608
rect 18321 8603 18387 8606
rect 20989 8603 21055 8606
rect 21173 8666 21239 8669
rect 23933 8666 23999 8669
rect 21173 8664 23999 8666
rect 21173 8608 21178 8664
rect 21234 8608 23938 8664
rect 23994 8608 23999 8664
rect 21173 8606 23999 8608
rect 21173 8603 21239 8606
rect 23933 8603 23999 8606
rect 14782 8470 15394 8530
rect 16205 8530 16271 8533
rect 22185 8530 22251 8533
rect 16205 8528 22251 8530
rect 16205 8472 16210 8528
rect 16266 8472 22190 8528
rect 22246 8472 22251 8528
rect 16205 8470 22251 8472
rect 12084 8468 12131 8470
rect 12065 8467 12131 8468
rect 12893 8467 12959 8470
rect 13721 8467 13787 8470
rect 16205 8467 16271 8470
rect 22185 8467 22251 8470
rect 22737 8530 22803 8533
rect 27520 8530 28000 8560
rect 22737 8528 28000 8530
rect 22737 8472 22742 8528
rect 22798 8472 28000 8528
rect 22737 8470 28000 8472
rect 22737 8467 22803 8470
rect 3328 8394 3388 8467
rect 27520 8440 28000 8470
rect 1718 8334 3388 8394
rect 9673 8394 9739 8397
rect 17309 8394 17375 8397
rect 21817 8394 21883 8397
rect 9673 8392 16498 8394
rect 9673 8336 9678 8392
rect 9734 8336 16498 8392
rect 9673 8334 16498 8336
rect 9673 8331 9739 8334
rect 5533 8258 5599 8261
rect 2638 8256 5599 8258
rect 2638 8200 5538 8256
rect 5594 8200 5599 8256
rect 2638 8198 5599 8200
rect 2497 8122 2563 8125
rect 2638 8122 2698 8198
rect 5533 8195 5599 8198
rect 10685 8258 10751 8261
rect 13813 8258 13879 8261
rect 10685 8256 13879 8258
rect 10685 8200 10690 8256
rect 10746 8200 13818 8256
rect 13874 8200 13879 8256
rect 10685 8198 13879 8200
rect 10685 8195 10751 8198
rect 13813 8195 13879 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 2497 8120 2698 8122
rect 2497 8064 2502 8120
rect 2558 8064 2698 8120
rect 2497 8062 2698 8064
rect 2497 8059 2563 8062
rect 6913 7986 6979 7989
rect 2776 7984 6979 7986
rect 2776 7952 6918 7984
rect 2684 7928 6918 7952
rect 6974 7928 6979 7984
rect 2684 7926 6979 7928
rect 16438 7986 16498 8334
rect 17309 8392 21883 8394
rect 17309 8336 17314 8392
rect 17370 8336 21822 8392
rect 21878 8336 21883 8392
rect 17309 8334 21883 8336
rect 17309 8331 17375 8334
rect 21817 8331 21883 8334
rect 21950 8332 21956 8396
rect 22020 8394 22026 8396
rect 22921 8394 22987 8397
rect 22020 8392 22987 8394
rect 22020 8336 22926 8392
rect 22982 8336 22987 8392
rect 22020 8334 22987 8336
rect 22020 8332 22026 8334
rect 22921 8331 22987 8334
rect 23473 8394 23539 8397
rect 24761 8394 24827 8397
rect 23473 8392 24827 8394
rect 23473 8336 23478 8392
rect 23534 8336 24766 8392
rect 24822 8336 24827 8392
rect 23473 8334 24827 8336
rect 23473 8331 23539 8334
rect 24761 8331 24827 8334
rect 21173 8258 21239 8261
rect 23657 8258 23723 8261
rect 21173 8256 23723 8258
rect 21173 8200 21178 8256
rect 21234 8200 23662 8256
rect 23718 8200 23723 8256
rect 21173 8198 23723 8200
rect 21173 8195 21239 8198
rect 23657 8195 23723 8198
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 20253 8122 20319 8125
rect 24853 8122 24919 8125
rect 20253 8120 24919 8122
rect 20253 8064 20258 8120
rect 20314 8064 24858 8120
rect 24914 8064 24919 8120
rect 20253 8062 24919 8064
rect 20253 8059 20319 8062
rect 24853 8059 24919 8062
rect 25037 8122 25103 8125
rect 25630 8122 25636 8124
rect 25037 8120 25636 8122
rect 25037 8064 25042 8120
rect 25098 8064 25636 8120
rect 25037 8062 25636 8064
rect 25037 8059 25103 8062
rect 25630 8060 25636 8062
rect 25700 8060 25706 8124
rect 20897 7986 20963 7989
rect 22829 7986 22895 7989
rect 16438 7984 20963 7986
rect 16438 7928 20902 7984
rect 20958 7928 20963 7984
rect 16438 7926 20963 7928
rect 2684 7892 2836 7926
rect 6913 7923 6979 7926
rect 20897 7923 20963 7926
rect 21038 7984 22895 7986
rect 21038 7928 22834 7984
rect 22890 7928 22895 7984
rect 21038 7926 22895 7928
rect 0 7850 480 7880
rect 2684 7850 2744 7892
rect 2957 7852 3023 7853
rect 2957 7850 3004 7852
rect 0 7790 2744 7850
rect 2912 7848 3004 7850
rect 2912 7792 2962 7848
rect 2912 7790 3004 7792
rect 0 7760 480 7790
rect 2957 7788 3004 7790
rect 3068 7788 3074 7852
rect 3693 7850 3759 7853
rect 6494 7850 6500 7852
rect 3693 7848 6500 7850
rect 3693 7792 3698 7848
rect 3754 7792 6500 7848
rect 3693 7790 6500 7792
rect 2957 7787 3023 7788
rect 3693 7787 3759 7790
rect 6494 7788 6500 7790
rect 6564 7788 6570 7852
rect 7925 7850 7991 7853
rect 19885 7850 19951 7853
rect 7925 7848 19951 7850
rect 7925 7792 7930 7848
rect 7986 7792 19890 7848
rect 19946 7792 19951 7848
rect 7925 7790 19951 7792
rect 7925 7787 7991 7790
rect 19885 7787 19951 7790
rect 20161 7850 20227 7853
rect 21038 7850 21098 7926
rect 22829 7923 22895 7926
rect 23657 7986 23723 7989
rect 23657 7984 26250 7986
rect 23657 7928 23662 7984
rect 23718 7928 26250 7984
rect 23657 7926 26250 7928
rect 23657 7923 23723 7926
rect 20161 7848 21098 7850
rect 20161 7792 20166 7848
rect 20222 7792 21098 7848
rect 20161 7790 21098 7792
rect 20161 7787 20227 7790
rect 24894 7788 24900 7852
rect 24964 7850 24970 7852
rect 26049 7850 26115 7853
rect 24964 7848 26115 7850
rect 24964 7792 26054 7848
rect 26110 7792 26115 7848
rect 24964 7790 26115 7792
rect 26190 7850 26250 7926
rect 27520 7850 28000 7880
rect 26190 7790 28000 7850
rect 24964 7788 24970 7790
rect 26049 7787 26115 7790
rect 27520 7760 28000 7790
rect 2405 7714 2471 7717
rect 4429 7714 4495 7717
rect 2405 7712 4495 7714
rect 2405 7656 2410 7712
rect 2466 7656 4434 7712
rect 4490 7656 4495 7712
rect 2405 7654 4495 7656
rect 2405 7651 2471 7654
rect 4429 7651 4495 7654
rect 19425 7714 19491 7717
rect 23289 7714 23355 7717
rect 19425 7712 23355 7714
rect 19425 7656 19430 7712
rect 19486 7656 23294 7712
rect 23350 7656 23355 7712
rect 19425 7654 23355 7656
rect 19425 7651 19491 7654
rect 23289 7651 23355 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 3417 7578 3483 7581
rect 5349 7578 5415 7581
rect 1350 7576 3483 7578
rect 1350 7520 3422 7576
rect 3478 7520 3483 7576
rect 1350 7518 3483 7520
rect 0 7306 480 7336
rect 1350 7306 1410 7518
rect 3417 7515 3483 7518
rect 3558 7576 5415 7578
rect 3558 7520 5354 7576
rect 5410 7520 5415 7576
rect 3558 7518 5415 7520
rect 2037 7442 2103 7445
rect 3558 7442 3618 7518
rect 5349 7515 5415 7518
rect 7414 7516 7420 7580
rect 7484 7578 7490 7580
rect 7557 7578 7623 7581
rect 7484 7576 7623 7578
rect 7484 7520 7562 7576
rect 7618 7520 7623 7576
rect 7484 7518 7623 7520
rect 7484 7516 7490 7518
rect 7557 7515 7623 7518
rect 8569 7578 8635 7581
rect 12157 7578 12223 7581
rect 13997 7578 14063 7581
rect 21357 7578 21423 7581
rect 8569 7576 11162 7578
rect 8569 7520 8574 7576
rect 8630 7520 11162 7576
rect 8569 7518 11162 7520
rect 8569 7515 8635 7518
rect 5165 7444 5231 7445
rect 5165 7442 5212 7444
rect 2037 7440 3618 7442
rect 2037 7384 2042 7440
rect 2098 7384 3618 7440
rect 2037 7382 3618 7384
rect 5120 7440 5212 7442
rect 5120 7384 5170 7440
rect 5120 7382 5212 7384
rect 2037 7379 2103 7382
rect 5165 7380 5212 7382
rect 5276 7380 5282 7444
rect 7097 7442 7163 7445
rect 11102 7442 11162 7518
rect 12157 7576 14063 7578
rect 12157 7520 12162 7576
rect 12218 7520 14002 7576
rect 14058 7520 14063 7576
rect 12157 7518 14063 7520
rect 12157 7515 12223 7518
rect 13997 7515 14063 7518
rect 19198 7576 21423 7578
rect 19198 7520 21362 7576
rect 21418 7520 21423 7576
rect 19198 7518 21423 7520
rect 12433 7442 12499 7445
rect 19198 7442 19258 7518
rect 21357 7515 21423 7518
rect 7097 7440 10978 7442
rect 7097 7384 7102 7440
rect 7158 7384 10978 7440
rect 7097 7382 10978 7384
rect 11102 7440 12499 7442
rect 11102 7384 12438 7440
rect 12494 7384 12499 7440
rect 11102 7382 12499 7384
rect 5165 7379 5231 7380
rect 7097 7379 7163 7382
rect 7189 7306 7255 7309
rect 7373 7306 7439 7309
rect 0 7246 1410 7306
rect 5030 7304 7439 7306
rect 5030 7248 7194 7304
rect 7250 7248 7378 7304
rect 7434 7248 7439 7304
rect 5030 7246 7439 7248
rect 0 7216 480 7246
rect 5030 7170 5090 7246
rect 7189 7243 7255 7246
rect 7373 7243 7439 7246
rect 9213 7306 9279 7309
rect 10918 7306 10978 7382
rect 12433 7379 12499 7382
rect 13494 7382 19258 7442
rect 13494 7306 13554 7382
rect 19374 7380 19380 7444
rect 19444 7442 19450 7444
rect 19977 7442 20043 7445
rect 19444 7440 20043 7442
rect 19444 7384 19982 7440
rect 20038 7384 20043 7440
rect 19444 7382 20043 7384
rect 19444 7380 19450 7382
rect 19977 7379 20043 7382
rect 21541 7442 21607 7445
rect 23473 7442 23539 7445
rect 21541 7440 23539 7442
rect 21541 7384 21546 7440
rect 21602 7384 23478 7440
rect 23534 7384 23539 7440
rect 21541 7382 23539 7384
rect 21541 7379 21607 7382
rect 23473 7379 23539 7382
rect 9213 7304 10840 7306
rect 9213 7248 9218 7304
rect 9274 7248 10840 7304
rect 9213 7246 10840 7248
rect 10918 7246 13554 7306
rect 13629 7306 13695 7309
rect 14549 7306 14615 7309
rect 20713 7306 20779 7309
rect 13629 7304 20779 7306
rect 13629 7248 13634 7304
rect 13690 7248 14554 7304
rect 14610 7248 20718 7304
rect 20774 7248 20779 7304
rect 13629 7246 20779 7248
rect 9213 7243 9279 7246
rect 3604 7110 5090 7170
rect 5349 7170 5415 7173
rect 5349 7168 6746 7170
rect 5349 7112 5354 7168
rect 5410 7112 6746 7168
rect 5349 7110 6746 7112
rect 1577 7034 1643 7037
rect 3604 7034 3664 7110
rect 5349 7107 5415 7110
rect 1577 7032 3664 7034
rect 1577 6976 1582 7032
rect 1638 6976 3664 7032
rect 1577 6974 3664 6976
rect 1577 6971 1643 6974
rect 3734 6972 3740 7036
rect 3804 7034 3810 7036
rect 4061 7034 4127 7037
rect 6686 7034 6746 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 7925 7034 7991 7037
rect 8845 7034 8911 7037
rect 3804 7032 4127 7034
rect 3804 6976 4066 7032
rect 4122 6976 4127 7032
rect 3804 6974 4127 6976
rect 3804 6972 3810 6974
rect 4061 6971 4127 6974
rect 5030 6974 6562 7034
rect 6686 7032 8911 7034
rect 6686 6976 7930 7032
rect 7986 6976 8850 7032
rect 8906 6976 8911 7032
rect 6686 6974 8911 6976
rect 10780 7034 10840 7246
rect 13629 7243 13695 7246
rect 14549 7243 14615 7246
rect 20713 7243 20779 7246
rect 21817 7306 21883 7309
rect 27520 7306 28000 7336
rect 21817 7304 28000 7306
rect 21817 7248 21822 7304
rect 21878 7248 28000 7304
rect 21817 7246 28000 7248
rect 21817 7243 21883 7246
rect 27520 7216 28000 7246
rect 10961 7170 11027 7173
rect 13169 7170 13235 7173
rect 10961 7168 13235 7170
rect 10961 7112 10966 7168
rect 11022 7112 13174 7168
rect 13230 7112 13235 7168
rect 10961 7110 13235 7112
rect 10961 7107 11027 7110
rect 13169 7107 13235 7110
rect 14181 7170 14247 7173
rect 19333 7170 19399 7173
rect 14181 7168 19399 7170
rect 14181 7112 14186 7168
rect 14242 7112 19338 7168
rect 19394 7112 19399 7168
rect 14181 7110 19399 7112
rect 14181 7107 14247 7110
rect 19333 7107 19399 7110
rect 21633 7170 21699 7173
rect 23473 7170 23539 7173
rect 21633 7168 23539 7170
rect 21633 7112 21638 7168
rect 21694 7112 23478 7168
rect 23534 7112 23539 7168
rect 21633 7110 23539 7112
rect 21633 7107 21699 7110
rect 23473 7107 23539 7110
rect 26182 7108 26188 7172
rect 26252 7170 26258 7172
rect 26417 7170 26483 7173
rect 26252 7168 26483 7170
rect 26252 7112 26422 7168
rect 26478 7112 26483 7168
rect 26252 7110 26483 7112
rect 26252 7108 26258 7110
rect 26417 7107 26483 7110
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 14273 7034 14339 7037
rect 10780 7032 14339 7034
rect 10780 6976 14278 7032
rect 14334 6976 14339 7032
rect 10780 6974 14339 6976
rect 3509 6898 3575 6901
rect 4838 6898 4844 6900
rect 3509 6896 4844 6898
rect 3509 6840 3514 6896
rect 3570 6840 4844 6896
rect 3509 6838 4844 6840
rect 3509 6835 3575 6838
rect 4838 6836 4844 6838
rect 4908 6836 4914 6900
rect 0 6762 480 6792
rect 2405 6762 2471 6765
rect 5030 6762 5090 6974
rect 5257 6898 5323 6901
rect 5257 6896 6424 6898
rect 5257 6840 5262 6896
rect 5318 6840 6424 6896
rect 5257 6838 6424 6840
rect 5257 6835 5323 6838
rect 6085 6764 6151 6765
rect 6085 6762 6132 6764
rect 0 6702 1410 6762
rect 0 6672 480 6702
rect 1350 6626 1410 6702
rect 2405 6760 5090 6762
rect 2405 6704 2410 6760
rect 2466 6704 5090 6760
rect 2405 6702 5090 6704
rect 6040 6760 6132 6762
rect 6040 6704 6090 6760
rect 6040 6702 6132 6704
rect 2405 6699 2471 6702
rect 6085 6700 6132 6702
rect 6196 6700 6202 6764
rect 6085 6699 6151 6700
rect 4981 6626 5047 6629
rect 1350 6624 5047 6626
rect 1350 6568 4986 6624
rect 5042 6568 5047 6624
rect 1350 6566 5047 6568
rect 6364 6626 6424 6838
rect 6502 6762 6562 6974
rect 7925 6971 7991 6974
rect 8845 6971 8911 6974
rect 14273 6971 14339 6974
rect 14733 7034 14799 7037
rect 16849 7034 16915 7037
rect 14733 7032 16915 7034
rect 14733 6976 14738 7032
rect 14794 6976 16854 7032
rect 16910 6976 16915 7032
rect 14733 6974 16915 6976
rect 14733 6971 14799 6974
rect 16849 6971 16915 6974
rect 18413 7034 18479 7037
rect 19149 7034 19215 7037
rect 19425 7034 19491 7037
rect 18413 7032 19491 7034
rect 18413 6976 18418 7032
rect 18474 6976 19154 7032
rect 19210 6976 19430 7032
rect 19486 6976 19491 7032
rect 18413 6974 19491 6976
rect 18413 6971 18479 6974
rect 19149 6971 19215 6974
rect 19425 6971 19491 6974
rect 20897 7034 20963 7037
rect 22921 7034 22987 7037
rect 20897 7032 22987 7034
rect 20897 6976 20902 7032
rect 20958 6976 22926 7032
rect 22982 6976 22987 7032
rect 20897 6974 22987 6976
rect 20897 6971 20963 6974
rect 22921 6971 22987 6974
rect 24894 6972 24900 7036
rect 24964 7034 24970 7036
rect 25681 7034 25747 7037
rect 24964 7032 25747 7034
rect 24964 6976 25686 7032
rect 25742 6976 25747 7032
rect 24964 6974 25747 6976
rect 24964 6972 24970 6974
rect 25681 6971 25747 6974
rect 6821 6898 6887 6901
rect 17953 6898 18019 6901
rect 6821 6896 18019 6898
rect 6821 6840 6826 6896
rect 6882 6840 17958 6896
rect 18014 6840 18019 6896
rect 6821 6838 18019 6840
rect 6821 6835 6887 6838
rect 17953 6835 18019 6838
rect 18086 6836 18092 6900
rect 18156 6898 18162 6900
rect 20805 6898 20871 6901
rect 18156 6896 20871 6898
rect 18156 6840 20810 6896
rect 20866 6840 20871 6896
rect 18156 6838 20871 6840
rect 18156 6836 18162 6838
rect 20805 6835 20871 6838
rect 21449 6898 21515 6901
rect 21766 6898 21772 6900
rect 21449 6896 21772 6898
rect 21449 6840 21454 6896
rect 21510 6840 21772 6896
rect 21449 6838 21772 6840
rect 21449 6835 21515 6838
rect 21766 6836 21772 6838
rect 21836 6836 21842 6900
rect 22645 6898 22711 6901
rect 25037 6898 25103 6901
rect 22645 6896 25103 6898
rect 22645 6840 22650 6896
rect 22706 6840 25042 6896
rect 25098 6840 25103 6896
rect 22645 6838 25103 6840
rect 22645 6835 22711 6838
rect 25037 6835 25103 6838
rect 10409 6762 10475 6765
rect 6502 6760 10475 6762
rect 6502 6704 10414 6760
rect 10470 6704 10475 6760
rect 6502 6702 10475 6704
rect 10409 6699 10475 6702
rect 10593 6762 10659 6765
rect 13353 6762 13419 6765
rect 20897 6762 20963 6765
rect 10593 6760 13419 6762
rect 10593 6704 10598 6760
rect 10654 6704 13358 6760
rect 13414 6704 13419 6760
rect 10593 6702 13419 6704
rect 10593 6699 10659 6702
rect 13353 6699 13419 6702
rect 14782 6760 20963 6762
rect 14782 6704 20902 6760
rect 20958 6704 20963 6760
rect 14782 6702 20963 6704
rect 14782 6626 14842 6702
rect 20897 6699 20963 6702
rect 21173 6762 21239 6765
rect 24025 6762 24091 6765
rect 27520 6762 28000 6792
rect 21173 6760 24091 6762
rect 21173 6704 21178 6760
rect 21234 6704 24030 6760
rect 24086 6704 24091 6760
rect 21173 6702 24091 6704
rect 21173 6699 21239 6702
rect 24025 6699 24091 6702
rect 24718 6702 28000 6762
rect 6364 6566 14842 6626
rect 16757 6626 16823 6629
rect 20529 6626 20595 6629
rect 22277 6626 22343 6629
rect 16757 6624 22343 6626
rect 16757 6568 16762 6624
rect 16818 6568 20534 6624
rect 20590 6568 22282 6624
rect 22338 6568 22343 6624
rect 16757 6566 22343 6568
rect 4981 6563 5047 6566
rect 16757 6563 16823 6566
rect 20529 6563 20595 6566
rect 22277 6563 22343 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 8109 6492 8175 6493
rect 8109 6490 8156 6492
rect 8064 6488 8156 6490
rect 8064 6432 8114 6488
rect 8064 6430 8156 6432
rect 8109 6428 8156 6430
rect 8220 6428 8226 6492
rect 9806 6428 9812 6492
rect 9876 6490 9882 6492
rect 9949 6490 10015 6493
rect 9876 6488 10015 6490
rect 9876 6432 9954 6488
rect 10010 6432 10015 6488
rect 9876 6430 10015 6432
rect 9876 6428 9882 6430
rect 8109 6427 8175 6428
rect 9949 6427 10015 6430
rect 10501 6490 10567 6493
rect 10726 6490 10732 6492
rect 10501 6488 10732 6490
rect 10501 6432 10506 6488
rect 10562 6432 10732 6488
rect 10501 6430 10732 6432
rect 10501 6427 10567 6430
rect 10726 6428 10732 6430
rect 10796 6428 10802 6492
rect 12198 6428 12204 6492
rect 12268 6490 12274 6492
rect 12525 6490 12591 6493
rect 14733 6490 14799 6493
rect 17902 6490 17908 6492
rect 12268 6488 12591 6490
rect 12268 6432 12530 6488
rect 12586 6432 12591 6488
rect 12268 6430 12591 6432
rect 12268 6428 12274 6430
rect 12525 6427 12591 6430
rect 13862 6488 14799 6490
rect 13862 6432 14738 6488
rect 14794 6432 14799 6488
rect 13862 6430 14799 6432
rect 7189 6354 7255 6357
rect 13862 6354 13922 6430
rect 14733 6427 14799 6430
rect 15334 6430 17908 6490
rect 7189 6352 13922 6354
rect 7189 6296 7194 6352
rect 7250 6296 13922 6352
rect 7189 6294 13922 6296
rect 14089 6354 14155 6357
rect 15334 6354 15394 6430
rect 17902 6428 17908 6430
rect 17972 6428 17978 6492
rect 18045 6490 18111 6493
rect 21173 6490 21239 6493
rect 18045 6488 21239 6490
rect 18045 6432 18050 6488
rect 18106 6432 21178 6488
rect 21234 6432 21239 6488
rect 18045 6430 21239 6432
rect 18045 6427 18111 6430
rect 21173 6427 21239 6430
rect 14089 6352 15394 6354
rect 14089 6296 14094 6352
rect 14150 6296 15394 6352
rect 14089 6294 15394 6296
rect 16573 6354 16639 6357
rect 18229 6354 18295 6357
rect 16573 6352 18295 6354
rect 16573 6296 16578 6352
rect 16634 6296 18234 6352
rect 18290 6296 18295 6352
rect 16573 6294 18295 6296
rect 7189 6291 7255 6294
rect 14089 6291 14155 6294
rect 16573 6291 16639 6294
rect 18229 6291 18295 6294
rect 20846 6292 20852 6356
rect 20916 6354 20922 6356
rect 21541 6354 21607 6357
rect 21766 6354 21772 6356
rect 20916 6352 21772 6354
rect 20916 6296 21546 6352
rect 21602 6296 21772 6352
rect 20916 6294 21772 6296
rect 20916 6292 20922 6294
rect 21541 6291 21607 6294
rect 21766 6292 21772 6294
rect 21836 6292 21842 6356
rect 23422 6292 23428 6356
rect 23492 6354 23498 6356
rect 24718 6354 24778 6702
rect 27520 6672 28000 6702
rect 23492 6294 24778 6354
rect 23492 6292 23498 6294
rect 1853 6218 1919 6221
rect 2589 6218 2655 6221
rect 8753 6218 8819 6221
rect 1853 6216 8819 6218
rect 1853 6160 1858 6216
rect 1914 6160 2594 6216
rect 2650 6160 8758 6216
rect 8814 6160 8819 6216
rect 1853 6158 8819 6160
rect 1853 6155 1919 6158
rect 2589 6155 2655 6158
rect 8753 6155 8819 6158
rect 9949 6218 10015 6221
rect 17718 6218 17724 6220
rect 9949 6216 17724 6218
rect 9949 6160 9954 6216
rect 10010 6160 17724 6216
rect 9949 6158 17724 6160
rect 9949 6155 10015 6158
rect 17718 6156 17724 6158
rect 17788 6156 17794 6220
rect 19057 6218 19123 6221
rect 21265 6218 21331 6221
rect 19057 6216 21331 6218
rect 19057 6160 19062 6216
rect 19118 6160 21270 6216
rect 21326 6160 21331 6216
rect 19057 6158 21331 6160
rect 19057 6155 19123 6158
rect 21265 6155 21331 6158
rect 21725 6218 21791 6221
rect 24577 6218 24643 6221
rect 21725 6216 24643 6218
rect 21725 6160 21730 6216
rect 21786 6160 24582 6216
rect 24638 6160 24643 6216
rect 21725 6158 24643 6160
rect 21725 6155 21791 6158
rect 24577 6155 24643 6158
rect 0 6082 480 6112
rect 2681 6082 2747 6085
rect 0 6080 2747 6082
rect 0 6024 2686 6080
rect 2742 6024 2747 6080
rect 0 6022 2747 6024
rect 0 5992 480 6022
rect 2681 6019 2747 6022
rect 5349 6082 5415 6085
rect 7414 6082 7420 6084
rect 5349 6080 7420 6082
rect 5349 6024 5354 6080
rect 5410 6024 7420 6080
rect 5349 6022 7420 6024
rect 5349 6019 5415 6022
rect 7414 6020 7420 6022
rect 7484 6020 7490 6084
rect 13302 6020 13308 6084
rect 13372 6082 13378 6084
rect 15469 6082 15535 6085
rect 13372 6080 15535 6082
rect 13372 6024 15474 6080
rect 15530 6024 15535 6080
rect 13372 6022 15535 6024
rect 13372 6020 13378 6022
rect 15469 6019 15535 6022
rect 20805 6082 20871 6085
rect 22001 6082 22067 6085
rect 20805 6080 22067 6082
rect 20805 6024 20810 6080
rect 20866 6024 22006 6080
rect 22062 6024 22067 6080
rect 20805 6022 22067 6024
rect 20805 6019 20871 6022
rect 22001 6019 22067 6022
rect 23933 6082 23999 6085
rect 27520 6082 28000 6112
rect 23933 6080 28000 6082
rect 23933 6024 23938 6080
rect 23994 6024 28000 6080
rect 23933 6022 28000 6024
rect 23933 6019 23999 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 27520 5992 28000 6022
rect 19610 5951 19930 5952
rect 3417 5946 3483 5949
rect 8845 5946 8911 5949
rect 15285 5946 15351 5949
rect 18413 5946 18479 5949
rect 3417 5944 8911 5946
rect 3417 5888 3422 5944
rect 3478 5888 8850 5944
rect 8906 5888 8911 5944
rect 3417 5886 8911 5888
rect 3417 5883 3483 5886
rect 8845 5883 8911 5886
rect 10688 5886 15210 5946
rect 5165 5810 5231 5813
rect 6177 5810 6243 5813
rect 5165 5808 6243 5810
rect 5165 5752 5170 5808
rect 5226 5752 6182 5808
rect 6238 5752 6243 5808
rect 5165 5750 6243 5752
rect 5165 5747 5231 5750
rect 6177 5747 6243 5750
rect 8293 5810 8359 5813
rect 10688 5810 10748 5886
rect 8293 5808 10748 5810
rect 8293 5752 8298 5808
rect 8354 5752 10748 5808
rect 8293 5750 10748 5752
rect 11881 5810 11947 5813
rect 13721 5810 13787 5813
rect 11881 5808 13787 5810
rect 11881 5752 11886 5808
rect 11942 5752 13726 5808
rect 13782 5752 13787 5808
rect 11881 5750 13787 5752
rect 15150 5810 15210 5886
rect 15285 5944 18479 5946
rect 15285 5888 15290 5944
rect 15346 5888 18418 5944
rect 18474 5888 18479 5944
rect 15285 5886 18479 5888
rect 15285 5883 15351 5886
rect 18413 5883 18479 5886
rect 21265 5946 21331 5949
rect 26233 5946 26299 5949
rect 21265 5944 26299 5946
rect 21265 5888 21270 5944
rect 21326 5888 26238 5944
rect 26294 5888 26299 5944
rect 21265 5886 26299 5888
rect 21265 5883 21331 5886
rect 26233 5883 26299 5886
rect 20253 5810 20319 5813
rect 15150 5808 20319 5810
rect 15150 5752 20258 5808
rect 20314 5752 20319 5808
rect 15150 5750 20319 5752
rect 8293 5747 8359 5750
rect 11881 5747 11947 5750
rect 13721 5747 13787 5750
rect 20253 5747 20319 5750
rect 21357 5810 21423 5813
rect 26233 5810 26299 5813
rect 21357 5808 26299 5810
rect 21357 5752 21362 5808
rect 21418 5752 26238 5808
rect 26294 5752 26299 5808
rect 21357 5750 26299 5752
rect 21357 5747 21423 5750
rect 26233 5747 26299 5750
rect 12801 5674 12867 5677
rect 4846 5672 12867 5674
rect 4846 5616 12806 5672
rect 12862 5616 12867 5672
rect 4846 5614 12867 5616
rect 0 5538 480 5568
rect 4846 5538 4906 5614
rect 12801 5611 12867 5614
rect 12985 5674 13051 5677
rect 13905 5674 13971 5677
rect 18229 5674 18295 5677
rect 21817 5674 21883 5677
rect 12985 5672 21883 5674
rect 12985 5616 12990 5672
rect 13046 5616 13910 5672
rect 13966 5616 18234 5672
rect 18290 5616 21822 5672
rect 21878 5616 21883 5672
rect 12985 5614 21883 5616
rect 12985 5611 13051 5614
rect 13905 5611 13971 5614
rect 18229 5611 18295 5614
rect 21817 5611 21883 5614
rect 23289 5674 23355 5677
rect 23289 5672 24732 5674
rect 23289 5616 23294 5672
rect 23350 5616 24732 5672
rect 23289 5614 24732 5616
rect 23289 5611 23355 5614
rect 0 5478 4906 5538
rect 7189 5540 7255 5541
rect 7189 5536 7236 5540
rect 7300 5538 7306 5540
rect 7465 5538 7531 5541
rect 10317 5538 10383 5541
rect 7189 5480 7194 5536
rect 0 5448 480 5478
rect 7189 5476 7236 5480
rect 7300 5478 7346 5538
rect 7465 5536 10383 5538
rect 7465 5480 7470 5536
rect 7526 5480 10322 5536
rect 10378 5480 10383 5536
rect 7465 5478 10383 5480
rect 7300 5476 7306 5478
rect 7189 5475 7255 5476
rect 7465 5475 7531 5478
rect 10317 5475 10383 5478
rect 10501 5538 10567 5541
rect 13261 5538 13327 5541
rect 10501 5536 13327 5538
rect 10501 5480 10506 5536
rect 10562 5480 13266 5536
rect 13322 5480 13327 5536
rect 10501 5478 13327 5480
rect 24672 5538 24732 5614
rect 27520 5538 28000 5568
rect 24672 5478 28000 5538
rect 10501 5475 10567 5478
rect 13261 5475 13327 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 27520 5448 28000 5478
rect 24277 5407 24597 5408
rect 9622 5340 9628 5404
rect 9692 5402 9698 5404
rect 9692 5342 11714 5402
rect 9692 5340 9698 5342
rect 2313 5266 2379 5269
rect 3049 5266 3115 5269
rect 5717 5266 5783 5269
rect 2313 5264 5783 5266
rect 2313 5208 2318 5264
rect 2374 5208 3054 5264
rect 3110 5208 5722 5264
rect 5778 5208 5783 5264
rect 2313 5206 5783 5208
rect 2313 5203 2379 5206
rect 3049 5203 3115 5206
rect 5717 5203 5783 5206
rect 8017 5266 8083 5269
rect 11513 5266 11579 5269
rect 8017 5264 11579 5266
rect 8017 5208 8022 5264
rect 8078 5208 11518 5264
rect 11574 5208 11579 5264
rect 8017 5206 11579 5208
rect 11654 5266 11714 5342
rect 17718 5340 17724 5404
rect 17788 5402 17794 5404
rect 20989 5402 21055 5405
rect 17788 5400 21055 5402
rect 17788 5344 20994 5400
rect 21050 5344 21055 5400
rect 17788 5342 21055 5344
rect 17788 5340 17794 5342
rect 20989 5339 21055 5342
rect 22093 5402 22159 5405
rect 23657 5402 23723 5405
rect 24025 5404 24091 5405
rect 22093 5400 23723 5402
rect 22093 5344 22098 5400
rect 22154 5344 23662 5400
rect 23718 5344 23723 5400
rect 22093 5342 23723 5344
rect 22093 5339 22159 5342
rect 23657 5339 23723 5342
rect 23974 5340 23980 5404
rect 24044 5402 24091 5404
rect 24044 5400 24136 5402
rect 24086 5344 24136 5400
rect 24044 5342 24136 5344
rect 24044 5340 24091 5342
rect 24025 5339 24091 5340
rect 23013 5266 23079 5269
rect 11654 5264 23079 5266
rect 11654 5208 23018 5264
rect 23074 5208 23079 5264
rect 11654 5206 23079 5208
rect 8017 5203 8083 5206
rect 11513 5203 11579 5206
rect 23013 5203 23079 5206
rect 9990 5068 9996 5132
rect 10060 5130 10066 5132
rect 10869 5130 10935 5133
rect 10060 5128 10935 5130
rect 10060 5072 10874 5128
rect 10930 5072 10935 5128
rect 10060 5070 10935 5072
rect 10060 5068 10066 5070
rect 10869 5067 10935 5070
rect 13077 5130 13143 5133
rect 20713 5130 20779 5133
rect 13077 5128 20779 5130
rect 13077 5072 13082 5128
rect 13138 5072 20718 5128
rect 20774 5072 20779 5128
rect 13077 5070 20779 5072
rect 13077 5067 13143 5070
rect 20713 5067 20779 5070
rect 21633 5130 21699 5133
rect 22185 5130 22251 5133
rect 21633 5128 22251 5130
rect 21633 5072 21638 5128
rect 21694 5072 22190 5128
rect 22246 5072 22251 5128
rect 21633 5070 22251 5072
rect 21633 5067 21699 5070
rect 22185 5067 22251 5070
rect 0 4994 480 5024
rect 8937 4994 9003 4997
rect 0 4992 9003 4994
rect 0 4936 8942 4992
rect 8998 4936 9003 4992
rect 0 4934 9003 4936
rect 0 4904 480 4934
rect 8937 4931 9003 4934
rect 12065 4994 12131 4997
rect 15510 4994 15516 4996
rect 12065 4992 15516 4994
rect 12065 4936 12070 4992
rect 12126 4936 15516 4992
rect 12065 4934 15516 4936
rect 12065 4931 12131 4934
rect 15510 4932 15516 4934
rect 15580 4932 15586 4996
rect 20161 4994 20227 4997
rect 24945 4994 25011 4997
rect 20161 4992 25011 4994
rect 20161 4936 20166 4992
rect 20222 4936 24950 4992
rect 25006 4936 25011 4992
rect 20161 4934 25011 4936
rect 20161 4931 20227 4934
rect 24945 4931 25011 4934
rect 25497 4994 25563 4997
rect 27520 4994 28000 5024
rect 25497 4992 28000 4994
rect 25497 4936 25502 4992
rect 25558 4936 28000 4992
rect 25497 4934 28000 4936
rect 25497 4931 25563 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 27520 4904 28000 4934
rect 19610 4863 19930 4864
rect 9489 4858 9555 4861
rect 11605 4858 11671 4861
rect 19149 4858 19215 4861
rect 9489 4856 10058 4858
rect 9489 4800 9494 4856
rect 9550 4800 10058 4856
rect 9489 4798 10058 4800
rect 9489 4795 9555 4798
rect 2773 4722 2839 4725
rect 4153 4722 4219 4725
rect 2773 4720 4219 4722
rect 2773 4664 2778 4720
rect 2834 4664 4158 4720
rect 4214 4664 4219 4720
rect 2773 4662 4219 4664
rect 2773 4659 2839 4662
rect 4153 4659 4219 4662
rect 7557 4722 7623 4725
rect 9998 4722 10058 4798
rect 11605 4856 19215 4858
rect 11605 4800 11610 4856
rect 11666 4800 19154 4856
rect 19210 4800 19215 4856
rect 11605 4798 19215 4800
rect 11605 4795 11671 4798
rect 19149 4795 19215 4798
rect 20253 4858 20319 4861
rect 25405 4858 25471 4861
rect 20253 4856 25471 4858
rect 20253 4800 20258 4856
rect 20314 4800 25410 4856
rect 25466 4800 25471 4856
rect 20253 4798 25471 4800
rect 20253 4795 20319 4798
rect 25405 4795 25471 4798
rect 15285 4722 15351 4725
rect 7557 4720 9506 4722
rect 7557 4664 7562 4720
rect 7618 4664 9506 4720
rect 7557 4662 9506 4664
rect 9998 4720 15351 4722
rect 9998 4664 15290 4720
rect 15346 4664 15351 4720
rect 9998 4662 15351 4664
rect 7557 4659 7623 4662
rect 4061 4586 4127 4589
rect 9213 4586 9279 4589
rect 4061 4584 9279 4586
rect 4061 4528 4066 4584
rect 4122 4528 9218 4584
rect 9274 4528 9279 4584
rect 4061 4526 9279 4528
rect 9446 4586 9506 4662
rect 15285 4659 15351 4662
rect 15653 4722 15719 4725
rect 17125 4722 17191 4725
rect 15653 4720 17191 4722
rect 15653 4664 15658 4720
rect 15714 4664 17130 4720
rect 17186 4664 17191 4720
rect 15653 4662 17191 4664
rect 15653 4659 15719 4662
rect 17125 4659 17191 4662
rect 21265 4722 21331 4725
rect 25037 4722 25103 4725
rect 21265 4720 25103 4722
rect 21265 4664 21270 4720
rect 21326 4664 25042 4720
rect 25098 4664 25103 4720
rect 21265 4662 25103 4664
rect 21265 4659 21331 4662
rect 25037 4659 25103 4662
rect 14089 4586 14155 4589
rect 9446 4584 14155 4586
rect 9446 4528 14094 4584
rect 14150 4528 14155 4584
rect 9446 4526 14155 4528
rect 4061 4523 4127 4526
rect 9213 4523 9279 4526
rect 14089 4523 14155 4526
rect 14549 4586 14615 4589
rect 17677 4586 17743 4589
rect 14549 4584 17743 4586
rect 14549 4528 14554 4584
rect 14610 4528 17682 4584
rect 17738 4528 17743 4584
rect 14549 4526 17743 4528
rect 14549 4523 14615 4526
rect 17677 4523 17743 4526
rect 17861 4586 17927 4589
rect 22461 4586 22527 4589
rect 17861 4584 22527 4586
rect 17861 4528 17866 4584
rect 17922 4528 22466 4584
rect 22522 4528 22527 4584
rect 17861 4526 22527 4528
rect 17861 4523 17927 4526
rect 22461 4523 22527 4526
rect 22645 4586 22711 4589
rect 22645 4584 24732 4586
rect 22645 4528 22650 4584
rect 22706 4528 24732 4584
rect 22645 4526 24732 4528
rect 22645 4523 22711 4526
rect 0 4450 480 4480
rect 1853 4450 1919 4453
rect 0 4448 1919 4450
rect 0 4392 1858 4448
rect 1914 4392 1919 4448
rect 0 4390 1919 4392
rect 0 4360 480 4390
rect 1853 4387 1919 4390
rect 8569 4450 8635 4453
rect 9765 4450 9831 4453
rect 9990 4450 9996 4452
rect 8569 4448 9996 4450
rect 8569 4392 8574 4448
rect 8630 4392 9770 4448
rect 9826 4392 9996 4448
rect 8569 4390 9996 4392
rect 8569 4387 8635 4390
rect 9765 4387 9831 4390
rect 9990 4388 9996 4390
rect 10060 4388 10066 4452
rect 10317 4450 10383 4453
rect 14273 4450 14339 4453
rect 14549 4450 14615 4453
rect 10317 4448 14615 4450
rect 10317 4392 10322 4448
rect 10378 4392 14278 4448
rect 14334 4392 14554 4448
rect 14610 4392 14615 4448
rect 10317 4390 14615 4392
rect 10317 4387 10383 4390
rect 14273 4387 14339 4390
rect 14549 4387 14615 4390
rect 19517 4450 19583 4453
rect 20110 4450 20116 4452
rect 19517 4448 20116 4450
rect 19517 4392 19522 4448
rect 19578 4392 20116 4448
rect 19517 4390 20116 4392
rect 19517 4387 19583 4390
rect 20110 4388 20116 4390
rect 20180 4388 20186 4452
rect 20662 4388 20668 4452
rect 20732 4450 20738 4452
rect 21173 4450 21239 4453
rect 20732 4448 21239 4450
rect 20732 4392 21178 4448
rect 21234 4392 21239 4448
rect 20732 4390 21239 4392
rect 20732 4388 20738 4390
rect 21173 4387 21239 4390
rect 22645 4450 22711 4453
rect 23841 4450 23907 4453
rect 22645 4448 23907 4450
rect 22645 4392 22650 4448
rect 22706 4392 23846 4448
rect 23902 4392 23907 4448
rect 22645 4390 23907 4392
rect 24672 4450 24732 4526
rect 27520 4450 28000 4480
rect 24672 4390 28000 4450
rect 22645 4387 22711 4390
rect 23841 4387 23907 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 27520 4360 28000 4390
rect 24277 4319 24597 4320
rect 9213 4314 9279 4317
rect 11053 4314 11119 4317
rect 9213 4312 11119 4314
rect 9213 4256 9218 4312
rect 9274 4256 11058 4312
rect 11114 4256 11119 4312
rect 9213 4254 11119 4256
rect 9213 4251 9279 4254
rect 11053 4251 11119 4254
rect 18505 4314 18571 4317
rect 18505 4312 24042 4314
rect 18505 4256 18510 4312
rect 18566 4256 24042 4312
rect 18505 4254 24042 4256
rect 18505 4251 18571 4254
rect 2221 4178 2287 4181
rect 6361 4178 6427 4181
rect 2221 4176 6427 4178
rect 2221 4120 2226 4176
rect 2282 4120 6366 4176
rect 6422 4120 6427 4176
rect 2221 4118 6427 4120
rect 2221 4115 2287 4118
rect 6361 4115 6427 4118
rect 9673 4178 9739 4181
rect 11094 4178 11100 4180
rect 9673 4176 11100 4178
rect 9673 4120 9678 4176
rect 9734 4120 11100 4176
rect 9673 4118 11100 4120
rect 9673 4115 9739 4118
rect 11094 4116 11100 4118
rect 11164 4116 11170 4180
rect 12065 4178 12131 4181
rect 14641 4178 14707 4181
rect 12065 4176 14707 4178
rect 12065 4120 12070 4176
rect 12126 4120 14646 4176
rect 14702 4120 14707 4176
rect 12065 4118 14707 4120
rect 12065 4115 12131 4118
rect 14641 4115 14707 4118
rect 15009 4178 15075 4181
rect 22461 4178 22527 4181
rect 15009 4176 22527 4178
rect 15009 4120 15014 4176
rect 15070 4120 22466 4176
rect 22522 4120 22527 4176
rect 15009 4118 22527 4120
rect 15009 4115 15075 4118
rect 22461 4115 22527 4118
rect 22737 4178 22803 4181
rect 23381 4178 23447 4181
rect 22737 4176 23447 4178
rect 22737 4120 22742 4176
rect 22798 4120 23386 4176
rect 23442 4120 23447 4176
rect 22737 4118 23447 4120
rect 23982 4178 24042 4254
rect 24945 4178 25011 4181
rect 23982 4176 25011 4178
rect 23982 4120 24950 4176
rect 25006 4120 25011 4176
rect 23982 4118 25011 4120
rect 22737 4115 22803 4118
rect 23381 4115 23447 4118
rect 24945 4115 25011 4118
rect 3877 4042 3943 4045
rect 11513 4042 11579 4045
rect 3877 4040 11579 4042
rect 3877 3984 3882 4040
rect 3938 3984 11518 4040
rect 11574 3984 11579 4040
rect 3877 3982 11579 3984
rect 3877 3979 3943 3982
rect 11513 3979 11579 3982
rect 12525 4042 12591 4045
rect 15745 4042 15811 4045
rect 12525 4040 15811 4042
rect 12525 3984 12530 4040
rect 12586 3984 15750 4040
rect 15806 3984 15811 4040
rect 12525 3982 15811 3984
rect 12525 3979 12591 3982
rect 15745 3979 15811 3982
rect 20713 4042 20779 4045
rect 25037 4042 25103 4045
rect 20713 4040 25103 4042
rect 20713 3984 20718 4040
rect 20774 3984 25042 4040
rect 25098 3984 25103 4040
rect 20713 3982 25103 3984
rect 20713 3979 20779 3982
rect 25037 3979 25103 3982
rect 25313 4042 25379 4045
rect 27061 4042 27127 4045
rect 25313 4040 27127 4042
rect 25313 3984 25318 4040
rect 25374 3984 27066 4040
rect 27122 3984 27127 4040
rect 25313 3982 27127 3984
rect 25313 3979 25379 3982
rect 27061 3979 27127 3982
rect 7557 3906 7623 3909
rect 8477 3906 8543 3909
rect 7557 3904 8543 3906
rect 7557 3848 7562 3904
rect 7618 3848 8482 3904
rect 8538 3848 8543 3904
rect 7557 3846 8543 3848
rect 7557 3843 7623 3846
rect 8477 3843 8543 3846
rect 11789 3906 11855 3909
rect 16757 3906 16823 3909
rect 11789 3904 16823 3906
rect 11789 3848 11794 3904
rect 11850 3848 16762 3904
rect 16818 3848 16823 3904
rect 11789 3846 16823 3848
rect 11789 3843 11855 3846
rect 16757 3843 16823 3846
rect 21030 3844 21036 3908
rect 21100 3906 21106 3908
rect 21357 3906 21423 3909
rect 21100 3904 21423 3906
rect 21100 3848 21362 3904
rect 21418 3848 21423 3904
rect 21100 3846 21423 3848
rect 21100 3844 21106 3846
rect 21357 3843 21423 3846
rect 24209 3906 24275 3909
rect 26509 3906 26575 3909
rect 24209 3904 26575 3906
rect 24209 3848 24214 3904
rect 24270 3848 26514 3904
rect 26570 3848 26575 3904
rect 24209 3846 26575 3848
rect 24209 3843 24275 3846
rect 26509 3843 26575 3846
rect 10277 3840 10597 3841
rect 0 3770 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 4153 3770 4219 3773
rect 0 3768 4219 3770
rect 0 3712 4158 3768
rect 4214 3712 4219 3768
rect 0 3710 4219 3712
rect 0 3680 480 3710
rect 4153 3707 4219 3710
rect 4521 3770 4587 3773
rect 6126 3770 6132 3772
rect 4521 3768 6132 3770
rect 4521 3712 4526 3768
rect 4582 3712 6132 3768
rect 4521 3710 6132 3712
rect 4521 3707 4587 3710
rect 6126 3708 6132 3710
rect 6196 3708 6202 3772
rect 8293 3770 8359 3773
rect 9438 3770 9444 3772
rect 8293 3768 9444 3770
rect 8293 3712 8298 3768
rect 8354 3712 9444 3768
rect 8293 3710 9444 3712
rect 8293 3707 8359 3710
rect 9438 3708 9444 3710
rect 9508 3708 9514 3772
rect 13670 3708 13676 3772
rect 13740 3770 13746 3772
rect 15377 3770 15443 3773
rect 13740 3768 15443 3770
rect 13740 3712 15382 3768
rect 15438 3712 15443 3768
rect 13740 3710 15443 3712
rect 13740 3708 13746 3710
rect 15377 3707 15443 3710
rect 16297 3770 16363 3773
rect 18045 3770 18111 3773
rect 16297 3768 18111 3770
rect 16297 3712 16302 3768
rect 16358 3712 18050 3768
rect 18106 3712 18111 3768
rect 16297 3710 18111 3712
rect 16297 3707 16363 3710
rect 18045 3707 18111 3710
rect 20621 3770 20687 3773
rect 21541 3770 21607 3773
rect 20621 3768 21607 3770
rect 20621 3712 20626 3768
rect 20682 3712 21546 3768
rect 21602 3712 21607 3768
rect 20621 3710 21607 3712
rect 20621 3707 20687 3710
rect 21541 3707 21607 3710
rect 21766 3708 21772 3772
rect 21836 3770 21842 3772
rect 25221 3770 25287 3773
rect 27520 3770 28000 3800
rect 21836 3710 24962 3770
rect 21836 3708 21842 3710
rect 5165 3634 5231 3637
rect 6453 3634 6519 3637
rect 5165 3632 6519 3634
rect 5165 3576 5170 3632
rect 5226 3576 6458 3632
rect 6514 3576 6519 3632
rect 5165 3574 6519 3576
rect 5165 3571 5231 3574
rect 6453 3571 6519 3574
rect 8017 3634 8083 3637
rect 9489 3634 9555 3637
rect 8017 3632 9555 3634
rect 8017 3576 8022 3632
rect 8078 3576 9494 3632
rect 9550 3576 9555 3632
rect 8017 3574 9555 3576
rect 8017 3571 8083 3574
rect 9489 3571 9555 3574
rect 14273 3634 14339 3637
rect 17769 3634 17835 3637
rect 23473 3634 23539 3637
rect 14273 3632 23539 3634
rect 14273 3576 14278 3632
rect 14334 3576 17774 3632
rect 17830 3576 23478 3632
rect 23534 3576 23539 3632
rect 14273 3574 23539 3576
rect 14273 3571 14339 3574
rect 17769 3571 17835 3574
rect 23473 3571 23539 3574
rect 7833 3498 7899 3501
rect 11789 3498 11855 3501
rect 14365 3500 14431 3501
rect 14365 3498 14412 3500
rect 7833 3496 11855 3498
rect 7833 3440 7838 3496
rect 7894 3440 11794 3496
rect 11850 3440 11855 3496
rect 7833 3438 11855 3440
rect 14320 3496 14412 3498
rect 14320 3440 14370 3496
rect 14320 3438 14412 3440
rect 7833 3435 7899 3438
rect 11789 3435 11855 3438
rect 14365 3436 14412 3438
rect 14476 3436 14482 3500
rect 18137 3498 18203 3501
rect 20989 3498 21055 3501
rect 18137 3496 21055 3498
rect 18137 3440 18142 3496
rect 18198 3440 20994 3496
rect 21050 3440 21055 3496
rect 18137 3438 21055 3440
rect 14365 3435 14431 3436
rect 18137 3435 18203 3438
rect 20989 3435 21055 3438
rect 8569 3362 8635 3365
rect 9581 3362 9647 3365
rect 8569 3360 9647 3362
rect 8569 3304 8574 3360
rect 8630 3304 9586 3360
rect 9642 3304 9647 3360
rect 8569 3302 9647 3304
rect 8569 3299 8635 3302
rect 9581 3299 9647 3302
rect 9765 3362 9831 3365
rect 12065 3362 12131 3365
rect 9765 3360 12131 3362
rect 9765 3304 9770 3360
rect 9826 3304 12070 3360
rect 12126 3304 12131 3360
rect 9765 3302 12131 3304
rect 9765 3299 9831 3302
rect 12065 3299 12131 3302
rect 12249 3362 12315 3365
rect 14549 3362 14615 3365
rect 19977 3362 20043 3365
rect 12249 3360 14615 3362
rect 12249 3304 12254 3360
rect 12310 3304 14554 3360
rect 14610 3304 14615 3360
rect 12249 3302 14615 3304
rect 12249 3299 12315 3302
rect 14549 3299 14615 3302
rect 15702 3360 20043 3362
rect 15702 3304 19982 3360
rect 20038 3304 20043 3360
rect 15702 3302 20043 3304
rect 5610 3296 5930 3297
rect 0 3226 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 3141 3226 3207 3229
rect 10777 3226 10843 3229
rect 14457 3228 14523 3229
rect 0 3224 3207 3226
rect 0 3168 3146 3224
rect 3202 3168 3207 3224
rect 0 3166 3207 3168
rect 0 3136 480 3166
rect 3141 3163 3207 3166
rect 6502 3224 10843 3226
rect 6502 3168 10782 3224
rect 10838 3168 10843 3224
rect 6502 3166 10843 3168
rect 657 3090 723 3093
rect 6502 3090 6562 3166
rect 10777 3163 10843 3166
rect 14406 3164 14412 3228
rect 14476 3226 14523 3228
rect 14476 3224 14568 3226
rect 14518 3168 14568 3224
rect 14476 3166 14568 3168
rect 14476 3164 14523 3166
rect 14457 3163 14523 3164
rect 657 3088 6562 3090
rect 657 3032 662 3088
rect 718 3032 6562 3088
rect 657 3030 6562 3032
rect 657 3027 723 3030
rect 6678 3028 6684 3092
rect 6748 3090 6754 3092
rect 6821 3090 6887 3093
rect 6748 3088 6887 3090
rect 6748 3032 6826 3088
rect 6882 3032 6887 3088
rect 6748 3030 6887 3032
rect 6748 3028 6754 3030
rect 6821 3027 6887 3030
rect 8937 3090 9003 3093
rect 11237 3090 11303 3093
rect 8937 3088 11303 3090
rect 8937 3032 8942 3088
rect 8998 3032 11242 3088
rect 11298 3032 11303 3088
rect 8937 3030 11303 3032
rect 8937 3027 9003 3030
rect 11237 3027 11303 3030
rect 14549 3090 14615 3093
rect 15702 3090 15762 3302
rect 19977 3299 20043 3302
rect 21265 3362 21331 3365
rect 23422 3362 23428 3364
rect 21265 3360 23428 3362
rect 21265 3304 21270 3360
rect 21326 3304 23428 3360
rect 21265 3302 23428 3304
rect 21265 3299 21331 3302
rect 23422 3300 23428 3302
rect 23492 3300 23498 3364
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 16205 3226 16271 3229
rect 18413 3226 18479 3229
rect 16205 3224 18479 3226
rect 16205 3168 16210 3224
rect 16266 3168 18418 3224
rect 18474 3168 18479 3224
rect 16205 3166 18479 3168
rect 16205 3163 16271 3166
rect 18413 3163 18479 3166
rect 18597 3226 18663 3229
rect 20989 3226 21055 3229
rect 18597 3224 21055 3226
rect 18597 3168 18602 3224
rect 18658 3168 20994 3224
rect 21050 3168 21055 3224
rect 18597 3166 21055 3168
rect 18597 3163 18663 3166
rect 20989 3163 21055 3166
rect 21173 3226 21239 3229
rect 24025 3226 24091 3229
rect 21173 3224 24091 3226
rect 21173 3168 21178 3224
rect 21234 3168 24030 3224
rect 24086 3168 24091 3224
rect 21173 3166 24091 3168
rect 24902 3226 24962 3710
rect 25221 3768 28000 3770
rect 25221 3712 25226 3768
rect 25282 3712 28000 3768
rect 25221 3710 28000 3712
rect 25221 3707 25287 3710
rect 27520 3680 28000 3710
rect 25405 3498 25471 3501
rect 27613 3498 27679 3501
rect 25405 3496 27679 3498
rect 25405 3440 25410 3496
rect 25466 3440 27618 3496
rect 27674 3440 27679 3496
rect 25405 3438 27679 3440
rect 25405 3435 25471 3438
rect 27613 3435 27679 3438
rect 27520 3226 28000 3256
rect 24902 3166 28000 3226
rect 21173 3163 21239 3166
rect 23982 3163 24091 3166
rect 14549 3088 15762 3090
rect 14549 3032 14554 3088
rect 14610 3032 15762 3088
rect 14549 3030 15762 3032
rect 15837 3090 15903 3093
rect 18505 3090 18571 3093
rect 23841 3090 23907 3093
rect 15837 3088 23907 3090
rect 15837 3032 15842 3088
rect 15898 3032 18510 3088
rect 18566 3032 23846 3088
rect 23902 3032 23907 3088
rect 15837 3030 23907 3032
rect 23982 3090 24042 3163
rect 27520 3136 28000 3166
rect 26233 3090 26299 3093
rect 23982 3088 26299 3090
rect 23982 3032 26238 3088
rect 26294 3032 26299 3088
rect 23982 3030 26299 3032
rect 14549 3027 14615 3030
rect 15837 3027 15903 3030
rect 18505 3027 18571 3030
rect 23841 3027 23907 3030
rect 26233 3027 26299 3030
rect 2957 2954 3023 2957
rect 3785 2954 3851 2957
rect 8569 2954 8635 2957
rect 2957 2952 8635 2954
rect 2957 2896 2962 2952
rect 3018 2896 3790 2952
rect 3846 2896 8574 2952
rect 8630 2896 8635 2952
rect 2957 2894 8635 2896
rect 2957 2891 3023 2894
rect 3785 2891 3851 2894
rect 8569 2891 8635 2894
rect 8753 2954 8819 2957
rect 13854 2954 13860 2956
rect 8753 2952 13860 2954
rect 8753 2896 8758 2952
rect 8814 2896 13860 2952
rect 8753 2894 13860 2896
rect 8753 2891 8819 2894
rect 13854 2892 13860 2894
rect 13924 2892 13930 2956
rect 13997 2954 14063 2957
rect 17401 2954 17467 2957
rect 13997 2952 17467 2954
rect 13997 2896 14002 2952
rect 14058 2896 17406 2952
rect 17462 2896 17467 2952
rect 13997 2894 17467 2896
rect 13997 2891 14063 2894
rect 17401 2891 17467 2894
rect 17534 2892 17540 2956
rect 17604 2954 17610 2956
rect 20713 2954 20779 2957
rect 17604 2952 20779 2954
rect 17604 2896 20718 2952
rect 20774 2896 20779 2952
rect 17604 2894 20779 2896
rect 17604 2892 17610 2894
rect 20713 2891 20779 2894
rect 21081 2954 21147 2957
rect 25129 2954 25195 2957
rect 21081 2952 25195 2954
rect 21081 2896 21086 2952
rect 21142 2896 25134 2952
rect 25190 2896 25195 2952
rect 21081 2894 25195 2896
rect 21081 2891 21147 2894
rect 25129 2891 25195 2894
rect 7925 2818 7991 2821
rect 9765 2818 9831 2821
rect 7925 2816 9831 2818
rect 7925 2760 7930 2816
rect 7986 2760 9770 2816
rect 9826 2760 9831 2816
rect 7925 2758 9831 2760
rect 7925 2755 7991 2758
rect 9765 2755 9831 2758
rect 13629 2818 13695 2821
rect 18045 2818 18111 2821
rect 13629 2816 18111 2818
rect 13629 2760 13634 2816
rect 13690 2760 18050 2816
rect 18106 2760 18111 2816
rect 13629 2758 18111 2760
rect 13629 2755 13695 2758
rect 18045 2755 18111 2758
rect 24025 2818 24091 2821
rect 25221 2818 25287 2821
rect 24025 2816 25287 2818
rect 24025 2760 24030 2816
rect 24086 2760 25226 2816
rect 25282 2760 25287 2816
rect 24025 2758 25287 2760
rect 24025 2755 24091 2758
rect 25221 2755 25287 2758
rect 10277 2752 10597 2753
rect 0 2682 480 2712
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 9213 2682 9279 2685
rect 0 2680 9279 2682
rect 0 2624 9218 2680
rect 9274 2624 9279 2680
rect 0 2622 9279 2624
rect 0 2592 480 2622
rect 9213 2619 9279 2622
rect 10685 2682 10751 2685
rect 13537 2682 13603 2685
rect 19425 2682 19491 2685
rect 10685 2680 11530 2682
rect 10685 2624 10690 2680
rect 10746 2624 11530 2680
rect 10685 2622 11530 2624
rect 10685 2619 10751 2622
rect 3693 2546 3759 2549
rect 8661 2546 8727 2549
rect 11237 2546 11303 2549
rect 3693 2544 6562 2546
rect 3693 2488 3698 2544
rect 3754 2488 6562 2544
rect 3693 2486 6562 2488
rect 3693 2483 3759 2486
rect 6502 2410 6562 2486
rect 8661 2544 11303 2546
rect 8661 2488 8666 2544
rect 8722 2488 11242 2544
rect 11298 2488 11303 2544
rect 8661 2486 11303 2488
rect 11470 2546 11530 2622
rect 13537 2680 19491 2682
rect 13537 2624 13542 2680
rect 13598 2624 19430 2680
rect 19486 2624 19491 2680
rect 13537 2622 19491 2624
rect 13537 2619 13603 2622
rect 19425 2619 19491 2622
rect 20069 2682 20135 2685
rect 22277 2682 22343 2685
rect 20069 2680 22343 2682
rect 20069 2624 20074 2680
rect 20130 2624 22282 2680
rect 22338 2624 22343 2680
rect 20069 2622 22343 2624
rect 20069 2619 20135 2622
rect 22277 2619 22343 2622
rect 23105 2682 23171 2685
rect 27520 2682 28000 2712
rect 23105 2680 28000 2682
rect 23105 2624 23110 2680
rect 23166 2624 28000 2680
rect 23105 2622 28000 2624
rect 23105 2619 23171 2622
rect 27520 2592 28000 2622
rect 17309 2546 17375 2549
rect 11470 2544 17375 2546
rect 11470 2488 17314 2544
rect 17370 2488 17375 2544
rect 11470 2486 17375 2488
rect 8661 2483 8727 2486
rect 11237 2483 11303 2486
rect 17309 2483 17375 2486
rect 17493 2546 17559 2549
rect 21909 2546 21975 2549
rect 24485 2546 24551 2549
rect 26417 2546 26483 2549
rect 17493 2544 20730 2546
rect 17493 2488 17498 2544
rect 17554 2488 20730 2544
rect 17493 2486 20730 2488
rect 17493 2483 17559 2486
rect 10593 2410 10659 2413
rect 6502 2408 10659 2410
rect 6502 2352 10598 2408
rect 10654 2352 10659 2408
rect 6502 2350 10659 2352
rect 10593 2347 10659 2350
rect 10777 2410 10843 2413
rect 14549 2410 14615 2413
rect 20529 2410 20595 2413
rect 10777 2408 14615 2410
rect 10777 2352 10782 2408
rect 10838 2352 14554 2408
rect 14610 2352 14615 2408
rect 10777 2350 14615 2352
rect 10777 2347 10843 2350
rect 14549 2347 14615 2350
rect 14782 2408 20595 2410
rect 14782 2352 20534 2408
rect 20590 2352 20595 2408
rect 14782 2350 20595 2352
rect 20670 2410 20730 2486
rect 21909 2544 26483 2546
rect 21909 2488 21914 2544
rect 21970 2488 24490 2544
rect 24546 2488 26422 2544
rect 26478 2488 26483 2544
rect 21909 2486 26483 2488
rect 21909 2483 21975 2486
rect 24485 2483 24551 2486
rect 26417 2483 26483 2486
rect 22737 2412 22803 2413
rect 20670 2350 22570 2410
rect 1577 2274 1643 2277
rect 5390 2274 5396 2276
rect 1577 2272 5396 2274
rect 1577 2216 1582 2272
rect 1638 2216 5396 2272
rect 1577 2214 5396 2216
rect 1577 2211 1643 2214
rect 5390 2212 5396 2214
rect 5460 2212 5466 2276
rect 9581 2274 9647 2277
rect 14782 2274 14842 2350
rect 20529 2347 20595 2350
rect 9581 2272 14842 2274
rect 9581 2216 9586 2272
rect 9642 2216 14842 2272
rect 9581 2214 14842 2216
rect 17309 2274 17375 2277
rect 20897 2274 20963 2277
rect 17309 2272 20963 2274
rect 17309 2216 17314 2272
rect 17370 2216 20902 2272
rect 20958 2216 20963 2272
rect 17309 2214 20963 2216
rect 22510 2274 22570 2350
rect 22686 2348 22692 2412
rect 22756 2410 22803 2412
rect 22756 2408 22848 2410
rect 22798 2352 22848 2408
rect 22756 2350 22848 2352
rect 22756 2348 22803 2350
rect 22737 2347 22803 2348
rect 23933 2274 23999 2277
rect 22510 2272 23999 2274
rect 22510 2216 23938 2272
rect 23994 2216 23999 2272
rect 22510 2214 23999 2216
rect 9581 2211 9647 2214
rect 17309 2211 17375 2214
rect 20897 2211 20963 2214
rect 23933 2211 23999 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 5993 2138 6059 2141
rect 11973 2138 12039 2141
rect 5993 2136 12039 2138
rect 5993 2080 5998 2136
rect 6054 2080 11978 2136
rect 12034 2080 12039 2136
rect 5993 2078 12039 2080
rect 5993 2075 6059 2078
rect 11973 2075 12039 2078
rect 0 2002 480 2032
rect 4061 2002 4127 2005
rect 0 2000 4127 2002
rect 0 1944 4066 2000
rect 4122 1944 4127 2000
rect 0 1942 4127 1944
rect 0 1912 480 1942
rect 4061 1939 4127 1942
rect 10961 2002 11027 2005
rect 18689 2002 18755 2005
rect 20989 2002 21055 2005
rect 10961 2000 17418 2002
rect 10961 1944 10966 2000
rect 11022 1944 17418 2000
rect 10961 1942 17418 1944
rect 10961 1939 11027 1942
rect 1945 1866 2011 1869
rect 13261 1866 13327 1869
rect 1945 1864 13327 1866
rect 1945 1808 1950 1864
rect 2006 1808 13266 1864
rect 13322 1808 13327 1864
rect 1945 1806 13327 1808
rect 1945 1803 2011 1806
rect 13261 1803 13327 1806
rect 13721 1866 13787 1869
rect 16849 1866 16915 1869
rect 13721 1864 16915 1866
rect 13721 1808 13726 1864
rect 13782 1808 16854 1864
rect 16910 1808 16915 1864
rect 13721 1806 16915 1808
rect 13721 1803 13787 1806
rect 16849 1803 16915 1806
rect 197 1730 263 1733
rect 11053 1730 11119 1733
rect 197 1728 11119 1730
rect 197 1672 202 1728
rect 258 1672 11058 1728
rect 11114 1672 11119 1728
rect 197 1670 11119 1672
rect 197 1667 263 1670
rect 11053 1667 11119 1670
rect 11237 1730 11303 1733
rect 17358 1730 17418 1942
rect 18689 2000 21055 2002
rect 18689 1944 18694 2000
rect 18750 1944 20994 2000
rect 21050 1944 21055 2000
rect 18689 1942 21055 1944
rect 18689 1939 18755 1942
rect 20989 1939 21055 1942
rect 24710 1940 24716 2004
rect 24780 2002 24786 2004
rect 27520 2002 28000 2032
rect 24780 1942 28000 2002
rect 24780 1940 24786 1942
rect 27520 1912 28000 1942
rect 17493 1866 17559 1869
rect 25773 1866 25839 1869
rect 17493 1864 25839 1866
rect 17493 1808 17498 1864
rect 17554 1808 25778 1864
rect 25834 1808 25839 1864
rect 17493 1806 25839 1808
rect 17493 1803 17559 1806
rect 25773 1803 25839 1806
rect 22829 1730 22895 1733
rect 11237 1728 17234 1730
rect 11237 1672 11242 1728
rect 11298 1672 17234 1728
rect 11237 1670 17234 1672
rect 17358 1728 22895 1730
rect 17358 1672 22834 1728
rect 22890 1672 22895 1728
rect 17358 1670 22895 1672
rect 11237 1667 11303 1670
rect 4061 1594 4127 1597
rect 15101 1594 15167 1597
rect 4061 1592 15167 1594
rect 4061 1536 4066 1592
rect 4122 1536 15106 1592
rect 15162 1536 15167 1592
rect 4061 1534 15167 1536
rect 17174 1594 17234 1670
rect 22829 1667 22895 1670
rect 23933 1730 23999 1733
rect 26141 1730 26207 1733
rect 23933 1728 26207 1730
rect 23933 1672 23938 1728
rect 23994 1672 26146 1728
rect 26202 1672 26207 1728
rect 23933 1670 26207 1672
rect 23933 1667 23999 1670
rect 26141 1667 26207 1670
rect 24669 1594 24735 1597
rect 17174 1592 24735 1594
rect 17174 1536 24674 1592
rect 24730 1536 24735 1592
rect 17174 1534 24735 1536
rect 4061 1531 4127 1534
rect 15101 1531 15167 1534
rect 24669 1531 24735 1534
rect 0 1458 480 1488
rect 4337 1458 4403 1461
rect 4889 1458 4955 1461
rect 18321 1458 18387 1461
rect 0 1456 4403 1458
rect 0 1400 4342 1456
rect 4398 1400 4403 1456
rect 0 1398 4403 1400
rect 0 1368 480 1398
rect 4337 1395 4403 1398
rect 4478 1456 18387 1458
rect 4478 1400 4894 1456
rect 4950 1400 18326 1456
rect 18382 1400 18387 1456
rect 4478 1398 18387 1400
rect 2497 1322 2563 1325
rect 4478 1322 4538 1398
rect 4889 1395 4955 1398
rect 18321 1395 18387 1398
rect 19333 1458 19399 1461
rect 22921 1458 22987 1461
rect 19333 1456 22987 1458
rect 19333 1400 19338 1456
rect 19394 1400 22926 1456
rect 22982 1400 22987 1456
rect 19333 1398 22987 1400
rect 19333 1395 19399 1398
rect 22921 1395 22987 1398
rect 23565 1458 23631 1461
rect 27520 1458 28000 1488
rect 23565 1456 28000 1458
rect 23565 1400 23570 1456
rect 23626 1400 28000 1456
rect 23565 1398 28000 1400
rect 23565 1395 23631 1398
rect 27520 1368 28000 1398
rect 2497 1320 4538 1322
rect 2497 1264 2502 1320
rect 2558 1264 4538 1320
rect 2497 1262 4538 1264
rect 6085 1322 6151 1325
rect 15193 1322 15259 1325
rect 18229 1322 18295 1325
rect 6085 1320 15259 1322
rect 6085 1264 6090 1320
rect 6146 1264 15198 1320
rect 15254 1264 15259 1320
rect 6085 1262 15259 1264
rect 2497 1259 2563 1262
rect 6085 1259 6151 1262
rect 15193 1259 15259 1262
rect 15334 1320 18295 1322
rect 15334 1264 18234 1320
rect 18290 1264 18295 1320
rect 15334 1262 18295 1264
rect 10593 1186 10659 1189
rect 10910 1186 10916 1188
rect 10593 1184 10916 1186
rect 10593 1128 10598 1184
rect 10654 1128 10916 1184
rect 10593 1126 10916 1128
rect 10593 1123 10659 1126
rect 10910 1124 10916 1126
rect 10980 1124 10986 1188
rect 11421 1186 11487 1189
rect 15334 1186 15394 1262
rect 18229 1259 18295 1262
rect 18413 1322 18479 1325
rect 25037 1322 25103 1325
rect 18413 1320 25103 1322
rect 18413 1264 18418 1320
rect 18474 1264 25042 1320
rect 25098 1264 25103 1320
rect 18413 1262 25103 1264
rect 18413 1259 18479 1262
rect 25037 1259 25103 1262
rect 17309 1186 17375 1189
rect 11421 1184 15394 1186
rect 11421 1128 11426 1184
rect 11482 1128 15394 1184
rect 11421 1126 15394 1128
rect 16990 1184 17375 1186
rect 16990 1128 17314 1184
rect 17370 1128 17375 1184
rect 16990 1126 17375 1128
rect 11421 1123 11487 1126
rect 9765 1050 9831 1053
rect 16990 1050 17050 1126
rect 17309 1123 17375 1126
rect 24025 1050 24091 1053
rect 9765 1048 17050 1050
rect 9765 992 9770 1048
rect 9826 992 17050 1048
rect 9765 990 17050 992
rect 17174 1048 24091 1050
rect 17174 992 24030 1048
rect 24086 992 24091 1048
rect 17174 990 24091 992
rect 9765 987 9831 990
rect 0 914 480 944
rect 4061 914 4127 917
rect 0 912 4127 914
rect 0 856 4066 912
rect 4122 856 4127 912
rect 0 854 4127 856
rect 0 824 480 854
rect 4061 851 4127 854
rect 7189 914 7255 917
rect 17174 914 17234 990
rect 24025 987 24091 990
rect 7189 912 17234 914
rect 7189 856 7194 912
rect 7250 856 17234 912
rect 7189 854 17234 856
rect 17401 914 17467 917
rect 27520 914 28000 944
rect 17401 912 28000 914
rect 17401 856 17406 912
rect 17462 856 28000 912
rect 17401 854 28000 856
rect 7189 851 7255 854
rect 17401 851 17467 854
rect 27520 824 28000 854
rect 1485 778 1551 781
rect 11881 778 11947 781
rect 17309 778 17375 781
rect 23381 778 23447 781
rect 1485 776 7666 778
rect 1485 720 1490 776
rect 1546 720 7666 776
rect 1485 718 7666 720
rect 1485 715 1551 718
rect 7465 642 7531 645
rect 614 640 7531 642
rect 614 584 7470 640
rect 7526 584 7531 640
rect 614 582 7531 584
rect 7606 642 7666 718
rect 11881 776 17234 778
rect 11881 720 11886 776
rect 11942 720 17234 776
rect 11881 718 17234 720
rect 11881 715 11947 718
rect 17033 642 17099 645
rect 7606 640 17099 642
rect 7606 584 17038 640
rect 17094 584 17099 640
rect 7606 582 17099 584
rect 17174 642 17234 718
rect 17309 776 23447 778
rect 17309 720 17314 776
rect 17370 720 23386 776
rect 23442 720 23447 776
rect 17309 718 23447 720
rect 17309 715 17375 718
rect 23381 715 23447 718
rect 24761 642 24827 645
rect 17174 640 24827 642
rect 17174 584 24766 640
rect 24822 584 24827 640
rect 17174 582 24827 584
rect 0 370 480 400
rect 614 370 674 582
rect 7465 579 7531 582
rect 17033 579 17099 582
rect 24761 579 24827 582
rect 6269 506 6335 509
rect 26049 506 26115 509
rect 6269 504 26115 506
rect 6269 448 6274 504
rect 6330 448 26054 504
rect 26110 448 26115 504
rect 6269 446 26115 448
rect 6269 443 6335 446
rect 26049 443 26115 446
rect 0 310 674 370
rect 3877 370 3943 373
rect 4981 370 5047 373
rect 15193 370 15259 373
rect 19425 370 19491 373
rect 3877 368 15026 370
rect 3877 312 3882 368
rect 3938 312 4986 368
rect 5042 312 15026 368
rect 3877 310 15026 312
rect 0 280 480 310
rect 3877 307 3943 310
rect 4981 307 5047 310
rect 4061 234 4127 237
rect 14825 234 14891 237
rect 4061 232 14891 234
rect 4061 176 4066 232
rect 4122 176 14830 232
rect 14886 176 14891 232
rect 4061 174 14891 176
rect 4061 171 4127 174
rect 14825 171 14891 174
rect 14966 98 15026 310
rect 15193 368 19491 370
rect 15193 312 15198 368
rect 15254 312 19430 368
rect 19486 312 19491 368
rect 15193 310 19491 312
rect 15193 307 15259 310
rect 19425 307 19491 310
rect 23289 370 23355 373
rect 27520 370 28000 400
rect 23289 368 28000 370
rect 23289 312 23294 368
rect 23350 312 28000 368
rect 23289 310 28000 312
rect 23289 307 23355 310
rect 27520 280 28000 310
rect 17033 234 17099 237
rect 23790 234 23796 236
rect 17033 232 23796 234
rect 17033 176 17038 232
rect 17094 176 23796 232
rect 17033 174 23796 176
rect 17033 171 17099 174
rect 23790 172 23796 174
rect 23860 172 23866 236
rect 20161 98 20227 101
rect 14966 96 20227 98
rect 14966 40 20166 96
rect 20222 40 20227 96
rect 14966 38 20227 40
rect 20161 35 20227 38
<< via3 >>
rect 21956 26556 22020 26620
rect 21036 26420 21100 26484
rect 12940 26284 13004 26348
rect 23612 26284 23676 26348
rect 3004 26148 3068 26212
rect 25084 26012 25148 26076
rect 3740 25876 3804 25940
rect 22324 25876 22388 25940
rect 2452 25740 2516 25804
rect 12204 25604 12268 25668
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 19380 25468 19444 25532
rect 25820 25468 25884 25532
rect 9628 25196 9692 25260
rect 21220 25332 21284 25396
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 23796 25060 23860 25124
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 1532 24652 1596 24716
rect 11100 24516 11164 24580
rect 14780 24788 14844 24852
rect 23428 24924 23492 24988
rect 16068 24788 16132 24852
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 17172 24380 17236 24444
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 2820 23836 2884 23900
rect 1900 23760 1964 23764
rect 1900 23704 1950 23760
rect 1950 23704 1964 23760
rect 1900 23700 1964 23704
rect 21404 23972 21468 24036
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 21772 23428 21836 23492
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 1900 22204 1964 22268
rect 3188 22204 3252 22268
rect 9444 22204 9508 22268
rect 23980 22204 24044 22268
rect 23980 21932 24044 21996
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 23980 21720 24044 21724
rect 23980 21664 23994 21720
rect 23994 21664 24044 21720
rect 23980 21660 24044 21664
rect 17172 21252 17236 21316
rect 20300 21388 20364 21452
rect 25268 21388 25332 21452
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 1900 21116 1964 21180
rect 5396 21116 5460 21180
rect 9812 20844 9876 20908
rect 20116 20708 20180 20772
rect 20852 20708 20916 20772
rect 23980 20768 24044 20772
rect 23980 20712 24030 20768
rect 24030 20712 24044 20768
rect 23980 20708 24044 20712
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 9996 20224 10060 20228
rect 9996 20168 10046 20224
rect 10046 20168 10060 20224
rect 9996 20164 10060 20168
rect 21220 20164 21284 20228
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 10732 20028 10796 20092
rect 12940 20088 13004 20092
rect 12940 20032 12954 20088
rect 12954 20032 13004 20088
rect 12940 20028 13004 20032
rect 22692 20088 22756 20092
rect 22692 20032 22742 20088
rect 22742 20032 22756 20088
rect 22692 20028 22756 20032
rect 9628 19892 9692 19956
rect 24900 19892 24964 19956
rect 22324 19756 22388 19820
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 21772 19484 21836 19548
rect 4476 19212 4540 19276
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 2820 19000 2884 19004
rect 2820 18944 2834 19000
rect 2834 18944 2884 19000
rect 2820 18940 2884 18944
rect 14780 18940 14844 19004
rect 5396 18804 5460 18868
rect 11468 18804 11532 18868
rect 7788 18668 7852 18732
rect 15884 18668 15948 18732
rect 22876 18668 22940 18732
rect 23980 18668 24044 18732
rect 20300 18532 20364 18596
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 7052 17988 7116 18052
rect 22324 17988 22388 18052
rect 23612 17988 23676 18052
rect 24716 17988 24780 18052
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5212 17912 5276 17916
rect 5212 17856 5226 17912
rect 5226 17856 5276 17912
rect 5212 17852 5276 17856
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 2820 17308 2884 17372
rect 13124 17368 13188 17372
rect 13124 17312 13138 17368
rect 13138 17312 13188 17368
rect 13124 17308 13188 17312
rect 23060 17172 23124 17236
rect 5212 16900 5276 16964
rect 19196 17036 19260 17100
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 4844 16764 4908 16828
rect 13860 16688 13924 16692
rect 13860 16632 13910 16688
rect 13910 16632 13924 16688
rect 13860 16628 13924 16632
rect 21772 16492 21836 16556
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 1532 16084 1596 16148
rect 11100 16084 11164 16148
rect 12020 16084 12084 16148
rect 14780 16220 14844 16284
rect 21956 16144 22020 16148
rect 21956 16088 22006 16144
rect 22006 16088 22020 16144
rect 21956 16084 22020 16088
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5396 15540 5460 15604
rect 22140 15464 22204 15468
rect 22140 15408 22154 15464
rect 22154 15408 22204 15464
rect 22140 15404 22204 15408
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 7788 15192 7852 15196
rect 7788 15136 7802 15192
rect 7802 15136 7852 15192
rect 7788 15132 7852 15136
rect 19380 15132 19444 15196
rect 21956 15268 22020 15332
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 13676 14996 13740 15060
rect 6316 14784 6380 14788
rect 6316 14728 6366 14784
rect 6366 14728 6380 14784
rect 6316 14724 6380 14728
rect 23060 14724 23124 14788
rect 25636 14724 25700 14788
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 12020 14588 12084 14652
rect 20300 14588 20364 14652
rect 23612 14588 23676 14652
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 9260 13968 9324 13972
rect 9260 13912 9310 13968
rect 9310 13912 9324 13968
rect 9260 13908 9324 13912
rect 14412 13908 14476 13972
rect 15332 13772 15396 13836
rect 20484 13772 20548 13836
rect 10916 13636 10980 13700
rect 14596 13636 14660 13700
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 23060 13228 23124 13292
rect 24716 13228 24780 13292
rect 25268 13228 25332 13292
rect 13492 13092 13556 13156
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 9996 12956 10060 13020
rect 10916 12956 10980 13020
rect 16068 13016 16132 13020
rect 16068 12960 16118 13016
rect 16118 12960 16132 13016
rect 16068 12956 16132 12960
rect 22692 12820 22756 12884
rect 25268 12820 25332 12884
rect 11468 12684 11532 12748
rect 10916 12548 10980 12612
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 2452 12200 2516 12204
rect 2452 12144 2466 12200
rect 2466 12144 2516 12200
rect 2452 12140 2516 12144
rect 6500 12200 6564 12204
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 6500 12144 6514 12200
rect 6514 12144 6564 12200
rect 6500 12140 6564 12144
rect 12020 12276 12084 12340
rect 16436 12412 16500 12476
rect 19196 12412 19260 12476
rect 25820 12276 25884 12340
rect 9260 12004 9324 12068
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 23612 12004 23676 12068
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 21404 11928 21468 11932
rect 21404 11872 21454 11928
rect 21454 11872 21468 11928
rect 21404 11868 21468 11872
rect 22140 11868 22204 11932
rect 6316 11596 6380 11660
rect 2820 11520 2884 11524
rect 2820 11464 2870 11520
rect 2870 11464 2884 11520
rect 2820 11460 2884 11464
rect 3924 11324 3988 11388
rect 22324 11596 22388 11660
rect 16804 11460 16868 11524
rect 19196 11520 19260 11524
rect 19196 11464 19246 11520
rect 19246 11464 19260 11520
rect 19196 11460 19260 11464
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 14596 11324 14660 11388
rect 15516 11324 15580 11388
rect 11284 11188 11348 11252
rect 21956 11324 22020 11388
rect 3924 11052 3988 11116
rect 16988 11052 17052 11116
rect 19380 11052 19444 11116
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 2084 10568 2148 10572
rect 2084 10512 2098 10568
rect 2098 10512 2148 10568
rect 2084 10508 2148 10512
rect 20484 10780 20548 10844
rect 25084 10976 25148 10980
rect 25084 10920 25098 10976
rect 25098 10920 25148 10976
rect 25084 10916 25148 10920
rect 26372 10916 26436 10980
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 10916 10236 10980 10300
rect 20300 10236 20364 10300
rect 5396 9888 5460 9892
rect 5396 9832 5410 9888
rect 5410 9832 5460 9888
rect 5396 9828 5460 9832
rect 6684 9828 6748 9892
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 7788 9692 7852 9756
rect 15332 9964 15396 10028
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 1716 9616 1780 9620
rect 1716 9560 1766 9616
rect 1766 9560 1780 9616
rect 1716 9556 1780 9560
rect 23428 9556 23492 9620
rect 24900 9556 24964 9620
rect 25452 9616 25516 9620
rect 25452 9560 25466 9616
rect 25466 9560 25516 9616
rect 25452 9556 25516 9560
rect 26004 9616 26068 9620
rect 26004 9560 26018 9616
rect 26018 9560 26068 9616
rect 26004 9556 26068 9560
rect 11100 9420 11164 9484
rect 14412 9284 14476 9348
rect 25268 9420 25332 9484
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 3004 9148 3068 9212
rect 9628 9148 9692 9212
rect 10916 9148 10980 9212
rect 20668 9148 20732 9212
rect 26740 9148 26804 9212
rect 4844 8740 4908 8804
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 20116 8876 20180 8940
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 3188 8528 3252 8532
rect 3188 8472 3202 8528
rect 3202 8472 3252 8528
rect 3188 8468 3252 8472
rect 4476 8468 4540 8532
rect 5212 8468 5276 8532
rect 12020 8528 12084 8532
rect 12020 8472 12070 8528
rect 12070 8472 12084 8528
rect 12020 8468 12084 8472
rect 19196 8740 19260 8804
rect 23796 8800 23860 8804
rect 23796 8744 23846 8800
rect 23846 8744 23860 8800
rect 23796 8740 23860 8744
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 21956 8332 22020 8396
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 25636 8060 25700 8124
rect 3004 7848 3068 7852
rect 3004 7792 3018 7848
rect 3018 7792 3068 7848
rect 3004 7788 3068 7792
rect 6500 7788 6564 7852
rect 24900 7788 24964 7852
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 7420 7516 7484 7580
rect 5212 7440 5276 7444
rect 5212 7384 5226 7440
rect 5226 7384 5276 7440
rect 5212 7380 5276 7384
rect 19380 7380 19444 7444
rect 3740 6972 3804 7036
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 26188 7108 26252 7172
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 4844 6836 4908 6900
rect 6132 6760 6196 6764
rect 6132 6704 6146 6760
rect 6146 6704 6196 6760
rect 6132 6700 6196 6704
rect 24900 6972 24964 7036
rect 18092 6836 18156 6900
rect 21772 6836 21836 6900
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 8156 6488 8220 6492
rect 8156 6432 8170 6488
rect 8170 6432 8220 6488
rect 8156 6428 8220 6432
rect 9812 6428 9876 6492
rect 10732 6428 10796 6492
rect 12204 6428 12268 6492
rect 17908 6428 17972 6492
rect 20852 6292 20916 6356
rect 21772 6292 21836 6356
rect 23428 6292 23492 6356
rect 17724 6156 17788 6220
rect 7420 6020 7484 6084
rect 13308 6020 13372 6084
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 7236 5536 7300 5540
rect 7236 5480 7250 5536
rect 7250 5480 7300 5536
rect 7236 5476 7300 5480
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 9628 5340 9692 5404
rect 17724 5340 17788 5404
rect 23980 5400 24044 5404
rect 23980 5344 24030 5400
rect 24030 5344 24044 5400
rect 23980 5340 24044 5344
rect 9996 5068 10060 5132
rect 15516 4932 15580 4996
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 9996 4388 10060 4452
rect 20116 4388 20180 4452
rect 20668 4388 20732 4452
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 11100 4116 11164 4180
rect 21036 3844 21100 3908
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 6132 3708 6196 3772
rect 9444 3708 9508 3772
rect 13676 3708 13740 3772
rect 21772 3708 21836 3772
rect 14412 3496 14476 3500
rect 14412 3440 14426 3496
rect 14426 3440 14476 3496
rect 14412 3436 14476 3440
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 14412 3224 14476 3228
rect 14412 3168 14462 3224
rect 14462 3168 14476 3224
rect 14412 3164 14476 3168
rect 6684 3028 6748 3092
rect 23428 3300 23492 3364
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 13860 2892 13924 2956
rect 17540 2892 17604 2956
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5396 2212 5460 2276
rect 22692 2408 22756 2412
rect 22692 2352 22742 2408
rect 22742 2352 22756 2408
rect 22692 2348 22756 2352
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 24716 1940 24780 2004
rect 10916 1124 10980 1188
rect 23796 172 23860 236
<< metal4 >>
rect 21955 26620 22021 26621
rect 21955 26556 21956 26620
rect 22020 26556 22021 26620
rect 21955 26555 22021 26556
rect 21035 26484 21101 26485
rect 21035 26420 21036 26484
rect 21100 26420 21101 26484
rect 21035 26419 21101 26420
rect 12939 26348 13005 26349
rect 12939 26284 12940 26348
rect 13004 26284 13005 26348
rect 12939 26283 13005 26284
rect 3003 26212 3069 26213
rect 3003 26148 3004 26212
rect 3068 26148 3069 26212
rect 3003 26147 3069 26148
rect 2451 25804 2517 25805
rect 2451 25740 2452 25804
rect 2516 25740 2517 25804
rect 2451 25739 2517 25740
rect 1531 24716 1597 24717
rect 1531 24652 1532 24716
rect 1596 24652 1597 24716
rect 1531 24651 1597 24652
rect 1534 22898 1594 24651
rect 1899 23764 1965 23765
rect 1899 23700 1900 23764
rect 1964 23700 1965 23764
rect 1899 23699 1965 23700
rect 1534 16149 1594 22662
rect 1902 22269 1962 23699
rect 1899 22268 1965 22269
rect 1899 22204 1900 22268
rect 1964 22204 1965 22268
rect 1899 22203 1965 22204
rect 1899 21180 1965 21181
rect 1899 21116 1900 21180
rect 1964 21116 1965 21180
rect 1899 21115 1965 21116
rect 1531 16148 1597 16149
rect 1531 16084 1532 16148
rect 1596 16084 1597 16148
rect 1531 16083 1597 16084
rect 1902 11250 1962 21115
rect 2454 12205 2514 25739
rect 2819 23900 2885 23901
rect 2819 23836 2820 23900
rect 2884 23836 2885 23900
rect 2819 23835 2885 23836
rect 2822 19005 2882 23835
rect 2819 19004 2885 19005
rect 2819 18940 2820 19004
rect 2884 18940 2885 19004
rect 2819 18939 2885 18940
rect 2819 17372 2885 17373
rect 2819 17308 2820 17372
rect 2884 17308 2885 17372
rect 2819 17307 2885 17308
rect 2451 12204 2517 12205
rect 2451 12140 2452 12204
rect 2516 12140 2517 12204
rect 2451 12139 2517 12140
rect 2822 11525 2882 17307
rect 2819 11524 2885 11525
rect 2819 11460 2820 11524
rect 2884 11460 2885 11524
rect 2819 11459 2885 11460
rect 1718 11190 1962 11250
rect 1718 9621 1778 11190
rect 1715 9620 1781 9621
rect 1715 9556 1716 9620
rect 1780 9556 1781 9620
rect 1715 9555 1781 9556
rect 3006 9213 3066 26147
rect 3739 25940 3805 25941
rect 3739 25876 3740 25940
rect 3804 25876 3805 25940
rect 3739 25875 3805 25876
rect 3187 22268 3253 22269
rect 3187 22204 3188 22268
rect 3252 22204 3253 22268
rect 3187 22203 3253 22204
rect 3003 9212 3069 9213
rect 3003 9148 3004 9212
rect 3068 9148 3069 9212
rect 3003 9147 3069 9148
rect 3190 8533 3250 22203
rect 3187 8532 3253 8533
rect 3187 8468 3188 8532
rect 3252 8468 3253 8532
rect 3187 8467 3253 8468
rect 3742 7037 3802 25875
rect 12203 25668 12269 25669
rect 5398 21181 5458 25382
rect 5610 25056 5931 25616
rect 10277 25600 10597 25616
rect 12203 25604 12204 25668
rect 12268 25604 12269 25668
rect 12203 25603 12269 25604
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 9627 25260 9693 25261
rect 9627 25258 9628 25260
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 9446 25198 9628 25258
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5395 21180 5461 21181
rect 5395 21116 5396 21180
rect 5460 21116 5461 21180
rect 5395 21115 5461 21116
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 4475 19276 4541 19277
rect 4475 19212 4476 19276
rect 4540 19212 4541 19276
rect 4475 19211 4541 19212
rect 3923 11388 3989 11389
rect 3923 11324 3924 11388
rect 3988 11324 3989 11388
rect 3923 11323 3989 11324
rect 3926 11117 3986 11323
rect 3923 11116 3989 11117
rect 3923 11052 3924 11116
rect 3988 11052 3989 11116
rect 3923 11051 3989 11052
rect 4478 8533 4538 19211
rect 5398 18869 5458 20622
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5395 18868 5461 18869
rect 5395 18804 5396 18868
rect 5460 18804 5461 18868
rect 5395 18803 5461 18804
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5211 17916 5277 17917
rect 5211 17852 5212 17916
rect 5276 17852 5277 17916
rect 5211 17851 5277 17852
rect 5214 16965 5274 17851
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5211 16964 5277 16965
rect 5211 16900 5212 16964
rect 5276 16900 5277 16964
rect 5211 16899 5277 16900
rect 4843 16828 4909 16829
rect 4843 16764 4844 16828
rect 4908 16764 4909 16828
rect 5214 16778 5274 16899
rect 4843 16763 4909 16764
rect 4846 12698 4906 16763
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5395 15604 5461 15605
rect 5395 15540 5396 15604
rect 5460 15540 5461 15604
rect 5395 15539 5461 15540
rect 4846 8805 4906 12462
rect 5398 9893 5458 15539
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5395 9892 5461 9893
rect 5395 9828 5396 9892
rect 5460 9828 5461 9892
rect 5395 9827 5461 9828
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 4843 8804 4909 8805
rect 4843 8740 4844 8804
rect 4908 8740 4909 8804
rect 4843 8739 4909 8740
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 4475 8532 4541 8533
rect 4475 8468 4476 8532
rect 4540 8468 4541 8532
rect 4475 8467 4541 8468
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5211 7444 5277 7445
rect 5211 7380 5212 7444
rect 5276 7380 5277 7444
rect 5211 7379 5277 7380
rect 5214 7258 5274 7379
rect 3739 7036 3805 7037
rect 3739 6972 3740 7036
rect 3804 6972 3805 7036
rect 3739 6971 3805 6972
rect 4843 6900 4909 6901
rect 4843 6836 4844 6900
rect 4908 6836 4909 6900
rect 4843 6835 4909 6836
rect 4846 1138 4906 6835
rect 5610 6560 5931 7584
rect 6134 6765 6194 21982
rect 6315 14788 6381 14789
rect 6315 14724 6316 14788
rect 6380 14724 6381 14788
rect 6315 14723 6381 14724
rect 6318 11661 6378 14723
rect 6499 12204 6565 12205
rect 6499 12140 6500 12204
rect 6564 12140 6565 12204
rect 6499 12139 6565 12140
rect 6315 11660 6381 11661
rect 6315 11596 6316 11660
rect 6380 11596 6381 11660
rect 6315 11595 6381 11596
rect 6502 7853 6562 12139
rect 6686 9893 6746 24702
rect 9446 22269 9506 25198
rect 9627 25196 9628 25198
rect 9692 25196 9693 25260
rect 9627 25195 9693 25196
rect 10277 24512 10597 25536
rect 11099 24580 11165 24581
rect 11099 24516 11100 24580
rect 11164 24516 11165 24580
rect 11099 24515 11165 24516
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 9443 22268 9509 22269
rect 9443 22204 9444 22268
rect 9508 22204 9509 22268
rect 9443 22203 9509 22204
rect 9814 20909 9874 21302
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 9811 20908 9877 20909
rect 9811 20844 9812 20908
rect 9876 20844 9877 20908
rect 9811 20843 9877 20844
rect 9627 19956 9693 19957
rect 9627 19892 9628 19956
rect 9692 19892 9693 19956
rect 9627 19891 9693 19892
rect 7051 18052 7117 18053
rect 7051 17988 7052 18052
rect 7116 17988 7117 18052
rect 7051 17987 7117 17988
rect 7054 12018 7114 17987
rect 6683 9892 6749 9893
rect 6683 9828 6684 9892
rect 6748 9828 6749 9892
rect 6683 9827 6749 9828
rect 7054 9754 7114 11782
rect 7054 9694 7298 9754
rect 6499 7852 6565 7853
rect 6499 7788 6500 7852
rect 6564 7788 6565 7852
rect 6499 7787 6565 7788
rect 6131 6764 6197 6765
rect 6131 6700 6132 6764
rect 6196 6700 6197 6764
rect 6131 6699 6197 6700
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 7238 5541 7298 9694
rect 7422 7581 7482 19262
rect 7787 18732 7853 18733
rect 7787 18668 7788 18732
rect 7852 18668 7853 18732
rect 7787 18667 7853 18668
rect 7790 18138 7850 18667
rect 7790 15197 7850 17902
rect 7787 15196 7853 15197
rect 7787 15132 7788 15196
rect 7852 15132 7853 15196
rect 7787 15131 7853 15132
rect 9259 13972 9325 13973
rect 9259 13908 9260 13972
rect 9324 13908 9325 13972
rect 9259 13907 9325 13908
rect 9262 12069 9322 13907
rect 9259 12068 9325 12069
rect 9259 12004 9260 12068
rect 9324 12004 9325 12068
rect 9259 12003 9325 12004
rect 7787 9692 7788 9742
rect 7852 9692 7853 9742
rect 7787 9691 7853 9692
rect 9630 9213 9690 19891
rect 9627 9212 9693 9213
rect 9627 9148 9628 9212
rect 9692 9148 9693 9212
rect 9627 9147 9693 9148
rect 7419 7580 7485 7581
rect 7419 7516 7420 7580
rect 7484 7516 7485 7580
rect 7419 7515 7485 7516
rect 7422 6085 7482 7515
rect 9814 6493 9874 20843
rect 9995 20228 10061 20229
rect 9995 20164 9996 20228
rect 10060 20164 10061 20228
rect 9995 20163 10061 20164
rect 9998 13021 10058 20163
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10731 20092 10797 20093
rect 10731 20028 10732 20092
rect 10796 20028 10797 20092
rect 10731 20027 10797 20028
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 9995 13020 10061 13021
rect 9995 12956 9996 13020
rect 10060 12956 10061 13020
rect 9995 12955 10061 12956
rect 9811 6492 9877 6493
rect 9811 6428 9812 6492
rect 9876 6428 9877 6492
rect 9811 6427 9877 6428
rect 7419 6084 7485 6085
rect 7419 6020 7420 6084
rect 7484 6020 7485 6084
rect 7419 6019 7485 6020
rect 7235 5540 7301 5541
rect 7235 5476 7236 5540
rect 7300 5476 7301 5540
rect 7235 5475 7301 5476
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 9627 5404 9693 5405
rect 9627 5340 9628 5404
rect 9692 5340 9693 5404
rect 9627 5339 9693 5340
rect 9630 5130 9690 5339
rect 9998 5133 10058 12955
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10734 6493 10794 20027
rect 11102 16149 11162 24515
rect 11467 18868 11533 18869
rect 11467 18818 11468 18868
rect 11532 18818 11533 18868
rect 11099 16148 11165 16149
rect 11099 16084 11100 16148
rect 11164 16084 11165 16148
rect 11099 16083 11165 16084
rect 11470 13970 11530 18582
rect 12019 16148 12085 16149
rect 12019 16084 12020 16148
rect 12084 16084 12085 16148
rect 12019 16083 12085 16084
rect 12022 14653 12082 16083
rect 12019 14652 12085 14653
rect 12019 14588 12020 14652
rect 12084 14588 12085 14652
rect 12019 14587 12085 14588
rect 11286 13910 11530 13970
rect 10915 13700 10981 13701
rect 10915 13636 10916 13700
rect 10980 13636 10981 13700
rect 10915 13635 10981 13636
rect 10918 13021 10978 13635
rect 10915 13020 10981 13021
rect 10915 12956 10916 13020
rect 10980 12956 10981 13020
rect 10915 12955 10981 12956
rect 10915 12612 10981 12613
rect 10915 12548 10916 12612
rect 10980 12548 10981 12612
rect 10915 12547 10981 12548
rect 10918 10301 10978 12547
rect 11286 11253 11346 13910
rect 11467 12748 11533 12749
rect 11467 12684 11468 12748
rect 11532 12684 11533 12748
rect 11467 12683 11533 12684
rect 11283 11252 11349 11253
rect 11283 11188 11284 11252
rect 11348 11188 11349 11252
rect 11283 11187 11349 11188
rect 11470 10658 11530 12683
rect 12019 12340 12085 12341
rect 12019 12276 12020 12340
rect 12084 12276 12085 12340
rect 12019 12275 12085 12276
rect 10915 10300 10981 10301
rect 10915 10236 10916 10300
rect 10980 10236 10981 10300
rect 10915 10235 10981 10236
rect 11099 9484 11165 9485
rect 11099 9420 11100 9484
rect 11164 9420 11165 9484
rect 11099 9419 11165 9420
rect 10915 9212 10981 9213
rect 10915 9148 10916 9212
rect 10980 9148 10981 9212
rect 10915 9147 10981 9148
rect 10731 6492 10797 6493
rect 10731 6428 10732 6492
rect 10796 6428 10797 6492
rect 10731 6427 10797 6428
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 9446 5070 9690 5130
rect 9995 5132 10061 5133
rect 9446 3773 9506 5070
rect 9995 5068 9996 5132
rect 10060 5068 10061 5132
rect 9995 5067 10061 5068
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 9443 3772 9509 3773
rect 9443 3708 9444 3772
rect 9508 3708 9509 3772
rect 9443 3707 9509 3708
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5395 2276 5461 2277
rect 5395 2212 5396 2276
rect 5460 2212 5461 2276
rect 5395 2211 5461 2212
rect 5398 1818 5458 2211
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 10918 1189 10978 9147
rect 11102 4181 11162 9419
rect 12022 8533 12082 12275
rect 12019 8532 12085 8533
rect 12019 8468 12020 8532
rect 12084 8468 12085 8532
rect 12019 8467 12085 8468
rect 12206 6493 12266 25603
rect 12942 20178 13002 26283
rect 14944 25056 15264 25616
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19379 25532 19445 25533
rect 19379 25468 19380 25532
rect 19444 25468 19445 25532
rect 19379 25467 19445 25468
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14779 24852 14845 24853
rect 14779 24788 14780 24852
rect 14844 24788 14845 24852
rect 14779 24787 14845 24788
rect 14782 19005 14842 24787
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14779 19004 14845 19005
rect 14779 18940 14780 19004
rect 14844 18940 14845 19004
rect 14779 18939 14845 18940
rect 14782 16285 14842 18939
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14779 16284 14845 16285
rect 14779 16220 14780 16284
rect 14844 16220 14845 16284
rect 14779 16219 14845 16220
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 13675 15060 13741 15061
rect 13675 14996 13676 15060
rect 13740 14996 13741 15060
rect 13675 14995 13741 14996
rect 13678 14058 13738 14995
rect 14414 13973 14474 14502
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14411 13972 14477 13973
rect 14411 13908 14412 13972
rect 14476 13908 14477 13972
rect 14411 13907 14477 13908
rect 14595 13700 14661 13701
rect 14595 13636 14596 13700
rect 14660 13636 14661 13700
rect 14595 13635 14661 13636
rect 13491 13092 13492 13142
rect 13556 13092 13557 13142
rect 13491 13091 13557 13092
rect 14598 12698 14658 13635
rect 14944 13088 15264 14112
rect 15331 13836 15397 13837
rect 15331 13772 15332 13836
rect 15396 13772 15397 13836
rect 15331 13771 15397 13772
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14598 11389 14658 12462
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14595 11388 14661 11389
rect 14595 11324 14596 11388
rect 14660 11324 14661 11388
rect 14595 11323 14661 11324
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 15334 10029 15394 13771
rect 15518 11389 15578 23342
rect 15883 18732 15949 18733
rect 15883 18668 15884 18732
rect 15948 18668 15949 18732
rect 15883 18667 15949 18668
rect 15886 12698 15946 18667
rect 16070 13021 16130 24702
rect 17171 24444 17237 24445
rect 17171 24380 17172 24444
rect 17236 24380 17237 24444
rect 17171 24379 17237 24380
rect 17174 21317 17234 24379
rect 17171 21316 17237 21317
rect 17171 21252 17172 21316
rect 17236 21252 17237 21316
rect 17171 21251 17237 21252
rect 16067 13020 16133 13021
rect 16067 12956 16068 13020
rect 16132 12956 16133 13020
rect 16067 12955 16133 12956
rect 16438 12477 16498 15182
rect 16435 12476 16501 12477
rect 16435 12412 16436 12476
rect 16500 12412 16501 12476
rect 16435 12411 16501 12412
rect 16806 11525 16866 17902
rect 19195 17100 19261 17101
rect 19195 17036 19196 17100
rect 19260 17036 19261 17100
rect 19195 17035 19261 17036
rect 19198 12477 19258 17035
rect 19382 15197 19442 25467
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 20299 18596 20365 18597
rect 20299 18532 20300 18596
rect 20364 18532 20365 18596
rect 20299 18531 20365 18532
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19379 15196 19445 15197
rect 19379 15132 19380 15196
rect 19444 15132 19445 15196
rect 19379 15131 19445 15132
rect 19195 12476 19261 12477
rect 19195 12412 19196 12476
rect 19260 12412 19261 12476
rect 19195 12411 19261 12412
rect 16803 11524 16869 11525
rect 16803 11460 16804 11524
rect 16868 11460 16869 11524
rect 16803 11459 16869 11460
rect 19195 11524 19261 11525
rect 19195 11460 19196 11524
rect 19260 11460 19261 11524
rect 19195 11459 19261 11460
rect 15515 11388 15581 11389
rect 15515 11324 15516 11388
rect 15580 11324 15581 11388
rect 15515 11323 15581 11324
rect 16987 11116 17053 11117
rect 16987 11052 16988 11116
rect 17052 11052 17053 11116
rect 16987 11051 17053 11052
rect 15331 10028 15397 10029
rect 15331 9964 15332 10028
rect 15396 9964 15397 10028
rect 16990 9978 17050 11051
rect 15331 9963 15397 9964
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14411 9348 14477 9349
rect 14411 9284 14412 9348
rect 14476 9284 14477 9348
rect 14411 9283 14477 9284
rect 12203 6492 12269 6493
rect 12203 6428 12204 6492
rect 12268 6428 12269 6492
rect 12203 6427 12269 6428
rect 13307 6084 13373 6085
rect 13307 6020 13308 6084
rect 13372 6020 13373 6084
rect 13307 6019 13373 6020
rect 11099 4180 11165 4181
rect 11099 4116 11100 4180
rect 11164 4116 11165 4180
rect 11099 4115 11165 4116
rect 13310 1818 13370 6019
rect 14414 3501 14474 9283
rect 14944 8736 15264 9760
rect 19198 8805 19258 11459
rect 19382 11117 19442 15131
rect 19610 14720 19930 15744
rect 20302 14738 20362 18531
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 20483 13836 20549 13837
rect 20483 13772 20484 13836
rect 20548 13772 20549 13836
rect 20483 13771 20549 13772
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19379 11116 19445 11117
rect 19379 11052 19380 11116
rect 19444 11052 19445 11116
rect 19379 11051 19445 11052
rect 19610 10368 19930 11392
rect 20486 10845 20546 13771
rect 20483 10844 20549 10845
rect 20483 10780 20484 10844
rect 20548 10780 20549 10844
rect 20483 10779 20549 10780
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 20299 10300 20365 10301
rect 20299 10236 20300 10300
rect 20364 10236 20365 10300
rect 20299 10235 20365 10236
rect 20302 9978 20362 10235
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19195 8804 19261 8805
rect 19195 8740 19196 8804
rect 19260 8740 19261 8804
rect 19195 8739 19261 8740
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 19382 7445 19442 8382
rect 19610 8192 19930 9216
rect 20670 9213 20730 22662
rect 20851 20772 20917 20773
rect 20851 20708 20852 20772
rect 20916 20708 20917 20772
rect 20851 20707 20917 20708
rect 20667 9212 20733 9213
rect 20667 9148 20668 9212
rect 20732 9148 20733 9212
rect 20667 9147 20733 9148
rect 20115 8940 20181 8941
rect 20115 8876 20116 8940
rect 20180 8876 20181 8940
rect 20115 8875 20181 8876
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19379 7444 19445 7445
rect 19379 7380 19380 7444
rect 19444 7380 19445 7444
rect 19379 7379 19445 7380
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 18091 6900 18157 6901
rect 18091 6836 18092 6900
rect 18156 6836 18157 6900
rect 18091 6835 18157 6836
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 17907 6492 17973 6493
rect 17907 6428 17908 6492
rect 17972 6490 17973 6492
rect 18094 6490 18154 6835
rect 17972 6430 18154 6490
rect 17972 6428 17973 6430
rect 17907 6427 17973 6428
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 15515 4996 15581 4997
rect 15515 4932 15516 4996
rect 15580 4932 15581 4996
rect 15515 4931 15581 4932
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14411 3500 14477 3501
rect 14411 3436 14412 3500
rect 14476 3436 14477 3500
rect 14411 3435 14477 3436
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14411 3228 14477 3229
rect 14411 3178 14412 3228
rect 14476 3178 14477 3228
rect 13859 2956 13925 2957
rect 13859 2892 13860 2956
rect 13924 2892 13925 2956
rect 13859 2891 13925 2892
rect 13862 2498 13922 2891
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 15518 1818 15578 4931
rect 17542 2957 17602 6342
rect 17723 6220 17789 6221
rect 17723 6156 17724 6220
rect 17788 6156 17789 6220
rect 17723 6155 17789 6156
rect 17726 5405 17786 6155
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 17723 5404 17789 5405
rect 17723 5340 17724 5404
rect 17788 5340 17789 5404
rect 17723 5339 17789 5340
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 20118 4453 20178 8875
rect 20854 6357 20914 20707
rect 20851 6356 20917 6357
rect 20851 6292 20852 6356
rect 20916 6292 20917 6356
rect 20851 6291 20917 6292
rect 20115 4452 20181 4453
rect 20115 4388 20116 4452
rect 20180 4388 20181 4452
rect 20115 4387 20181 4388
rect 21038 3909 21098 26419
rect 21219 25396 21285 25397
rect 21219 25332 21220 25396
rect 21284 25332 21285 25396
rect 21219 25331 21285 25332
rect 21222 20229 21282 25331
rect 21403 24036 21469 24037
rect 21403 23972 21404 24036
rect 21468 23972 21469 24036
rect 21403 23971 21469 23972
rect 21219 20228 21285 20229
rect 21219 20164 21220 20228
rect 21284 20164 21285 20228
rect 21219 20163 21285 20164
rect 21406 14650 21466 23971
rect 21771 23492 21837 23493
rect 21771 23428 21772 23492
rect 21836 23428 21837 23492
rect 21771 23427 21837 23428
rect 21774 19549 21834 23427
rect 21771 19548 21837 19549
rect 21771 19484 21772 19548
rect 21836 19484 21837 19548
rect 21771 19483 21837 19484
rect 21771 16556 21837 16557
rect 21771 16492 21772 16556
rect 21836 16492 21837 16556
rect 21771 16491 21837 16492
rect 21774 15330 21834 16491
rect 21958 16149 22018 26555
rect 23611 26348 23677 26349
rect 23611 26284 23612 26348
rect 23676 26284 23677 26348
rect 23611 26283 23677 26284
rect 22323 25940 22389 25941
rect 22323 25876 22324 25940
rect 22388 25876 22389 25940
rect 22323 25875 22389 25876
rect 22326 19821 22386 25875
rect 23427 24988 23493 24989
rect 23427 24924 23428 24988
rect 23492 24924 23493 24988
rect 23427 24923 23493 24924
rect 22323 19820 22389 19821
rect 22323 19756 22324 19820
rect 22388 19756 22389 19820
rect 22323 19755 22389 19756
rect 22323 18052 22389 18053
rect 22323 17988 22324 18052
rect 22388 17988 22389 18052
rect 22323 17987 22389 17988
rect 21955 16148 22021 16149
rect 21955 16084 21956 16148
rect 22020 16084 22021 16148
rect 21955 16083 22021 16084
rect 22139 15468 22205 15469
rect 22139 15404 22140 15468
rect 22204 15404 22205 15468
rect 22139 15403 22205 15404
rect 21955 15332 22021 15333
rect 21955 15330 21956 15332
rect 21774 15270 21956 15330
rect 21955 15268 21956 15270
rect 22020 15268 22021 15332
rect 21955 15267 22021 15268
rect 21406 14590 21834 14650
rect 21774 6901 21834 14590
rect 22142 11933 22202 15403
rect 22139 11932 22205 11933
rect 22139 11868 22140 11932
rect 22204 11868 22205 11932
rect 22139 11867 22205 11868
rect 22326 11661 22386 17987
rect 23059 17172 23060 17222
rect 23124 17172 23125 17222
rect 23059 17171 23125 17172
rect 23062 14789 23122 15182
rect 23059 14788 23125 14789
rect 23059 14724 23060 14788
rect 23124 14724 23125 14788
rect 23059 14723 23125 14724
rect 22694 12885 22754 13822
rect 22691 12884 22757 12885
rect 22691 12820 22692 12884
rect 22756 12820 22757 12884
rect 22691 12819 22757 12820
rect 22323 11660 22389 11661
rect 22323 11596 22324 11660
rect 22388 11596 22389 11660
rect 22323 11595 22389 11596
rect 21955 11388 22021 11389
rect 21955 11324 21956 11388
rect 22020 11324 22021 11388
rect 21955 11323 22021 11324
rect 21958 8397 22018 11323
rect 23430 9621 23490 24923
rect 23614 18053 23674 26283
rect 25454 26150 26066 26210
rect 25083 26076 25149 26077
rect 25083 26012 25084 26076
rect 25148 26012 25149 26076
rect 25083 26011 25149 26012
rect 23795 25124 23861 25125
rect 23795 25060 23796 25124
rect 23860 25060 23861 25124
rect 23795 25059 23861 25060
rect 23611 18052 23677 18053
rect 23611 17988 23612 18052
rect 23676 17988 23677 18052
rect 23798 18050 23858 25059
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 23979 22268 24045 22269
rect 23979 22204 23980 22268
rect 24044 22204 24045 22268
rect 23979 22203 24045 22204
rect 23982 21997 24042 22203
rect 23979 21996 24045 21997
rect 23979 21932 23980 21996
rect 24044 21932 24045 21996
rect 23979 21931 24045 21932
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 23979 21724 24045 21725
rect 23979 21660 23980 21724
rect 24044 21660 24045 21724
rect 23979 21659 24045 21660
rect 23982 20773 24042 21659
rect 23979 20772 24045 20773
rect 23979 20708 23980 20772
rect 24044 20708 24045 20772
rect 23979 20707 24045 20708
rect 23982 18733 24042 20707
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24899 19956 24965 19957
rect 24899 19892 24900 19956
rect 24964 19892 24965 19956
rect 24899 19891 24965 19892
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 23979 18732 24045 18733
rect 23979 18668 23980 18732
rect 24044 18668 24045 18732
rect 23979 18667 24045 18668
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 23798 17990 24042 18050
rect 23611 17987 23677 17988
rect 23611 14652 23677 14653
rect 23611 14588 23612 14652
rect 23676 14588 23677 14652
rect 23611 14587 23677 14588
rect 23614 12069 23674 14587
rect 23611 12068 23677 12069
rect 23611 12004 23612 12068
rect 23676 12004 23677 12068
rect 23611 12003 23677 12004
rect 23427 9620 23493 9621
rect 23427 9556 23428 9620
rect 23492 9556 23493 9620
rect 23427 9555 23493 9556
rect 23795 8804 23861 8805
rect 23795 8740 23796 8804
rect 23860 8740 23861 8804
rect 23795 8739 23861 8740
rect 21955 8396 22021 8397
rect 21955 8332 21956 8396
rect 22020 8332 22021 8396
rect 21955 8331 22021 8332
rect 21771 6900 21837 6901
rect 21771 6836 21772 6900
rect 21836 6836 21837 6900
rect 21771 6835 21837 6836
rect 21771 6356 21837 6357
rect 21771 6292 21772 6356
rect 21836 6292 21837 6356
rect 21771 6291 21837 6292
rect 23427 6356 23493 6357
rect 23427 6292 23428 6356
rect 23492 6292 23493 6356
rect 23427 6291 23493 6292
rect 21035 3908 21101 3909
rect 21035 3844 21036 3908
rect 21100 3844 21101 3908
rect 21035 3843 21101 3844
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 17539 2956 17605 2957
rect 17539 2892 17540 2956
rect 17604 2892 17605 2956
rect 17539 2891 17605 2892
rect 19610 2752 19930 3776
rect 21774 3773 21834 6291
rect 21771 3772 21837 3773
rect 21771 3708 21772 3772
rect 21836 3708 21837 3772
rect 21771 3707 21837 3708
rect 23430 3365 23490 6291
rect 23427 3364 23493 3365
rect 23427 3300 23428 3364
rect 23492 3300 23493 3364
rect 23427 3299 23493 3300
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 10915 1188 10981 1189
rect 10915 1124 10916 1188
rect 10980 1124 10981 1188
rect 10915 1123 10981 1124
rect 23798 237 23858 8739
rect 23982 5405 24042 17990
rect 24277 17440 24597 18464
rect 24715 18052 24781 18053
rect 24715 17988 24716 18052
rect 24780 17988 24781 18052
rect 24715 17987 24781 17988
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24718 13293 24778 17987
rect 24715 13292 24781 13293
rect 24715 13228 24716 13292
rect 24780 13228 24781 13292
rect 24715 13227 24781 13228
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24902 9621 24962 19891
rect 25086 10981 25146 26011
rect 25454 25618 25514 26150
rect 25819 25532 25885 25533
rect 25819 25468 25820 25532
rect 25884 25468 25885 25532
rect 25819 25467 25885 25468
rect 25267 21452 25333 21453
rect 25267 21388 25268 21452
rect 25332 21388 25333 21452
rect 25267 21387 25333 21388
rect 25270 13293 25330 21387
rect 25267 13292 25333 13293
rect 25267 13228 25268 13292
rect 25332 13228 25333 13292
rect 25267 13227 25333 13228
rect 25267 12884 25333 12885
rect 25267 12820 25268 12884
rect 25332 12820 25333 12884
rect 25267 12819 25333 12820
rect 25083 10980 25149 10981
rect 25083 10916 25084 10980
rect 25148 10916 25149 10980
rect 25083 10915 25149 10916
rect 24899 9620 24965 9621
rect 24899 9556 24900 9620
rect 24964 9556 24965 9620
rect 24899 9555 24965 9556
rect 25270 9485 25330 12819
rect 25454 9621 25514 21982
rect 25635 14788 25701 14789
rect 25635 14724 25636 14788
rect 25700 14724 25701 14788
rect 25635 14723 25701 14724
rect 25451 9620 25517 9621
rect 25451 9556 25452 9620
rect 25516 9556 25517 9620
rect 25451 9555 25517 9556
rect 25267 9484 25333 9485
rect 25267 9420 25268 9484
rect 25332 9420 25333 9484
rect 25267 9419 25333 9420
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 25638 8125 25698 14723
rect 25822 12341 25882 25467
rect 25819 12340 25885 12341
rect 25819 12276 25820 12340
rect 25884 12276 25885 12340
rect 25819 12275 25885 12276
rect 26006 9621 26066 26150
rect 26374 10981 26434 23342
rect 26371 10980 26437 10981
rect 26371 10916 26372 10980
rect 26436 10916 26437 10980
rect 26371 10915 26437 10916
rect 26003 9620 26069 9621
rect 26003 9556 26004 9620
rect 26068 9556 26069 9620
rect 26003 9555 26069 9556
rect 26742 9213 26802 19262
rect 26739 9212 26805 9213
rect 26739 9148 26740 9212
rect 26804 9148 26805 9212
rect 26739 9147 26805 9148
rect 25635 8124 25701 8125
rect 25635 8060 25636 8124
rect 25700 8060 25701 8124
rect 25635 8059 25701 8060
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24899 7036 24965 7037
rect 24899 6972 24900 7036
rect 24964 6972 24965 7036
rect 24899 6971 24965 6972
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 23979 5404 24045 5405
rect 23979 5340 23980 5404
rect 24044 5340 24045 5404
rect 23979 5339 24045 5340
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24902 2410 24962 6971
rect 24902 2350 25330 2410
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 24715 2004 24781 2005
rect 24715 1940 24716 2004
rect 24780 1940 24781 2004
rect 24715 1939 24781 1940
rect 24718 1818 24778 1939
rect 25270 1138 25330 2350
rect 23795 236 23861 237
rect 23795 172 23796 236
rect 23860 172 23861 236
rect 23795 171 23861 172
<< via4 >>
rect 1446 22662 1682 22898
rect 1998 10572 2234 10658
rect 1998 10508 2084 10572
rect 2084 10508 2148 10572
rect 2148 10508 2234 10572
rect 1998 10422 2234 10508
rect 2918 7852 3154 7938
rect 2918 7788 3004 7852
rect 3004 7788 3068 7852
rect 3068 7788 3154 7852
rect 2918 7702 3154 7788
rect 5310 25382 5546 25618
rect 6598 24702 6834 24938
rect 6046 21982 6282 22218
rect 5310 20622 5546 20858
rect 5126 16542 5362 16778
rect 4758 12462 4994 12698
rect 5126 8532 5362 8618
rect 5126 8468 5212 8532
rect 5212 8468 5276 8532
rect 5276 8468 5362 8532
rect 5126 8382 5362 8468
rect 5126 7022 5362 7258
rect 9726 21302 9962 21538
rect 7334 19262 7570 19498
rect 6966 11782 7202 12018
rect 7702 17902 7938 18138
rect 7702 9756 7938 9978
rect 7702 9742 7788 9756
rect 7788 9742 7852 9756
rect 7852 9742 7938 9756
rect 8070 6492 8306 6578
rect 8070 6428 8156 6492
rect 8156 6428 8220 6492
rect 8220 6428 8306 6492
rect 8070 6342 8306 6428
rect 11382 18804 11468 18818
rect 11468 18804 11532 18818
rect 11532 18804 11618 18818
rect 11382 18582 11618 18804
rect 11382 10422 11618 10658
rect 6046 3772 6282 3858
rect 9910 4452 10146 4538
rect 9910 4388 9996 4452
rect 9996 4388 10060 4452
rect 10060 4388 10146 4452
rect 9910 4302 10146 4388
rect 6046 3708 6132 3772
rect 6132 3708 6196 3772
rect 6196 3708 6282 3772
rect 6046 3622 6282 3708
rect 6598 3092 6834 3178
rect 6598 3028 6684 3092
rect 6684 3028 6748 3092
rect 6748 3028 6834 3092
rect 6598 2942 6834 3028
rect 5310 1582 5546 1818
rect 12854 20092 13090 20178
rect 12854 20028 12940 20092
rect 12940 20028 13004 20092
rect 13004 20028 13090 20092
rect 12854 19942 13090 20028
rect 15982 24852 16218 24938
rect 15982 24788 16068 24852
rect 16068 24788 16132 24852
rect 16132 24788 16218 24852
rect 15982 24702 16218 24788
rect 15430 23342 15666 23578
rect 13038 17372 13274 17458
rect 13038 17308 13124 17372
rect 13124 17308 13188 17372
rect 13188 17308 13274 17372
rect 13038 17222 13274 17308
rect 13774 16692 14010 16778
rect 13774 16628 13860 16692
rect 13860 16628 13924 16692
rect 13924 16628 14010 16692
rect 13774 16542 14010 16628
rect 14326 14502 14562 14738
rect 13590 13822 13826 14058
rect 13406 13156 13642 13378
rect 13406 13142 13492 13156
rect 13492 13142 13556 13156
rect 13556 13142 13642 13156
rect 14510 12462 14746 12698
rect 16718 17902 16954 18138
rect 16350 15182 16586 15418
rect 15798 12462 16034 12698
rect 20582 22662 20818 22898
rect 20214 21452 20450 21538
rect 20214 21388 20300 21452
rect 20300 21388 20364 21452
rect 20364 21388 20450 21452
rect 20214 21302 20450 21388
rect 20030 20772 20266 20858
rect 20030 20708 20116 20772
rect 20116 20708 20180 20772
rect 20180 20708 20266 20772
rect 20030 20622 20266 20708
rect 13590 3772 13826 3858
rect 13590 3708 13676 3772
rect 13676 3708 13740 3772
rect 13740 3708 13826 3772
rect 13590 3622 13826 3708
rect 16902 9742 17138 9978
rect 20214 14652 20450 14738
rect 20214 14588 20300 14652
rect 20300 14588 20364 14652
rect 20364 14588 20450 14652
rect 20214 14502 20450 14588
rect 20214 9742 20450 9978
rect 19294 8382 19530 8618
rect 17454 6342 17690 6578
rect 14326 3164 14412 3178
rect 14412 3164 14476 3178
rect 14476 3164 14562 3178
rect 14326 2942 14562 3164
rect 13774 2262 14010 2498
rect 20582 4452 20818 4538
rect 20582 4388 20668 4452
rect 20668 4388 20732 4452
rect 20732 4388 20818 4452
rect 20582 4302 20818 4388
rect 22606 20092 22842 20178
rect 22606 20028 22692 20092
rect 22692 20028 22756 20092
rect 22756 20028 22842 20092
rect 22606 19942 22842 20028
rect 22790 18732 23026 18818
rect 22790 18668 22876 18732
rect 22876 18668 22940 18732
rect 22940 18668 23026 18732
rect 22790 18582 23026 18668
rect 21318 11932 21554 12018
rect 21318 11868 21404 11932
rect 21404 11868 21468 11932
rect 21468 11868 21554 11932
rect 21318 11782 21554 11868
rect 22974 17236 23210 17458
rect 22974 17222 23060 17236
rect 23060 17222 23124 17236
rect 23124 17222 23210 17236
rect 22974 15182 23210 15418
rect 22606 13822 22842 14058
rect 22974 13292 23210 13378
rect 22974 13228 23060 13292
rect 23060 13228 23124 13292
rect 23124 13228 23210 13292
rect 22974 13142 23210 13228
rect 22606 2412 22842 2498
rect 22606 2348 22692 2412
rect 22692 2348 22756 2412
rect 22756 2348 22842 2412
rect 22606 2262 22842 2348
rect 13222 1582 13458 1818
rect 15430 1582 15666 1818
rect 4758 902 4994 1138
rect 25366 25382 25602 25618
rect 25366 21982 25602 22218
rect 26286 23342 26522 23578
rect 26654 19262 26890 19498
rect 24814 7852 25050 7938
rect 24814 7788 24900 7852
rect 24900 7788 24964 7852
rect 24964 7788 25050 7852
rect 24814 7702 25050 7788
rect 26102 7172 26338 7258
rect 26102 7108 26188 7172
rect 26188 7108 26252 7172
rect 26252 7108 26338 7172
rect 26102 7022 26338 7108
rect 24630 1582 24866 1818
rect 25182 902 25418 1138
<< metal5 >>
rect 5268 25618 25644 25660
rect 5268 25382 5310 25618
rect 5546 25382 25366 25618
rect 25602 25382 25644 25618
rect 5268 25340 25644 25382
rect 6556 24938 16260 24980
rect 6556 24702 6598 24938
rect 6834 24702 15982 24938
rect 16218 24702 16260 24938
rect 6556 24660 16260 24702
rect 15388 23578 26564 23620
rect 15388 23342 15430 23578
rect 15666 23342 26286 23578
rect 26522 23342 26564 23578
rect 15388 23300 26564 23342
rect 1404 22898 20860 22940
rect 1404 22662 1446 22898
rect 1682 22662 20582 22898
rect 20818 22662 20860 22898
rect 1404 22620 20860 22662
rect 6004 22218 25644 22260
rect 6004 21982 6046 22218
rect 6282 21982 25366 22218
rect 25602 21982 25644 22218
rect 6004 21940 25644 21982
rect 9684 21538 20492 21580
rect 9684 21302 9726 21538
rect 9962 21302 20214 21538
rect 20450 21302 20492 21538
rect 9684 21260 20492 21302
rect 5268 20858 20308 20900
rect 5268 20622 5310 20858
rect 5546 20622 20030 20858
rect 20266 20622 20308 20858
rect 5268 20580 20308 20622
rect 12812 20178 22884 20220
rect 12812 19942 12854 20178
rect 13090 19942 22606 20178
rect 22842 19942 22884 20178
rect 12812 19900 22884 19942
rect 7292 19498 26932 19540
rect 7292 19262 7334 19498
rect 7570 19262 26654 19498
rect 26890 19262 26932 19498
rect 7292 19220 26932 19262
rect 11340 18818 23068 18860
rect 11340 18582 11382 18818
rect 11618 18582 22790 18818
rect 23026 18582 23068 18818
rect 11340 18540 23068 18582
rect 7660 18138 16996 18180
rect 7660 17902 7702 18138
rect 7938 17902 16718 18138
rect 16954 17902 16996 18138
rect 7660 17860 16996 17902
rect 12996 17458 23252 17500
rect 12996 17222 13038 17458
rect 13274 17222 22974 17458
rect 23210 17222 23252 17458
rect 12996 17180 23252 17222
rect 5084 16778 14052 16820
rect 5084 16542 5126 16778
rect 5362 16542 13774 16778
rect 14010 16542 14052 16778
rect 5084 16500 14052 16542
rect 16308 15418 23252 15460
rect 16308 15182 16350 15418
rect 16586 15182 22974 15418
rect 23210 15182 23252 15418
rect 16308 15140 23252 15182
rect 14284 14738 20492 14780
rect 14284 14502 14326 14738
rect 14562 14502 20214 14738
rect 20450 14502 20492 14738
rect 14284 14460 20492 14502
rect 13548 14058 22884 14100
rect 13548 13822 13590 14058
rect 13826 13822 22606 14058
rect 22842 13822 22884 14058
rect 13548 13780 22884 13822
rect 13364 13378 23252 13420
rect 13364 13142 13406 13378
rect 13642 13142 22974 13378
rect 23210 13142 23252 13378
rect 13364 13100 23252 13142
rect 4716 12698 14788 12740
rect 4716 12462 4758 12698
rect 4994 12462 14510 12698
rect 14746 12462 14788 12698
rect 4716 12420 14788 12462
rect 15756 12698 16076 13100
rect 15756 12462 15798 12698
rect 16034 12462 16076 12698
rect 15756 12420 16076 12462
rect 6924 12018 21596 12060
rect 6924 11782 6966 12018
rect 7202 11782 21318 12018
rect 21554 11782 21596 12018
rect 6924 11740 21596 11782
rect 1956 10658 11660 10700
rect 1956 10422 1998 10658
rect 2234 10422 11382 10658
rect 11618 10422 11660 10658
rect 1956 10380 11660 10422
rect 7660 9978 20492 10020
rect 7660 9742 7702 9978
rect 7938 9742 16902 9978
rect 17138 9742 20214 9978
rect 20450 9742 20492 9978
rect 7660 9700 20492 9742
rect 5084 8618 19572 8660
rect 5084 8382 5126 8618
rect 5362 8382 19294 8618
rect 19530 8382 19572 8618
rect 5084 8340 19572 8382
rect 2876 7938 25092 7980
rect 2876 7702 2918 7938
rect 3154 7702 24814 7938
rect 25050 7702 25092 7938
rect 2876 7660 25092 7702
rect 5084 7258 26380 7300
rect 5084 7022 5126 7258
rect 5362 7022 26102 7258
rect 26338 7022 26380 7258
rect 5084 6980 26380 7022
rect 8028 6578 17732 6620
rect 8028 6342 8070 6578
rect 8306 6342 17454 6578
rect 17690 6342 17732 6578
rect 8028 6300 17732 6342
rect 9868 4538 20860 4580
rect 9868 4302 9910 4538
rect 10146 4302 20582 4538
rect 20818 4302 20860 4538
rect 9868 4260 20860 4302
rect 6004 3858 13868 3900
rect 6004 3622 6046 3858
rect 6282 3622 13590 3858
rect 13826 3622 13868 3858
rect 6004 3580 13868 3622
rect 6556 3178 14604 3220
rect 6556 2942 6598 3178
rect 6834 2942 14326 3178
rect 14562 2942 14604 3178
rect 6556 2900 14604 2942
rect 13732 2498 22884 2540
rect 13732 2262 13774 2498
rect 14010 2262 22606 2498
rect 22842 2262 22884 2498
rect 13732 2220 22884 2262
rect 5268 1818 13500 1860
rect 5268 1582 5310 1818
rect 5546 1582 13222 1818
rect 13458 1582 13500 1818
rect 5268 1540 13500 1582
rect 15388 1818 24908 1860
rect 15388 1582 15430 1818
rect 15666 1582 24630 1818
rect 24866 1582 24908 1818
rect 15388 1540 24908 1582
rect 4716 1138 25460 1180
rect 4716 902 4758 1138
rect 4994 902 25182 1138
rect 25418 902 25460 1138
rect 4716 860 25460 902
use scs8hd_fill_1  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_track_1.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_19
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l5_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_23
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_29
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A1
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4324 0 -1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A0
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_82
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_86
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_90
timestamp 1586364061
transform 1 0 9384 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_102
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_106
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_113
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _113_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_117
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_128
timestamp 1586364061
transform 1 0 12880 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_145
timestamp 1586364061
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_141
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_175
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_168
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_172
timestamp 1586364061
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_176
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_179
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_180
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_203
timestamp 1586364061
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _110_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_227
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_231
timestamp 1586364061
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_231
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_235
timestamp 1586364061
transform 1 0 22724 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 22908 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 22540 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _111_
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_239
timestamp 1586364061
transform 1 0 23092 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_243
timestamp 1586364061
transform 1 0 23460 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_239
timestamp 1586364061
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 23276 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 23644 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_254
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_258
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _108_
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_266
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_270
timestamp 1586364061
transform 1 0 25944 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 26128 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_274
timestamp 1586364061
transform 1 0 26312 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_buf_1  mux_bottom_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_10
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A0
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__S
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_46
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_70
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_74
timestamp 1586364061
transform 1 0 7912 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_78
timestamp 1586364061
transform 1 0 8280 0 -1 3808
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_buf_1  mux_bottom_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11684 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_110
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_114
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_134
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_138
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use scs8hd_conb_1  _047_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_158
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1586364061
transform 1 0 15824 0 -1 3808
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 17388 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_169
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_173
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_186
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_192
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_203
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_207
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_211
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 22264 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 23460 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 23828 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_241
timestamp 1586364061
transform 1 0 23276 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_245
timestamp 1586364061
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_258
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 25024 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_262
timestamp 1586364061
transform 1 0 25208 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25392 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_266
timestamp 1586364061
transform 1 0 25576 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25760 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_270
timestamp 1586364061
transform 1 0 25944 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 26128 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__S
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__S
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_17
timestamp 1586364061
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A1
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_21
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_81
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_85
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 314 592
use scs8hd_conb_1  _046_
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_103
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_109
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 13708 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_139
timestamp 1586364061
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_152
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_160
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_173
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1586364061
transform 1 0 21160 0 1 3808
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_210
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_214
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_227
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_231
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_234
timestamp 1586364061
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_238
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_254
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _096_
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 26128 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_266
timestamp 1586364061
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_270
timestamp 1586364061
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_274
timestamp 1586364061
transform 1 0 26312 0 1 3808
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A0
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__S
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__S
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6532 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_51
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_55
timestamp 1586364061
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_82
timestamp 1586364061
transform 1 0 8648 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_87
timestamp 1586364061
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_97
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 10212 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1586364061
transform 1 0 10396 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_115
timestamp 1586364061
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_128
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_132
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15456 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_158
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 15916 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_182
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_199
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_203
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_207
timestamp 1586364061
transform 1 0 20148 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_211
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_228
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 24472 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 24012 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_241
timestamp 1586364061
transform 1 0 23276 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_258
timestamp 1586364061
transform 1 0 24840 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25024 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_262
timestamp 1586364061
transform 1 0 25208 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 25392 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_266
timestamp 1586364061
transform 1 0 25576 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 25760 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_270
timestamp 1586364061
transform 1 0 25944 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 26128 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A1
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_19
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _048_
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_42
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_46
timestamp 1586364061
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_67
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _043_
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_80
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_84
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_94
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_115
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_119
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_136
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _114_
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_140
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_148
timestamp 1586364061
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_152
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_165
timestamp 1586364061
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_169
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_200
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_210
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_227
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_231
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_234
timestamp 1586364061
transform 1 0 22632 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_238
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 26128 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_266
timestamp 1586364061
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_270
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_274
timestamp 1586364061
transform 1 0 26312 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_8
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__S
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A0
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A1
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_25
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_21
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__S
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_36
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__S
timestamp 1586364061
transform 1 0 4600 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_2  _075_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_48
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_40
timestamp 1586364061
transform 1 0 4784 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__A0
timestamp 1586364061
transform 1 0 4968 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_56
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_52
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_59
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_55
timestamp 1586364061
transform 1 0 6164 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_69
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_65
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_60
timestamp 1586364061
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_conb_1  _049_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_6_86
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_82
timestamp 1586364061
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__A0
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__A1
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_96
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_92
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_90
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_112
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_118
timestamp 1586364061
transform 1 0 11960 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_127
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_120
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_122
timestamp 1586364061
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_158
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_153
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_149
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_162
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_167
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 16560 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_170
timestamp 1586364061
transform 1 0 16744 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_197
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_194
timestamp 1586364061
transform 1 0 18952 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _112_
timestamp 1586364061
transform 1 0 19320 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 866 592
use scs8hd_fill_1  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_214
timestamp 1586364061
transform 1 0 20792 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_210
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_227
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_228
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_234
timestamp 1586364061
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_231
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_238
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 24012 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_241
timestamp 1586364061
transform 1 0 23276 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_247
timestamp 1586364061
transform 1 0 23828 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_258
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_262
timestamp 1586364061
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_258
timestamp 1586364061
transform 1 0 24840 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25024 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_266
timestamp 1586364061
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_266
timestamp 1586364061
transform 1 0 25576 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25392 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_270
timestamp 1586364061
transform 1 0 25944 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_270
timestamp 1586364061
transform 1 0 25944 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 26128 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25760 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_274
timestamp 1586364061
transform 1 0 26312 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__S
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_11
timestamp 1586364061
transform 1 0 2116 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__A1
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6072 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 5888 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_46
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_50
timestamp 1586364061
transform 1 0 5704 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_63
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_81
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_85
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_90
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10396 0 -1 7072
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_120
timestamp 1586364061
transform 1 0 12144 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_137
timestamp 1586364061
transform 1 0 13708 0 -1 7072
box -38 -48 314 592
use scs8hd_buf_2  _115_
timestamp 1586364061
transform 1 0 15456 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_142
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_146
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_150
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 16560 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_160
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_164
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_187
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_191
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_208
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_228
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 24012 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 24748 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_241
timestamp 1586364061
transform 1 0 23276 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_247
timestamp 1586364061
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_253
timestamp 1586364061
transform 1 0 24380 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_259
timestamp 1586364061
transform 1 0 24932 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _101_
timestamp 1586364061
transform 1 0 25116 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_265
timestamp 1586364061
transform 1 0 25484 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 25668 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_269
timestamp 1586364061
transform 1 0 25852 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__A1
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_273
timestamp 1586364061
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__S
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_14
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_18
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__S
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__A0
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_48
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_52
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_56
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_78
timestamp 1586364061
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_82
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_97
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_101
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_149
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_166
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_170
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_200
timestamp 1586364061
transform 1 0 19504 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_210
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_214
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_227
timestamp 1586364061
transform 1 0 21988 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_231
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_234
timestamp 1586364061
transform 1 0 22632 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_238
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 406 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 24196 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_242
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_249
timestamp 1586364061
transform 1 0 24012 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_253
timestamp 1586364061
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 25300 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__A0
timestamp 1586364061
transform 1 0 25668 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 26036 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__A1
timestamp 1586364061
transform 1 0 26404 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_261
timestamp 1586364061
transform 1 0 25116 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_265
timestamp 1586364061
transform 1 0 25484 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_273
timestamp 1586364061
transform 1 0 26220 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__A0
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  FILLER_10_9
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_2  _074_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A1
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A0
timestamp 1586364061
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A1
timestamp 1586364061
transform 1 0 4968 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_40
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_70
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_74
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_90
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_98
timestamp 1586364061
transform 1 0 10120 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 10304 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_111
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_115
timestamp 1586364061
transform 1 0 11684 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_138
timestamp 1586364061
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_142
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_146
timestamp 1586364061
transform 1 0 14536 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_150
timestamp 1586364061
transform 1 0 14904 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17204 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_173
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_177
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _109_
timestamp 1586364061
transform 1 0 19320 0 -1 8160
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 17756 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 18768 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17572 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_194
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 22448 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_228
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 24012 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 23460 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__A0
timestamp 1586364061
transform 1 0 24564 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_241
timestamp 1586364061
transform 1 0 23276 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_245
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_253
timestamp 1586364061
transform 1 0 24380 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_257
timestamp 1586364061
transform 1 0 24748 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__A1
timestamp 1586364061
transform 1 0 24932 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _097_
timestamp 1586364061
transform 1 0 25116 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_265
timestamp 1586364061
transform 1 0 25484 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_269
timestamp 1586364061
transform 1 0 25852 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__A1
timestamp 1586364061
transform 1 0 26036 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_273
timestamp 1586364061
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1472 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A0
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__A1
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_13
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_17
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A0
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A1
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_30
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__S
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__S
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_47
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_60
timestamp 1586364061
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_95
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_108
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_116
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_120
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_128
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_151
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_172
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_176
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_203
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_207
timestamp 1586364061
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 22080 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 21528 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 21896 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_224
timestamp 1586364061
transform 1 0 21712 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24104 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_248
timestamp 1586364061
transform 1 0 23920 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_252
timestamp 1586364061
transform 1 0 24288 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_256
timestamp 1586364061
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_260
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_264
timestamp 1586364061
transform 1 0 25392 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__A0
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_268
timestamp 1586364061
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__A0
timestamp 1586364061
transform 1 0 25576 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_272
timestamp 1586364061
transform 1 0 26128 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 25944 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_276
timestamp 1586364061
transform 1 0 26496 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 26312 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_conb_1  _041_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__S
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__S
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__A1
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__A0
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_45
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_49
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_53
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_57
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_77
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_81
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_85
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_90
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_96
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_132
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_173
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_177
timestamp 1586364061
transform 1 0 17388 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 18768 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19136 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_198
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19504 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 22264 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22908 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_228
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_235
timestamp 1586364061
transform 1 0 22724 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23460 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 23276 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 23920 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 24288 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 24656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_246
timestamp 1586364061
transform 1 0 23736 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_250
timestamp 1586364061
transform 1 0 24104 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_254
timestamp 1586364061
transform 1 0 24472 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_258
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25024 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_262
timestamp 1586364061
transform 1 0 25208 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25392 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_266
timestamp 1586364061
transform 1 0 25576 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25760 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_270
timestamp 1586364061
transform 1 0 25944 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 26128 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 3312 0 1 9248
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_20
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_47
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_43
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_50
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_56
timestamp 1586364061
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_52
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_69
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_63
timestamp 1586364061
transform 1 0 6900 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_67
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_60
timestamp 1586364061
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_87
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_84
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_80
timestamp 1586364061
transform 1 0 8464 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_14_109
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_107
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1586364061
transform 1 0 10304 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_113
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_115
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_111
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_13_119
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_126
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_126
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_conb_1  _045_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_131
timestamp 1586364061
transform 1 0 13156 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_130
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_14_147
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_143
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_151
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_157
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_153
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_169
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_180
timestamp 1586364061
transform 1 0 17664 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_197
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_207
timestamp 1586364061
transform 1 0 20148 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_203
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_211
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_214
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_210
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_228
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_227
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_231
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 22264 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 22540 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _039_
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_235
timestamp 1586364061
transform 1 0 22724 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_235
timestamp 1586364061
transform 1 0 22724 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 22908 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 22908 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_239
timestamp 1586364061
transform 1 0 23092 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 23276 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_243
timestamp 1586364061
transform 1 0 23460 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_buf_1  mux_right_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23552 0 -1 10336
box -38 -48 314 592
use scs8hd_buf_1  mux_right_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_248
timestamp 1586364061
transform 1 0 23920 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24012 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_252
timestamp 1586364061
transform 1 0 24288 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 24380 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24104 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24564 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  mux_right_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24564 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_262
timestamp 1586364061
transform 1 0 25208 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_258
timestamp 1586364061
transform 1 0 24840 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_261
timestamp 1586364061
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25024 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_266
timestamp 1586364061
transform 1 0 25576 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_265
timestamp 1586364061
transform 1 0 25484 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 25392 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 25300 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_270
timestamp 1586364061
transform 1 0 25944 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 25760 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 26036 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_274
timestamp 1586364061
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_273
timestamp 1586364061
transform 1 0 26220 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_buf_2  _070_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 1786 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_35
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_76
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_80
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_94
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use scs8hd_conb_1  _044_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12972 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13340 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_126
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_131
timestamp 1586364061
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_15_158
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_162
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_210
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_214
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 22908 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_227
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_231
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_235
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _095_
timestamp 1586364061
transform 1 0 24564 0 1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 23276 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23828 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_239
timestamp 1586364061
transform 1 0 23092 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_243
timestamp 1586364061
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_249
timestamp 1586364061
transform 1 0 24012 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_259
timestamp 1586364061
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_267 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25668 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_275
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _037_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_55
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_59
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_81
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_87
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_97
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_120
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_124
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_128
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_138
timestamp 1586364061
transform 1 0 13800 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_142
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_146
timestamp 1586364061
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_150
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_157
timestamp 1586364061
transform 1 0 15548 0 -1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 16192 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_162
timestamp 1586364061
transform 1 0 16008 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18952 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 18768 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_203
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_207
timestamp 1586364061
transform 1 0 20148 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 22448 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_228
timestamp 1586364061
transform 1 0 22080 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _094_
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 23644 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24012 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 24380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_241
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_247
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 25116 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25484 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_259
timestamp 1586364061
transform 1 0 24932 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_267
timestamp 1586364061
transform 1 0 25668 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_14
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_18
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _073_
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_41
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_45
timestamp 1586364061
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_81
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_85
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_89
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_119
timestamp 1586364061
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12972 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_148
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_152
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_203
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_207
timestamp 1586364061
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_211
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_216
timestamp 1586364061
transform 1 0 20976 0 1 11424
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_221
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_234
timestamp 1586364061
transform 1 0 22632 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_238
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_261
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_258
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _093_
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_266
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_270
timestamp 1586364061
transform 1 0 25944 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 26128 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_274
timestamp 1586364061
transform 1 0 26312 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_conb_1  _036_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_12
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _072_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__A0
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_40
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__A0
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_60
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_73
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_77
timestamp 1586364061
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use scs8hd_conb_1  _042_
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9936 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_98
timestamp 1586364061
transform 1 0 10120 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10304 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_109
timestamp 1586364061
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_136
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_140
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_148
timestamp 1586364061
transform 1 0 14720 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_144
timestamp 1586364061
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_158
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1586364061
transform 1 0 16192 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 16008 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_173
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_177
timestamp 1586364061
transform 1 0 17388 0 -1 12512
box -38 -48 130 592
use scs8hd_conb_1  _040_
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_180
timestamp 1586364061
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_187
timestamp 1586364061
transform 1 0 18308 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_191
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_204
timestamp 1586364061
transform 1 0 19872 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1586364061
transform 1 0 21804 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 21344 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 22816 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_219
timestamp 1586364061
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_222
timestamp 1586364061
transform 1 0 21528 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_234
timestamp 1586364061
transform 1 0 22632 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_238
timestamp 1586364061
transform 1 0 23000 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23368 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 24380 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 23184 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 24748 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_255
timestamp 1586364061
transform 1 0 24564 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _092_
timestamp 1586364061
transform 1 0 24932 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25484 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_267
timestamp 1586364061
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__S
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__S
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_17
timestamp 1586364061
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_29
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_25
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_21
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__A1
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_36
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_49
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_53
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8280 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_76
timestamp 1586364061
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_92
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_109
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_105
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_116
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_112
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_119
timestamp 1586364061
transform 1 0 12052 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_123
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_136
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 13800 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_148
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_144
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_140
timestamp 1586364061
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_142
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_158
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_155
timestamp 1586364061
transform 1 0 15364 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_160
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 15732 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 15916 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_174
timestamp 1586364061
transform 1 0 17112 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_170
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_177
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17296 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 16928 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17480 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 18308 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_191
timestamp 1586364061
transform 1 0 18676 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_189
timestamp 1586364061
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_212
timestamp 1586364061
transform 1 0 20608 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_204
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_208
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 22816 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_229
timestamp 1586364061
transform 1 0 22172 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_233
timestamp 1586364061
transform 1 0 22540 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_234
timestamp 1586364061
transform 1 0 22632 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_238
timestamp 1586364061
transform 1 0 23000 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 23184 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_255
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_254
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 24748 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 24380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_261
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_258
timestamp 1586364061
transform 1 0 24840 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _090_
timestamp 1586364061
transform 1 0 25208 0 1 12512
box -38 -48 406 592
use scs8hd_buf_2  _089_
timestamp 1586364061
transform 1 0 24932 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_271
timestamp 1586364061
transform 1 0 26036 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_267
timestamp 1586364061
transform 1 0 25668 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_270 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25944 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_266
timestamp 1586364061
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25852 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25484 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_276
timestamp 1586364061
transform 1 0 26496 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_14
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_18
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_22
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_34
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_38
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_55
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 6992 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_83
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_87
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_91
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_120
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_136
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_149
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_153
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_170
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_174
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_178
timestamp 1586364061
transform 1 0 17480 0 1 13600
box -38 -48 314 592
use scs8hd_conb_1  _032_
timestamp 1586364061
transform 1 0 18400 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 18216 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_191
timestamp 1586364061
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_195
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_21_218
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1586364061
transform 1 0 21896 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 21712 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 22908 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_222
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_235
timestamp 1586364061
transform 1 0 22724 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_239
timestamp 1586364061
transform 1 0 23092 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_254
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 314 592
use scs8hd_buf_2  _088_
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 26128 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_259
timestamp 1586364061
transform 1 0 24932 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_266
timestamp 1586364061
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_270
timestamp 1586364061
transform 1 0 25944 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_274
timestamp 1586364061
transform 1 0 26312 0 1 13600
box -38 -48 314 592
use scs8hd_buf_1  mux_left_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_53
timestamp 1586364061
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_57
timestamp 1586364061
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_2  _071_
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_65
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_69
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 11960 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 11776 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_112
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_137
timestamp 1586364061
transform 1 0 13708 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14260 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 13892 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_157
timestamp 1586364061
transform 1 0 15548 0 -1 14688
box -38 -48 406 592
use scs8hd_conb_1  _038_
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16468 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 15916 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_186
timestamp 1586364061
transform 1 0 18216 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_194
timestamp 1586364061
transform 1 0 18952 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_1  mux_top_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_210
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_218
timestamp 1586364061
transform 1 0 21160 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 22264 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 21344 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 21896 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_222
timestamp 1586364061
transform 1 0 21528 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_228
timestamp 1586364061
transform 1 0 22080 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1586364061
transform 1 0 24748 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 24564 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_249
timestamp 1586364061
transform 1 0 24012 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_253
timestamp 1586364061
transform 1 0 24380 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25760 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 26128 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_266
timestamp 1586364061
transform 1 0 25576 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_270
timestamp 1586364061
transform 1 0 25944 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_274
timestamp 1586364061
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_1  mux_left_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_6
timestamp 1586364061
transform 1 0 1656 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_10
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_23
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_50
timestamp 1586364061
transform 1 0 5704 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_54
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_58
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1586364061
transform 1 0 6992 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 1786 592
use scs8hd_conb_1  _050_
timestamp 1586364061
transform 1 0 11040 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_100
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_104
timestamp 1586364061
transform 1 0 10672 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_111
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_115
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_119
timestamp 1586364061
transform 1 0 12052 0 1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 1786 592
use scs8hd_buf_1  mux_top_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_139
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_146
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_152
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19964 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19780 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_201
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _091_
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 22264 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_224
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_228
timestamp 1586364061
transform 1 0 22080 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_236
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_240
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_254
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_261
timestamp 1586364061
transform 1 0 25116 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_258
timestamp 1586364061
transform 1 0 24840 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _086_
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_266
timestamp 1586364061
transform 1 0 25576 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_270
timestamp 1586364061
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 26128 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_274
timestamp 1586364061
transform 1 0 26312 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_buf_1  mux_left_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_6
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_12
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4692 0 -1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4508 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_58
timestamp 1586364061
transform 1 0 6440 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 6624 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_62
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_66
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_70
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_74
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _062_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_97
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10580 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_101
timestamp 1586364061
transform 1 0 10396 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_124
timestamp 1586364061
transform 1 0 12512 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_128
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_149
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_158
timestamp 1586364061
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 15456 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 15732 0 -1 15776
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18216 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 17664 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 19228 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_182
timestamp 1586364061
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_195
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use scs8hd_conb_1  _035_
timestamp 1586364061
transform 1 0 19780 0 -1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 19596 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_199
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_210
timestamp 1586364061
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 22448 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 22264 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_224
timestamp 1586364061
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_228
timestamp 1586364061
transform 1 0 22080 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 24380 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 24748 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_255
timestamp 1586364061
transform 1 0 24564 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_2  _084_
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 25484 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_267
timestamp 1586364061
transform 1 0 25668 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2024 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_19
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 3036 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_23
timestamp 1586364061
transform 1 0 3220 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_36
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_40
timestamp 1586364061
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_81
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_85
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_89
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _028_
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11040 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_102
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_106
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_136
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_149
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_153
timestamp 1586364061
transform 1 0 15180 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_162
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _029_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_187
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_191
timestamp 1586364061
transform 1 0 18676 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_214
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21620 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 22724 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_219
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_237
timestamp 1586364061
transform 1 0 22908 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23092 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_241
timestamp 1586364061
transform 1 0 23276 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_254
timestamp 1586364061
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use scs8hd_buf_2  _085_
timestamp 1586364061
transform 1 0 25208 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 26128 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_258
timestamp 1586364061
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_266
timestamp 1586364061
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_270
timestamp 1586364061
transform 1 0 25944 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_274
timestamp 1586364061
transform 1 0 26312 0 1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_26_6
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_1  mux_left_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_12
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_27_29
timestamp 1586364061
transform 1 0 3772 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_36
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_33
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_40
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use scs8hd_fill_1  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_55
timestamp 1586364061
transform 1 0 6164 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_51
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6348 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6440 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 6532 0 -1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_66
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_60
timestamp 1586364061
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_buf_2  _068_
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_70
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_78
timestamp 1586364061
transform 1 0 8280 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1586364061
transform 1 0 8280 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_87
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_86
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_82
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_91
timestamp 1586364061
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_97
timestamp 1586364061
transform 1 0 10028 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10304 0 -1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_119
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_125
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_136
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_146
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_142
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_148
timestamp 1586364061
transform 1 0 14720 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_144
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_140
timestamp 1586364061
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14536 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_151
timestamp 1586364061
transform 1 0 14996 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _033_
timestamp 1586364061
transform 1 0 15364 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 15456 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_158
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15640 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_162
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_171
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17020 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1586364061
transform 1 0 17204 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_188
timestamp 1586364061
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_184
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_197
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_192
timestamp 1586364061
transform 1 0 18768 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 19044 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_206
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_210
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_225
timestamp 1586364061
transform 1 0 21804 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_26_228
timestamp 1586364061
transform 1 0 22080 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 21896 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_236
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_229
timestamp 1586364061
transform 1 0 22172 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_234
timestamp 1586364061
transform 1 0 22632 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 22448 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 22264 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _087_
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22724 0 -1 16864
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 24656 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_254
timestamp 1586364061
transform 1 0 24472 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_254
timestamp 1586364061
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_258
timestamp 1586364061
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_258
timestamp 1586364061
transform 1 0 24840 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _083_
timestamp 1586364061
transform 1 0 25208 0 -1 16864
box -38 -48 406 592
use scs8hd_buf_2  _082_
timestamp 1586364061
transform 1 0 25208 0 1 16864
box -38 -48 406 592
use scs8hd_decap_6  FILLER_27_270
timestamp 1586364061
transform 1 0 25944 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_266
timestamp 1586364061
transform 1 0 25576 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_270
timestamp 1586364061
transform 1 0 25944 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_266
timestamp 1586364061
transform 1 0 25576 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 25760 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 25760 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_274
timestamp 1586364061
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_1  mux_left_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_6
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_10
timestamp 1586364061
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 4324 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_37
timestamp 1586364061
transform 1 0 4508 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_50
timestamp 1586364061
transform 1 0 5704 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_54
timestamp 1586364061
transform 1 0 6072 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_67
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_73
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11132 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 11500 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11960 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_107
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_111
timestamp 1586364061
transform 1 0 11316 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_115
timestamp 1586364061
transform 1 0 11684 0 -1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12144 0 -1 17952
box -38 -48 866 592
use scs8hd_buf_1  mux_top_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13708 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 13340 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 14168 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_140
timestamp 1586364061
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_144
timestamp 1586364061
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_148
timestamp 1586364061
transform 1 0 14720 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17204 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_173
timestamp 1586364061
transform 1 0 17020 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_177
timestamp 1586364061
transform 1 0 17388 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 17756 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17572 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19136 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__A1
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_194
timestamp 1586364061
transform 1 0 18952 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_198
timestamp 1586364061
transform 1 0 19320 0 -1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use scs8hd_buf_1  mux_right_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19780 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 19596 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__A0
timestamp 1586364061
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_210
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 22724 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 22448 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_228
timestamp 1586364061
transform 1 0 22080 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_234
timestamp 1586364061
transform 1 0 22632 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 24656 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_254
timestamp 1586364061
transform 1 0 24472 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_2  _081_
timestamp 1586364061
transform 1 0 25208 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 25024 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_258
timestamp 1586364061
transform 1 0 24840 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_266
timestamp 1586364061
transform 1 0 25576 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_274
timestamp 1586364061
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 1786 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_28
timestamp 1586364061
transform 1 0 3680 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_67
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_80
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_84
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_97
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _031_
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_143
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_148
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17020 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_188
timestamp 1586364061
transform 1 0 18400 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_buf_1  mux_right_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18124 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_192
timestamp 1586364061
transform 1 0 18768 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18584 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18952 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_215
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 21620 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 22632 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_219
timestamp 1586364061
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_236
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_254
timestamp 1586364061
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use scs8hd_buf_2  _080_
timestamp 1586364061
transform 1 0 25208 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_258
timestamp 1586364061
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_266
timestamp 1586364061
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_270
timestamp 1586364061
transform 1 0 25944 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_276
timestamp 1586364061
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use scs8hd_buf_1  mux_left_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_11
timestamp 1586364061
transform 1 0 2116 0 -1 19040
box -38 -48 314 592
use scs8hd_buf_2  _069_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__S
timestamp 1586364061
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_40
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_65
timestamp 1586364061
transform 1 0 7084 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_71
timestamp 1586364061
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use scs8hd_buf_2  _064_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10212 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_88
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_97
timestamp 1586364061
transform 1 0 10028 0 -1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 10580 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_101
timestamp 1586364061
transform 1 0 10396 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1586364061
transform 1 0 13340 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_124
timestamp 1586364061
transform 1 0 12512 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_128
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 314 592
use scs8hd_buf_1  mux_top_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 14352 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 14720 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_142
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_146
timestamp 1586364061
transform 1 0 14536 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_150
timestamp 1586364061
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_157
timestamp 1586364061
transform 1 0 15548 0 -1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 15732 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_161
timestamp 1586364061
transform 1 0 15916 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_165
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 18676 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_185
timestamp 1586364061
transform 1 0 18124 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_189
timestamp 1586364061
transform 1 0 18492 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_210
timestamp 1586364061
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 22448 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_229
timestamp 1586364061
transform 1 0 22172 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 24380 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 24748 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_255
timestamp 1586364061
transform 1 0 24564 0 -1 19040
box -38 -48 222 592
use scs8hd_buf_2  _079_
timestamp 1586364061
transform 1 0 24932 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 1786 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 3680 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_26
timestamp 1586364061
transform 1 0 3496 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_30
timestamp 1586364061
transform 1 0 3864 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_buf_2  _065_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 7360 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_66
timestamp 1586364061
transform 1 0 7176 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_70
timestamp 1586364061
transform 1 0 7544 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_94
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1586364061
transform 1 0 13156 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12696 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_128
timestamp 1586364061
transform 1 0 12880 0 1 19040
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 15088 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 14904 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_140
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_144
timestamp 1586364061
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_148
timestamp 1586364061
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  mux_right_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A0
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__S
timestamp 1586364061
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_161
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_165
timestamp 1586364061
transform 1 0 16284 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_169
timestamp 1586364061
transform 1 0 16652 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18676 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A1
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 18492 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_188
timestamp 1586364061
transform 1 0 18400 0 1 19040
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20056 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 19688 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_200
timestamp 1586364061
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_204
timestamp 1586364061
transform 1 0 19872 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_217
timestamp 1586364061
transform 1 0 21068 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21252 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21620 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_221
timestamp 1586364061
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_225
timestamp 1586364061
transform 1 0 21804 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_236
timestamp 1586364061
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_240
timestamp 1586364061
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_254
timestamp 1586364061
transform 1 0 24472 0 1 19040
box -38 -48 406 592
use scs8hd_buf_2  _078_
timestamp 1586364061
transform 1 0 25208 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 24932 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_258
timestamp 1586364061
transform 1 0 24840 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_261
timestamp 1586364061
transform 1 0 25116 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_266
timestamp 1586364061
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_270
timestamp 1586364061
transform 1 0 25944 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_276
timestamp 1586364061
transform 1 0 26496 0 1 19040
box -38 -48 130 592
use scs8hd_conb_1  _053_
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__A0
timestamp 1586364061
transform 1 0 1932 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_11
timestamp 1586364061
transform 1 0 2116 0 -1 20128
box -38 -48 314 592
use scs8hd_buf_2  _067_
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 4600 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_36
timestamp 1586364061
transform 1 0 4416 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__S
timestamp 1586364061
transform 1 0 4968 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_40
timestamp 1586364061
transform 1 0 4784 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7912 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_66
timestamp 1586364061
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_70
timestamp 1586364061
transform 1 0 7544 0 -1 20128
box -38 -48 222 592
use scs8hd_conb_1  _051_
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 10212 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_83
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_96
timestamp 1586364061
transform 1 0 9936 0 -1 20128
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12052 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11684 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_101
timestamp 1586364061
transform 1 0 10396 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_113
timestamp 1586364061
transform 1 0 11500 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_121
timestamp 1586364061
transform 1 0 12236 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_125
timestamp 1586364061
transform 1 0 12604 0 -1 20128
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1586364061
transform 1 0 17020 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A0
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16836 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_163
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_168
timestamp 1586364061
transform 1 0 16560 0 -1 20128
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 18400 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__A1
timestamp 1586364061
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_182
timestamp 1586364061
transform 1 0 17848 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_186
timestamp 1586364061
transform 1 0 18216 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20240 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 19596 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_199
timestamp 1586364061
transform 1 0 19412 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_203
timestamp 1586364061
transform 1 0 19780 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_207
timestamp 1586364061
transform 1 0 20148 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_210
timestamp 1586364061
transform 1 0 20424 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 22816 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_234
timestamp 1586364061
transform 1 0 22632 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_238
timestamp 1586364061
transform 1 0 23000 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1586364061
transform 1 0 23368 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 24380 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 24748 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 23184 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_255
timestamp 1586364061
transform 1 0 24564 0 -1 20128
box -38 -48 222 592
use scs8hd_buf_2  _077_
timestamp 1586364061
transform 1 0 24932 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__A1
timestamp 1586364061
transform 1 0 1748 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__A1
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1586364061
transform 1 0 1932 0 -1 21216
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_4_
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_18
timestamp 1586364061
transform 1 0 2760 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_18
timestamp 1586364061
transform 1 0 2760 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A1
timestamp 1586364061
transform 1 0 2944 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__S
timestamp 1586364061
transform 1 0 2944 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_22
timestamp 1586364061
transform 1 0 3128 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_22
timestamp 1586364061
transform 1 0 3128 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A0
timestamp 1586364061
transform 1 0 3312 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_26
timestamp 1586364061
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 3680 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 3864 0 1 20128
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_34_45
timestamp 1586364061
transform 1 0 5244 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_41
timestamp 1586364061
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_49
timestamp 1586364061
transform 1 0 5612 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 5428 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 5060 0 -1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1586364061
transform 1 0 5612 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_58
timestamp 1586364061
transform 1 0 6440 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_62
timestamp 1586364061
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_68
timestamp 1586364061
transform 1 0 7360 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6624 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7176 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6992 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7176 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_79
timestamp 1586364061
transform 1 0 8372 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_75
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8188 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7544 0 1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7728 0 1 20128
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_34_87
timestamp 1586364061
transform 1 0 9108 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_83
timestamp 1586364061
transform 1 0 8740 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 8924 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_91
timestamp 1586364061
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_95
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_91
timestamp 1586364061
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1586364061
transform 1 0 10212 0 1 20128
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9752 0 -1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__A0
timestamp 1586364061
transform 1 0 11684 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_108
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_112
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_113
timestamp 1586364061
transform 1 0 11500 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12236 0 -1 21216
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_137
timestamp 1586364061
transform 1 0 13708 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_134
timestamp 1586364061
transform 1 0 13432 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_130
timestamp 1586364061
transform 1 0 13064 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_136
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_132
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 13524 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 13892 0 -1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 866 592
use scs8hd_buf_2  _133_
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_149
timestamp 1586364061
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_156
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_153
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_149
timestamp 1586364061
transform 1 0 14812 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__A1
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_168
timestamp 1586364061
transform 1 0 16560 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_163
timestamp 1586364061
transform 1 0 16100 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_33_160
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__S
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A1
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1586364061
transform 1 0 16376 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_176
timestamp 1586364061
transform 1 0 17296 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_172
timestamp 1586364061
transform 1 0 16928 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_175
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 16744 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__A0
timestamp 1586364061
transform 1 0 17112 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__A0
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_187
timestamp 1586364061
transform 1 0 18308 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_182
timestamp 1586364061
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__S
timestamp 1586364061
transform 1 0 17664 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1586364061
transform 1 0 17664 0 -1 21216
box -38 -48 866 592
use scs8hd_conb_1  _034_
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_193
timestamp 1586364061
transform 1 0 18860 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_189
timestamp 1586364061
transform 1 0 18492 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_191
timestamp 1586364061
transform 1 0 18676 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 18676 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__S
timestamp 1586364061
transform 1 0 18492 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19044 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1586364061
transform 1 0 19228 0 -1 21216
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_34_206
timestamp 1586364061
transform 1 0 20056 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20240 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_210
timestamp 1586364061
transform 1 0 20424 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_214
timestamp 1586364061
transform 1 0 20792 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_218
timestamp 1586364061
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20976 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 21068 0 -1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 21712 0 -1 21216
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1586364061
transform 1 0 21528 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 22540 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 21528 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 22908 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_231
timestamp 1586364061
transform 1 0 22356 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_235
timestamp 1586364061
transform 1 0 22724 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_219
timestamp 1586364061
transform 1 0 21252 0 -1 21216
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23644 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 24012 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_239
timestamp 1586364061
transform 1 0 23092 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_243
timestamp 1586364061
transform 1 0 23460 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_247
timestamp 1586364061
transform 1 0 23828 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_264
timestamp 1586364061
transform 1 0 25392 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_260
timestamp 1586364061
transform 1 0 25024 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_264
timestamp 1586364061
transform 1 0 25392 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25208 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 25576 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_272
timestamp 1586364061
transform 1 0 26128 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_33_272
timestamp 1586364061
transform 1 0 26128 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_268
timestamp 1586364061
transform 1 0 25760 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 25944 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_276
timestamp 1586364061
transform 1 0 26496 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_6_
timestamp 1586364061
transform 1 0 1840 0 1 21216
box -38 -48 866 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__A1
timestamp 1586364061
transform 1 0 1656 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__A0
timestamp 1586364061
transform 1 0 2852 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_17
timestamp 1586364061
transform 1 0 2668 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1586364061
transform 1 0 3404 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 3220 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_21
timestamp 1586364061
transform 1 0 3036 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_34
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_38
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6440 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 6072 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7452 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 6992 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_60
timestamp 1586364061
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_66
timestamp 1586364061
transform 1 0 7176 0 1 21216
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_90
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_95
timestamp 1586364061
transform 1 0 9844 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11500 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11868 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_107
timestamp 1586364061
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_111
timestamp 1586364061
transform 1 0 11316 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_115
timestamp 1586364061
transform 1 0 11684 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_119
timestamp 1586364061
transform 1 0 12052 0 1 21216
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 13064 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 12696 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_128
timestamp 1586364061
transform 1 0 12880 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 15272 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_151
timestamp 1586364061
transform 1 0 14996 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__S
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_160
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 18584 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 18400 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_209
timestamp 1586364061
transform 1 0 20332 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_213
timestamp 1586364061
transform 1 0 20700 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 22632 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22080 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_226
timestamp 1586364061
transform 1 0 21896 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_236
timestamp 1586364061
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_240
timestamp 1586364061
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_254
timestamp 1586364061
transform 1 0 24472 0 1 21216
box -38 -48 222 592
use scs8hd_buf_2  _076_
timestamp 1586364061
transform 1 0 25208 0 1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 25760 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_258
timestamp 1586364061
transform 1 0 24840 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_266
timestamp 1586364061
transform 1 0 25576 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_270
timestamp 1586364061
transform 1 0 25944 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_276
timestamp 1586364061
transform 1 0 26496 0 1 21216
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1586364061
transform 1 0 1840 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2852 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__A0
timestamp 1586364061
transform 1 0 1656 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_17
timestamp 1586364061
transform 1 0 2668 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 4232 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_21
timestamp 1586364061
transform 1 0 3036 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1586364061
transform 1 0 6440 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5428 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5888 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_45
timestamp 1586364061
transform 1 0 5244 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_49
timestamp 1586364061
transform 1 0 5612 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_54
timestamp 1586364061
transform 1 0 6072 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_67
timestamp 1586364061
transform 1 0 7268 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_73
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_2  _056_
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10212 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_88
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_97
timestamp 1586364061
transform 1 0 10028 0 -1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_101
timestamp 1586364061
transform 1 0 10396 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1586364061
transform 1 0 13524 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 13248 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_127
timestamp 1586364061
transform 1 0 12788 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_131
timestamp 1586364061
transform 1 0 13156 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_134
timestamp 1586364061
transform 1 0 13432 0 -1 22304
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14536 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14904 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_144
timestamp 1586364061
transform 1 0 14352 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_148
timestamp 1586364061
transform 1 0 14720 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_152
timestamp 1586364061
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17204 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_173
timestamp 1586364061
transform 1 0 17020 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_177
timestamp 1586364061
transform 1 0 17388 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1586364061
transform 1 0 18124 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 19136 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 17940 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 17572 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_181
timestamp 1586364061
transform 1 0 17756 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_194
timestamp 1586364061
transform 1 0 18952 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_198
timestamp 1586364061
transform 1 0 19320 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_2  _125_
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21068 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20240 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 19504 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_206
timestamp 1586364061
transform 1 0 20056 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_210
timestamp 1586364061
transform 1 0 20424 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 22632 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22080 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 22448 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_226
timestamp 1586364061
transform 1 0 21896 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_230
timestamp 1586364061
transform 1 0 22264 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23644 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24012 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_243
timestamp 1586364061
transform 1 0 23460 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_247
timestamp 1586364061
transform 1 0 23828 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_260
timestamp 1586364061
transform 1 0 25024 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_36_272
timestamp 1586364061
transform 1 0 26128 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_2  _066_
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2668 0 1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_11
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4232 0 1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 3680 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 4048 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_26
timestamp 1586364061
transform 1 0 3496 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_30
timestamp 1586364061
transform 1 0 3864 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 8096 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_78
timestamp 1586364061
transform 1 0 8280 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 8648 0 1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 8464 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _135_
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 11040 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 10672 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_101
timestamp 1586364061
transform 1 0 10396 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_106
timestamp 1586364061
transform 1 0 10856 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_114
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_118
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_132
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_136
timestamp 1586364061
transform 1 0 13616 0 1 22304
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14076 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_140
timestamp 1586364061
transform 1 0 13984 0 1 22304
box -38 -48 130 592
use scs8hd_buf_2  _129_
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 16560 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_162
timestamp 1586364061
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_166
timestamp 1586364061
transform 1 0 16376 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_170
timestamp 1586364061
transform 1 0 16744 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_175
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_179
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_193
timestamp 1586364061
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_197
timestamp 1586364061
transform 1 0 19228 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1586364061
transform 1 0 21160 0 1 22304
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1586364061
transform 1 0 19596 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 20976 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_210
timestamp 1586364061
transform 1 0 20424 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_214
timestamp 1586364061
transform 1 0 20792 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_227
timestamp 1586364061
transform 1 0 21988 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_231
timestamp 1586364061
transform 1 0 22356 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_234
timestamp 1586364061
transform 1 0 22632 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_238
timestamp 1586364061
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use scs8hd_conb_1  _030_
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 314 592
use scs8hd_buf_2  _120_
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 24196 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_242
timestamp 1586364061
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_249
timestamp 1586364061
transform 1 0 24012 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_260
timestamp 1586364061
transform 1 0 25024 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_37_272
timestamp 1586364061
transform 1 0 26128 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_276
timestamp 1586364061
transform 1 0 26496 0 1 22304
box -38 -48 130 592
use scs8hd_buf_1  mux_left_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2392 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 2208 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__S
timestamp 1586364061
transform 1 0 1840 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_6
timestamp 1586364061
transform 1 0 1656 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_10
timestamp 1586364061
transform 1 0 2024 0 -1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 4692 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4324 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_37
timestamp 1586364061
transform 1 0 4508 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4876 0 -1 23392
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 7820 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7176 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_60
timestamp 1586364061
transform 1 0 6624 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_64
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_72
timestamp 1586364061
transform 1 0 7728 0 -1 23392
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_88
timestamp 1586364061
transform 1 0 9200 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1586364061
transform 1 0 11224 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_102
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_107
timestamp 1586364061
transform 1 0 10948 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_119
timestamp 1586364061
transform 1 0 12052 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12788 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12604 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12236 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13800 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_123
timestamp 1586364061
transform 1 0 12420 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_136
timestamp 1586364061
transform 1 0 13616 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_2  _121_
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14168 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14536 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_140
timestamp 1586364061
transform 1 0 13984 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_144
timestamp 1586364061
transform 1 0 14352 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_148
timestamp 1586364061
transform 1 0 14720 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_158
timestamp 1586364061
transform 1 0 15640 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 16468 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15824 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 16284 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_162
timestamp 1586364061
transform 1 0 16008 0 -1 23392
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1586364061
transform 1 0 18952 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 18676 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_186
timestamp 1586364061
transform 1 0 18216 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_193
timestamp 1586364061
transform 1 0 18860 0 -1 23392
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 20516 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20148 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_203
timestamp 1586364061
transform 1 0 19780 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_209
timestamp 1586364061
transform 1 0 20332 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_213
timestamp 1586364061
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 22448 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 21896 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 22264 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_224
timestamp 1586364061
transform 1 0 21712 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_228
timestamp 1586364061
transform 1 0 22080 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_2  _117_
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 23460 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_241
timestamp 1586364061
transform 1 0 23276 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_245
timestamp 1586364061
transform 1 0 23644 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_253
timestamp 1586364061
transform 1 0 24380 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_259
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_271
timestamp 1586364061
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1586364061
transform 1 0 1656 0 -1 24480
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 866 592
use scs8hd_decap_4  FILLER_40_19
timestamp 1586364061
transform 1 0 2852 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_19
timestamp 1586364061
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 2668 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__S
timestamp 1586364061
transform 1 0 2668 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_29
timestamp 1586364061
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_25
timestamp 1586364061
transform 1 0 3404 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_23
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3220 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__S
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_36
timestamp 1586364061
transform 1 0 4416 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_36
timestamp 1586364061
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 4232 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 4600 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_49
timestamp 1586364061
transform 1 0 5612 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_40
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4968 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1586364061
transform 1 0 4784 0 -1 24480
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 23392
box -38 -48 866 592
use scs8hd_decap_3  FILLER_40_57
timestamp 1586364061
transform 1 0 6348 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_53
timestamp 1586364061
transform 1 0 5980 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__A0
timestamp 1586364061
transform 1 0 6164 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5796 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _057_
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 8096 0 1 23392
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6624 0 -1 24480
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_70
timestamp 1586364061
transform 1 0 7544 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_79
timestamp 1586364061
transform 1 0 8372 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_83
timestamp 1586364061
transform 1 0 8740 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_87
timestamp 1586364061
transform 1 0 9108 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8924 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_91
timestamp 1586364061
transform 1 0 9476 0 -1 24480
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_97
timestamp 1586364061
transform 1 0 10028 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_95
timestamp 1586364061
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 10028 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 9844 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_99
timestamp 1586364061
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10212 0 -1 24480
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10396 0 -1 24480
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_103
timestamp 1586364061
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_114
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_120
timestamp 1586364061
transform 1 0 12144 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_124
timestamp 1586364061
transform 1 0 12512 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_127
timestamp 1586364061
transform 1 0 12788 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_137
timestamp 1586364061
transform 1 0 13708 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_146
timestamp 1586364061
transform 1 0 14536 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_3  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_39_146
timestamp 1586364061
transform 1 0 14536 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_142
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13892 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14352 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_150
timestamp 1586364061
transform 1 0 14904 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_149
timestamp 1586364061
transform 1 0 14812 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15180 0 1 23392
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 17112 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A0
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16744 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 17112 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_172
timestamp 1586364061
transform 1 0 16928 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_176
timestamp 1586364061
transform 1 0 17296 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_40_163
timestamp 1586364061
transform 1 0 16100 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_168
timestamp 1586364061
transform 1 0 16560 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_172
timestamp 1586364061
transform 1 0 16928 0 -1 24480
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1586364061
transform 1 0 18676 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__S
timestamp 1586364061
transform 1 0 18124 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 18492 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_180
timestamp 1586364061
transform 1 0 17664 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_183
timestamp 1586364061
transform 1 0 17940 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_187
timestamp 1586364061
transform 1 0 18308 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_204
timestamp 1586364061
transform 1 0 19872 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_200
timestamp 1586364061
transform 1 0 19504 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_207
timestamp 1586364061
transform 1 0 20148 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_203
timestamp 1586364061
transform 1 0 19780 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20148 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 19964 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_213
timestamp 1586364061
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_209
timestamp 1586364061
transform 1 0 20332 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 20516 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20332 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1586364061
transform 1 0 20516 0 1 23392
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_4  FILLER_40_228
timestamp 1586364061
transform 1 0 22080 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_224
timestamp 1586364061
transform 1 0 21712 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_224
timestamp 1586364061
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 21896 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21528 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 21896 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _126_
timestamp 1586364061
transform 1 0 22080 0 1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_39_236
timestamp 1586364061
transform 1 0 22816 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 22632 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _122_
timestamp 1586364061
transform 1 0 22448 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_236
timestamp 1586364061
transform 1 0 22816 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _116_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _118_
timestamp 1586364061
transform 1 0 24472 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_6  FILLER_40_248
timestamp 1586364061
transform 1 0 23920 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_274
timestamp 1586364061
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_270
timestamp 1586364061
transform 1 0 25944 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_258
timestamp 1586364061
transform 1 0 24840 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _060_
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 406 592
use scs8hd_buf_2  _063_
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 2300 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_7
timestamp 1586364061
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_11
timestamp 1586364061
transform 1 0 2116 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_19
timestamp 1586364061
transform 1 0 2852 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4508 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 3036 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 4048 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3680 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_23
timestamp 1586364061
transform 1 0 3220 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_30
timestamp 1586364061
transform 1 0 3864 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_34
timestamp 1586364061
transform 1 0 4232 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_46
timestamp 1586364061
transform 1 0 5336 0 1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_41_58
timestamp 1586364061
transform 1 0 6440 0 1 24480
box -38 -48 130 592
use scs8hd_conb_1  _052_
timestamp 1586364061
transform 1 0 7084 0 1 24480
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1586364061
transform 1 0 8096 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 7544 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_68
timestamp 1586364061
transform 1 0 7360 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_72
timestamp 1586364061
transform 1 0 7728 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1586364061
transform 1 0 9660 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 9476 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 9108 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_85
timestamp 1586364061
transform 1 0 8924 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_89
timestamp 1586364061
transform 1 0 9292 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _134_
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10948 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_102
timestamp 1586364061
transform 1 0 10488 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_106
timestamp 1586364061
transform 1 0 10856 0 1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_41_109
timestamp 1586364061
transform 1 0 11132 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_114
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 13432 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13800 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_132
timestamp 1586364061
transform 1 0 13248 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_136
timestamp 1586364061
transform 1 0 13616 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 14352 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 14168 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_140
timestamp 1586364061
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_153
timestamp 1586364061
transform 1 0 15180 0 1 24480
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1586364061
transform 1 0 16376 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A1
timestamp 1586364061
transform 1 0 16192 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 17388 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_163
timestamp 1586364061
transform 1 0 16100 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_175
timestamp 1586364061
transform 1 0 17204 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19044 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__A1
timestamp 1586364061
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_179
timestamp 1586364061
transform 1 0 17572 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_193
timestamp 1586364061
transform 1 0 18860 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_197
timestamp 1586364061
transform 1 0 19228 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19596 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 21160 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 20608 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19412 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_210
timestamp 1586364061
transform 1 0 20424 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_214
timestamp 1586364061
transform 1 0 20792 0 1 24480
box -38 -48 406 592
use scs8hd_buf_2  _123_
timestamp 1586364061
transform 1 0 21620 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 22264 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_227
timestamp 1586364061
transform 1 0 21988 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 774 592
use scs8hd_buf_2  _119_
timestamp 1586364061
transform 1 0 23828 0 1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_240
timestamp 1586364061
transform 1 0 23184 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_251
timestamp 1586364061
transform 1 0 24196 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_255
timestamp 1586364061
transform 1 0 24564 0 1 24480
box -38 -48 406 592
use scs8hd_conb_1  _054_
timestamp 1586364061
transform 1 0 24932 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_262
timestamp 1586364061
transform 1 0 25208 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_41_274
timestamp 1586364061
transform 1 0 26312 0 1 24480
box -38 -48 314 592
use scs8hd_buf_2  _059_
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_2  _061_
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__A1
timestamp 1586364061
transform 1 0 1932 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__A0
timestamp 1586364061
transform 1 0 2300 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_7
timestamp 1586364061
transform 1 0 1748 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_11
timestamp 1586364061
transform 1 0 2116 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_19
timestamp 1586364061
transform 1 0 2852 0 -1 25568
box -38 -48 222 592
use scs8hd_buf_2  _058_
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4600 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3036 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__A1
timestamp 1586364061
transform 1 0 3772 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_23
timestamp 1586364061
transform 1 0 3220 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_36
timestamp 1586364061
transform 1 0 4416 0 -1 25568
box -38 -48 222 592
use scs8hd_conb_1  _055_
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4968 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_40
timestamp 1586364061
transform 1 0 4784 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_47
timestamp 1586364061
transform 1 0 5428 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_42_59
timestamp 1586364061
transform 1 0 6532 0 -1 25568
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1586364061
transform 1 0 7544 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 7360 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_67
timestamp 1586364061
transform 1 0 7268 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_79
timestamp 1586364061
transform 1 0 8372 0 -1 25568
box -38 -48 222 592
use scs8hd_buf_2  _131_
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8556 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 9476 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_83
timestamp 1586364061
transform 1 0 8740 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  FILLER_42_98
timestamp 1586364061
transform 1 0 10120 0 -1 25568
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10948 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10396 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_103
timestamp 1586364061
transform 1 0 10580 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_116
timestamp 1586364061
transform 1 0 11776 0 -1 25568
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 13616 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_120
timestamp 1586364061
transform 1 0 12144 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_134
timestamp 1586364061
transform 1 0 13432 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_138
timestamp 1586364061
transform 1 0 13800 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 13984 0 -1 25568
box -38 -48 222 592
use scs8hd_buf_2  _127_
timestamp 1586364061
transform 1 0 14168 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_146
timestamp 1586364061
transform 1 0 14536 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14720 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_150
timestamp 1586364061
transform 1 0 14904 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15088 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_154
timestamp 1586364061
transform 1 0 15272 0 -1 25568
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_buf_2  _130_
timestamp 1586364061
transform 1 0 15548 0 -1 25568
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16652 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__S
timestamp 1586364061
transform 1 0 16376 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_161
timestamp 1586364061
transform 1 0 15916 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_165
timestamp 1586364061
transform 1 0 16284 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_178
timestamp 1586364061
transform 1 0 17480 0 -1 25568
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__A0
timestamp 1586364061
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_182
timestamp 1586364061
transform 1 0 17848 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_196
timestamp 1586364061
transform 1 0 19136 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_203
timestamp 1586364061
transform 1 0 19780 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_200
timestamp 1586364061
transform 1 0 19504 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19596 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_208
timestamp 1586364061
transform 1 0 20240 0 -1 25568
box -38 -48 222 592
use scs8hd_buf_2  _128_
timestamp 1586364061
transform 1 0 19872 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_4  FILLER_42_212
timestamp 1586364061
transform 1 0 20608 0 -1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20424 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_216
timestamp 1586364061
transform 1 0 20976 0 -1 25568
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_buf_2  _124_
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_2  _132_
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 21712 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_222
timestamp 1586364061
transform 1 0 21528 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_226
timestamp 1586364061
transform 1 0 21896 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_234
timestamp 1586364061
transform 1 0 22632 0 -1 25568
box -38 -48 1142 592
use scs8hd_buf_1  mux_right_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_246
timestamp 1586364061
transform 1 0 23736 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_252
timestamp 1586364061
transform 1 0 24288 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_264
timestamp 1586364061
transform 1 0 25392 0 -1 25568
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_42_276
timestamp 1586364061
transform 1 0 26496 0 -1 25568
box -38 -48 130 592
<< labels >>
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_34_
port 0 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_35_
port 1 nsew default input
rlabel metal2 s 1214 0 1270 480 6 bottom_left_grid_pin_36_
port 2 nsew default input
rlabel metal2 s 1766 0 1822 480 6 bottom_left_grid_pin_37_
port 3 nsew default input
rlabel metal2 s 2318 0 2374 480 6 bottom_left_grid_pin_38_
port 4 nsew default input
rlabel metal2 s 2870 0 2926 480 6 bottom_left_grid_pin_39_
port 5 nsew default input
rlabel metal2 s 3422 0 3478 480 6 bottom_left_grid_pin_40_
port 6 nsew default input
rlabel metal2 s 3974 0 4030 480 6 bottom_left_grid_pin_41_
port 7 nsew default input
rlabel metal2 s 5078 0 5134 480 6 ccff_head
port 8 nsew default input
rlabel metal2 s 5630 0 5686 480 6 ccff_tail
port 9 nsew default tristate
rlabel metal3 s 0 280 480 400 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[10]
port 11 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[11]
port 12 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[12]
port 13 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[13]
port 14 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[14]
port 15 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[15]
port 16 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[16]
port 17 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[17]
port 18 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[18]
port 19 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[19]
port 20 nsew default input
rlabel metal3 s 0 824 480 944 6 chanx_left_in[1]
port 21 nsew default input
rlabel metal3 s 0 1368 480 1488 6 chanx_left_in[2]
port 22 nsew default input
rlabel metal3 s 0 1912 480 2032 6 chanx_left_in[3]
port 23 nsew default input
rlabel metal3 s 0 2592 480 2712 6 chanx_left_in[4]
port 24 nsew default input
rlabel metal3 s 0 3136 480 3256 6 chanx_left_in[5]
port 25 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[6]
port 26 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[7]
port 27 nsew default input
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[8]
port 28 nsew default input
rlabel metal3 s 0 5448 480 5568 6 chanx_left_in[9]
port 29 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_out[0]
port 30 nsew default tristate
rlabel metal3 s 0 17688 480 17808 6 chanx_left_out[10]
port 31 nsew default tristate
rlabel metal3 s 0 18368 480 18488 6 chanx_left_out[11]
port 32 nsew default tristate
rlabel metal3 s 0 18912 480 19032 6 chanx_left_out[12]
port 33 nsew default tristate
rlabel metal3 s 0 19456 480 19576 6 chanx_left_out[13]
port 34 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[14]
port 35 nsew default tristate
rlabel metal3 s 0 20680 480 20800 6 chanx_left_out[15]
port 36 nsew default tristate
rlabel metal3 s 0 21224 480 21344 6 chanx_left_out[16]
port 37 nsew default tristate
rlabel metal3 s 0 21768 480 21888 6 chanx_left_out[17]
port 38 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[18]
port 39 nsew default tristate
rlabel metal3 s 0 22992 480 23112 6 chanx_left_out[19]
port 40 nsew default tristate
rlabel metal3 s 0 12520 480 12640 6 chanx_left_out[1]
port 41 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 chanx_left_out[2]
port 42 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[3]
port 43 nsew default tristate
rlabel metal3 s 0 14288 480 14408 6 chanx_left_out[4]
port 44 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 chanx_left_out[5]
port 45 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[6]
port 46 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[7]
port 47 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[8]
port 48 nsew default tristate
rlabel metal3 s 0 17144 480 17264 6 chanx_left_out[9]
port 49 nsew default tristate
rlabel metal3 s 27520 280 28000 400 6 chanx_right_in[0]
port 50 nsew default input
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_in[10]
port 51 nsew default input
rlabel metal3 s 27520 6672 28000 6792 6 chanx_right_in[11]
port 52 nsew default input
rlabel metal3 s 27520 7216 28000 7336 6 chanx_right_in[12]
port 53 nsew default input
rlabel metal3 s 27520 7760 28000 7880 6 chanx_right_in[13]
port 54 nsew default input
rlabel metal3 s 27520 8440 28000 8560 6 chanx_right_in[14]
port 55 nsew default input
rlabel metal3 s 27520 8984 28000 9104 6 chanx_right_in[15]
port 56 nsew default input
rlabel metal3 s 27520 9528 28000 9648 6 chanx_right_in[16]
port 57 nsew default input
rlabel metal3 s 27520 10072 28000 10192 6 chanx_right_in[17]
port 58 nsew default input
rlabel metal3 s 27520 10752 28000 10872 6 chanx_right_in[18]
port 59 nsew default input
rlabel metal3 s 27520 11296 28000 11416 6 chanx_right_in[19]
port 60 nsew default input
rlabel metal3 s 27520 824 28000 944 6 chanx_right_in[1]
port 61 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 chanx_right_in[2]
port 62 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 chanx_right_in[3]
port 63 nsew default input
rlabel metal3 s 27520 2592 28000 2712 6 chanx_right_in[4]
port 64 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 chanx_right_in[5]
port 65 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 chanx_right_in[6]
port 66 nsew default input
rlabel metal3 s 27520 4360 28000 4480 6 chanx_right_in[7]
port 67 nsew default input
rlabel metal3 s 27520 4904 28000 5024 6 chanx_right_in[8]
port 68 nsew default input
rlabel metal3 s 27520 5448 28000 5568 6 chanx_right_in[9]
port 69 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_out[0]
port 70 nsew default tristate
rlabel metal3 s 27520 17688 28000 17808 6 chanx_right_out[10]
port 71 nsew default tristate
rlabel metal3 s 27520 18368 28000 18488 6 chanx_right_out[11]
port 72 nsew default tristate
rlabel metal3 s 27520 18912 28000 19032 6 chanx_right_out[12]
port 73 nsew default tristate
rlabel metal3 s 27520 19456 28000 19576 6 chanx_right_out[13]
port 74 nsew default tristate
rlabel metal3 s 27520 20000 28000 20120 6 chanx_right_out[14]
port 75 nsew default tristate
rlabel metal3 s 27520 20680 28000 20800 6 chanx_right_out[15]
port 76 nsew default tristate
rlabel metal3 s 27520 21224 28000 21344 6 chanx_right_out[16]
port 77 nsew default tristate
rlabel metal3 s 27520 21768 28000 21888 6 chanx_right_out[17]
port 78 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_out[18]
port 79 nsew default tristate
rlabel metal3 s 27520 22992 28000 23112 6 chanx_right_out[19]
port 80 nsew default tristate
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_out[1]
port 81 nsew default tristate
rlabel metal3 s 27520 13064 28000 13184 6 chanx_right_out[2]
port 82 nsew default tristate
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_out[3]
port 83 nsew default tristate
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_out[4]
port 84 nsew default tristate
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_out[5]
port 85 nsew default tristate
rlabel metal3 s 27520 15376 28000 15496 6 chanx_right_out[6]
port 86 nsew default tristate
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_out[7]
port 87 nsew default tristate
rlabel metal3 s 27520 16600 28000 16720 6 chanx_right_out[8]
port 88 nsew default tristate
rlabel metal3 s 27520 17144 28000 17264 6 chanx_right_out[9]
port 89 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[0]
port 90 nsew default input
rlabel metal2 s 11702 0 11758 480 6 chany_bottom_in[10]
port 91 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[11]
port 92 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[12]
port 93 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[13]
port 94 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[14]
port 95 nsew default input
rlabel metal2 s 14370 0 14426 480 6 chany_bottom_in[15]
port 96 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[16]
port 97 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_in[17]
port 98 nsew default input
rlabel metal2 s 16026 0 16082 480 6 chany_bottom_in[18]
port 99 nsew default input
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_in[19]
port 100 nsew default input
rlabel metal2 s 6734 0 6790 480 6 chany_bottom_in[1]
port 101 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[2]
port 102 nsew default input
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_in[3]
port 103 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[4]
port 104 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[5]
port 105 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[6]
port 106 nsew default input
rlabel metal2 s 10046 0 10102 480 6 chany_bottom_in[7]
port 107 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[8]
port 108 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[9]
port 109 nsew default input
rlabel metal2 s 17130 0 17186 480 6 chany_bottom_out[0]
port 110 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[10]
port 111 nsew default tristate
rlabel metal2 s 23202 0 23258 480 6 chany_bottom_out[11]
port 112 nsew default tristate
rlabel metal2 s 23754 0 23810 480 6 chany_bottom_out[12]
port 113 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[13]
port 114 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 chany_bottom_out[14]
port 115 nsew default tristate
rlabel metal2 s 25410 0 25466 480 6 chany_bottom_out[15]
port 116 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[16]
port 117 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[17]
port 118 nsew default tristate
rlabel metal2 s 27066 0 27122 480 6 chany_bottom_out[18]
port 119 nsew default tristate
rlabel metal2 s 27618 0 27674 480 6 chany_bottom_out[19]
port 120 nsew default tristate
rlabel metal2 s 17682 0 17738 480 6 chany_bottom_out[1]
port 121 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chany_bottom_out[2]
port 122 nsew default tristate
rlabel metal2 s 18786 0 18842 480 6 chany_bottom_out[3]
port 123 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chany_bottom_out[4]
port 124 nsew default tristate
rlabel metal2 s 19890 0 19946 480 6 chany_bottom_out[5]
port 125 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 chany_bottom_out[6]
port 126 nsew default tristate
rlabel metal2 s 20994 0 21050 480 6 chany_bottom_out[7]
port 127 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[8]
port 128 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[9]
port 129 nsew default tristate
rlabel metal2 s 4894 27520 4950 28000 6 chany_top_in[0]
port 130 nsew default input
rlabel metal2 s 10782 27520 10838 28000 6 chany_top_in[10]
port 131 nsew default input
rlabel metal2 s 11334 27520 11390 28000 6 chany_top_in[11]
port 132 nsew default input
rlabel metal2 s 11886 27520 11942 28000 6 chany_top_in[12]
port 133 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[13]
port 134 nsew default input
rlabel metal2 s 13082 27520 13138 28000 6 chany_top_in[14]
port 135 nsew default input
rlabel metal2 s 13634 27520 13690 28000 6 chany_top_in[15]
port 136 nsew default input
rlabel metal2 s 14278 27520 14334 28000 6 chany_top_in[16]
port 137 nsew default input
rlabel metal2 s 14830 27520 14886 28000 6 chany_top_in[17]
port 138 nsew default input
rlabel metal2 s 15382 27520 15438 28000 6 chany_top_in[18]
port 139 nsew default input
rlabel metal2 s 16026 27520 16082 28000 6 chany_top_in[19]
port 140 nsew default input
rlabel metal2 s 5538 27520 5594 28000 6 chany_top_in[1]
port 141 nsew default input
rlabel metal2 s 6090 27520 6146 28000 6 chany_top_in[2]
port 142 nsew default input
rlabel metal2 s 6642 27520 6698 28000 6 chany_top_in[3]
port 143 nsew default input
rlabel metal2 s 7286 27520 7342 28000 6 chany_top_in[4]
port 144 nsew default input
rlabel metal2 s 7838 27520 7894 28000 6 chany_top_in[5]
port 145 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chany_top_in[6]
port 146 nsew default input
rlabel metal2 s 9034 27520 9090 28000 6 chany_top_in[7]
port 147 nsew default input
rlabel metal2 s 9586 27520 9642 28000 6 chany_top_in[8]
port 148 nsew default input
rlabel metal2 s 10138 27520 10194 28000 6 chany_top_in[9]
port 149 nsew default input
rlabel metal2 s 16578 27520 16634 28000 6 chany_top_out[0]
port 150 nsew default tristate
rlabel metal2 s 22374 27520 22430 28000 6 chany_top_out[10]
port 151 nsew default tristate
rlabel metal2 s 23018 27520 23074 28000 6 chany_top_out[11]
port 152 nsew default tristate
rlabel metal2 s 23570 27520 23626 28000 6 chany_top_out[12]
port 153 nsew default tristate
rlabel metal2 s 24122 27520 24178 28000 6 chany_top_out[13]
port 154 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[14]
port 155 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[15]
port 156 nsew default tristate
rlabel metal2 s 25870 27520 25926 28000 6 chany_top_out[16]
port 157 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[17]
port 158 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[18]
port 159 nsew default tristate
rlabel metal2 s 27618 27520 27674 28000 6 chany_top_out[19]
port 160 nsew default tristate
rlabel metal2 s 17130 27520 17186 28000 6 chany_top_out[1]
port 161 nsew default tristate
rlabel metal2 s 17774 27520 17830 28000 6 chany_top_out[2]
port 162 nsew default tristate
rlabel metal2 s 18326 27520 18382 28000 6 chany_top_out[3]
port 163 nsew default tristate
rlabel metal2 s 18878 27520 18934 28000 6 chany_top_out[4]
port 164 nsew default tristate
rlabel metal2 s 19522 27520 19578 28000 6 chany_top_out[5]
port 165 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[6]
port 166 nsew default tristate
rlabel metal2 s 20626 27520 20682 28000 6 chany_top_out[7]
port 167 nsew default tristate
rlabel metal2 s 21270 27520 21326 28000 6 chany_top_out[8]
port 168 nsew default tristate
rlabel metal2 s 21822 27520 21878 28000 6 chany_top_out[9]
port 169 nsew default tristate
rlabel metal3 s 0 23536 480 23656 6 left_top_grid_pin_42_
port 170 nsew default input
rlabel metal3 s 0 24080 480 24200 6 left_top_grid_pin_43_
port 171 nsew default input
rlabel metal3 s 0 24760 480 24880 6 left_top_grid_pin_44_
port 172 nsew default input
rlabel metal3 s 0 25304 480 25424 6 left_top_grid_pin_45_
port 173 nsew default input
rlabel metal3 s 0 25848 480 25968 6 left_top_grid_pin_46_
port 174 nsew default input
rlabel metal3 s 0 26528 480 26648 6 left_top_grid_pin_47_
port 175 nsew default input
rlabel metal3 s 0 27072 480 27192 6 left_top_grid_pin_48_
port 176 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_49_
port 177 nsew default input
rlabel metal2 s 4526 0 4582 480 6 prog_clk
port 178 nsew default input
rlabel metal3 s 27520 23536 28000 23656 6 right_top_grid_pin_42_
port 179 nsew default input
rlabel metal3 s 27520 24080 28000 24200 6 right_top_grid_pin_43_
port 180 nsew default input
rlabel metal3 s 27520 24760 28000 24880 6 right_top_grid_pin_44_
port 181 nsew default input
rlabel metal3 s 27520 25304 28000 25424 6 right_top_grid_pin_45_
port 182 nsew default input
rlabel metal3 s 27520 25848 28000 25968 6 right_top_grid_pin_46_
port 183 nsew default input
rlabel metal3 s 27520 26528 28000 26648 6 right_top_grid_pin_47_
port 184 nsew default input
rlabel metal3 s 27520 27072 28000 27192 6 right_top_grid_pin_48_
port 185 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 right_top_grid_pin_49_
port 186 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_34_
port 187 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_35_
port 188 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_36_
port 189 nsew default input
rlabel metal2 s 2042 27520 2098 28000 6 top_left_grid_pin_37_
port 190 nsew default input
rlabel metal2 s 2594 27520 2650 28000 6 top_left_grid_pin_38_
port 191 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_39_
port 192 nsew default input
rlabel metal2 s 3790 27520 3846 28000 6 top_left_grid_pin_40_
port 193 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 top_left_grid_pin_41_
port 194 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 195 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 196 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
