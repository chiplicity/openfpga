magic
tech EFS8A
magscale 1 2
timestamp 1602873500
<< locali >>
rect 19015 23137 19142 23171
rect 23615 18785 23650 18819
rect 16359 17833 16405 17867
rect 16163 17697 16290 17731
rect 21275 14569 21281 14603
rect 21275 14501 21309 14569
rect 6411 14433 6538 14467
rect 7975 12257 8102 12291
rect 15485 11611 15519 11781
rect 15979 11169 16162 11203
rect 15945 10523 15979 10693
rect 21275 10217 21281 10251
rect 21275 10149 21309 10217
rect 12259 8041 12265 8075
rect 12259 7973 12293 8041
rect 7515 7905 7642 7939
rect 18981 7259 19015 7497
rect 7895 7225 8033 7259
rect 6699 6953 6837 6987
rect 11707 6953 11713 6987
rect 21275 6953 21281 6987
rect 11707 6885 11741 6953
rect 21275 6885 21309 6953
rect 6595 6817 6630 6851
rect 6963 6205 7090 6239
rect 10971 6103 11005 6171
rect 10971 6069 10977 6103
rect 10091 5729 10126 5763
rect 9321 4471 9355 4777
rect 16957 4641 17083 4675
rect 16957 4539 16991 4641
rect 3985 4199 4019 4233
rect 2835 4165 2973 4199
rect 3985 4165 4077 4199
rect 12541 4063 12575 4097
rect 12541 4029 12667 4063
rect 8401 3961 8527 3995
rect 8493 3927 8527 3961
rect 11339 3689 11345 3723
rect 17871 3689 17877 3723
rect 11339 3621 11373 3689
rect 17871 3621 17905 3689
rect 2915 3553 3042 3587
rect 12541 3553 12755 3587
rect 15761 3383 15795 3621
rect 2283 3145 2421 3179
rect 15577 2907 15611 3009
<< viali >>
rect 24777 24361 24811 24395
rect 24593 24225 24627 24259
rect 24777 23817 24811 23851
rect 25145 23817 25179 23851
rect 24593 23613 24627 23647
rect 24409 23477 24443 23511
rect 24777 23273 24811 23307
rect 15704 23137 15738 23171
rect 18981 23137 19015 23171
rect 24593 23137 24627 23171
rect 19211 23069 19245 23103
rect 15807 22933 15841 22967
rect 15669 22389 15703 22423
rect 19073 22389 19107 22423
rect 24593 22389 24627 22423
rect 24777 21641 24811 21675
rect 24593 21437 24627 21471
rect 25237 21301 25271 21335
rect 24777 21097 24811 21131
rect 24593 20961 24627 20995
rect 24363 20485 24397 20519
rect 25053 20485 25087 20519
rect 24292 20349 24326 20383
rect 24777 20213 24811 20247
rect 24777 20009 24811 20043
rect 24593 19873 24627 19907
rect 24547 19397 24581 19431
rect 25237 19397 25271 19431
rect 24476 19261 24510 19295
rect 24869 19125 24903 19159
rect 24777 18921 24811 18955
rect 23581 18785 23615 18819
rect 24593 18785 24627 18819
rect 22569 18717 22603 18751
rect 23719 18581 23753 18615
rect 24501 18377 24535 18411
rect 22707 18309 22741 18343
rect 24777 18309 24811 18343
rect 22636 18173 22670 18207
rect 23121 18173 23155 18207
rect 24593 18173 24627 18207
rect 25145 18173 25179 18207
rect 21557 18037 21591 18071
rect 23949 18037 23983 18071
rect 16405 17833 16439 17867
rect 16129 17697 16163 17731
rect 17785 17697 17819 17731
rect 21557 17697 21591 17731
rect 22845 17697 22879 17731
rect 24869 17697 24903 17731
rect 21833 17629 21867 17663
rect 24225 17629 24259 17663
rect 18153 17493 18187 17527
rect 23121 17493 23155 17527
rect 15945 17289 15979 17323
rect 17785 17289 17819 17323
rect 21557 17289 21591 17323
rect 24777 17289 24811 17323
rect 25421 17289 25455 17323
rect 14749 17085 14783 17119
rect 14933 17085 14967 17119
rect 16313 17085 16347 17119
rect 16497 17085 16531 17119
rect 18705 17085 18739 17119
rect 18889 17085 18923 17119
rect 20361 17085 20395 17119
rect 20545 17085 20579 17119
rect 21925 17085 21959 17119
rect 22109 17085 22143 17119
rect 23397 17085 23431 17119
rect 23765 17085 23799 17119
rect 25237 17085 25271 17119
rect 25789 17085 25823 17119
rect 16405 17017 16439 17051
rect 22753 17017 22787 17051
rect 23673 17017 23707 17051
rect 15301 16949 15335 16983
rect 19073 16949 19107 16983
rect 20729 16949 20763 16983
rect 23029 16949 23063 16983
rect 19947 16745 19981 16779
rect 15485 16677 15519 16711
rect 18245 16677 18279 16711
rect 19844 16609 19878 16643
rect 21649 16609 21683 16643
rect 23121 16609 23155 16643
rect 23397 16609 23431 16643
rect 25053 16609 25087 16643
rect 15393 16541 15427 16575
rect 15669 16541 15703 16575
rect 18153 16541 18187 16575
rect 18429 16541 18463 16575
rect 22293 16541 22327 16575
rect 24685 16541 24719 16575
rect 19257 16405 19291 16439
rect 15117 16201 15151 16235
rect 18521 16201 18555 16235
rect 19073 16201 19107 16235
rect 21557 16201 21591 16235
rect 21833 16201 21867 16235
rect 25743 16201 25777 16235
rect 23029 16133 23063 16167
rect 15945 16065 15979 16099
rect 17877 16065 17911 16099
rect 18061 16065 18095 16099
rect 19257 16065 19291 16099
rect 19533 16065 19567 16099
rect 20177 16065 20211 16099
rect 22109 16065 22143 16099
rect 22477 16065 22511 16099
rect 21072 15997 21106 16031
rect 23949 15997 23983 16031
rect 24133 15997 24167 16031
rect 25640 15997 25674 16031
rect 26065 15997 26099 16031
rect 14197 15929 14231 15963
rect 14749 15929 14783 15963
rect 15301 15929 15335 15963
rect 15393 15929 15427 15963
rect 19349 15929 19383 15963
rect 22201 15929 22235 15963
rect 24777 15929 24811 15963
rect 16221 15861 16255 15895
rect 16681 15861 16715 15895
rect 21143 15861 21177 15895
rect 23397 15861 23431 15895
rect 25053 15861 25087 15895
rect 18429 15657 18463 15691
rect 21649 15657 21683 15691
rect 13829 15589 13863 15623
rect 15485 15589 15519 15623
rect 16037 15589 16071 15623
rect 17509 15589 17543 15623
rect 18061 15589 18095 15623
rect 19073 15589 19107 15623
rect 21925 15589 21959 15623
rect 22477 15589 22511 15623
rect 24225 15521 24259 15555
rect 13737 15453 13771 15487
rect 14381 15453 14415 15487
rect 15393 15453 15427 15487
rect 17417 15453 17451 15487
rect 18981 15453 19015 15487
rect 21833 15453 21867 15487
rect 24777 15453 24811 15487
rect 19533 15385 19567 15419
rect 16497 15317 16531 15351
rect 13829 15113 13863 15147
rect 15301 15113 15335 15147
rect 15577 15113 15611 15147
rect 16313 15113 16347 15147
rect 17509 15113 17543 15147
rect 19073 15113 19107 15147
rect 20637 15113 20671 15147
rect 21833 15113 21867 15147
rect 23121 15113 23155 15147
rect 24685 15113 24719 15147
rect 25789 15113 25823 15147
rect 25375 15045 25409 15079
rect 13553 14977 13587 15011
rect 17141 14977 17175 15011
rect 18429 14977 18463 15011
rect 19625 14977 19659 15011
rect 23765 14977 23799 15011
rect 12725 14909 12759 14943
rect 13461 14909 13495 14943
rect 14381 14909 14415 14943
rect 22636 14909 22670 14943
rect 25304 14909 25338 14943
rect 14702 14841 14736 14875
rect 16497 14841 16531 14875
rect 16589 14841 16623 14875
rect 18153 14841 18187 14875
rect 18245 14841 18279 14875
rect 20821 14841 20855 14875
rect 20913 14841 20947 14875
rect 21465 14841 21499 14875
rect 22201 14841 22235 14875
rect 23857 14841 23891 14875
rect 24409 14841 24443 14875
rect 14289 14773 14323 14807
rect 17785 14773 17819 14807
rect 19441 14773 19475 14807
rect 20177 14773 20211 14807
rect 22707 14773 22741 14807
rect 23489 14773 23523 14807
rect 12771 14569 12805 14603
rect 13553 14569 13587 14603
rect 15577 14569 15611 14603
rect 17049 14569 17083 14603
rect 17417 14569 17451 14603
rect 18797 14569 18831 14603
rect 21281 14569 21315 14603
rect 21833 14569 21867 14603
rect 23765 14569 23799 14603
rect 16450 14501 16484 14535
rect 18198 14501 18232 14535
rect 22845 14501 22879 14535
rect 23397 14501 23431 14535
rect 24409 14501 24443 14535
rect 6377 14433 6411 14467
rect 12700 14433 12734 14467
rect 13645 14433 13679 14467
rect 14105 14433 14139 14467
rect 14381 14365 14415 14399
rect 16129 14365 16163 14399
rect 17877 14365 17911 14399
rect 19809 14365 19843 14399
rect 20913 14365 20947 14399
rect 22753 14365 22787 14399
rect 24317 14365 24351 14399
rect 24593 14365 24627 14399
rect 6607 14297 6641 14331
rect 14657 14229 14691 14263
rect 19073 14229 19107 14263
rect 22109 14229 22143 14263
rect 24041 14229 24075 14263
rect 17417 14025 17451 14059
rect 19901 14025 19935 14059
rect 20913 14025 20947 14059
rect 22661 14025 22695 14059
rect 24777 14025 24811 14059
rect 25789 14025 25823 14059
rect 12725 13957 12759 13991
rect 14933 13957 14967 13991
rect 16865 13957 16899 13991
rect 17785 13957 17819 13991
rect 18981 13957 19015 13991
rect 22937 13957 22971 13991
rect 15669 13889 15703 13923
rect 18429 13889 18463 13923
rect 19533 13889 19567 13923
rect 19993 13889 20027 13923
rect 24041 13889 24075 13923
rect 25053 13889 25087 13923
rect 13093 13821 13127 13855
rect 14013 13821 14047 13855
rect 15853 13821 15887 13855
rect 16313 13821 16347 13855
rect 21741 13821 21775 13855
rect 23397 13821 23431 13855
rect 25304 13821 25338 13855
rect 14375 13753 14409 13787
rect 18521 13753 18555 13787
rect 20355 13753 20389 13787
rect 22062 13753 22096 13787
rect 23765 13753 23799 13787
rect 23857 13753 23891 13787
rect 6469 13685 6503 13719
rect 13461 13685 13495 13719
rect 13829 13685 13863 13719
rect 16129 13685 16163 13719
rect 21281 13685 21315 13719
rect 21557 13685 21591 13719
rect 25375 13685 25409 13719
rect 16221 13481 16255 13515
rect 17693 13481 17727 13515
rect 14381 13413 14415 13447
rect 17094 13413 17128 13447
rect 18705 13413 18739 13447
rect 22661 13413 22695 13447
rect 23213 13413 23247 13447
rect 24225 13413 24259 13447
rect 12633 13345 12667 13379
rect 13921 13345 13955 13379
rect 14197 13345 14231 13379
rect 20913 13345 20947 13379
rect 21373 13345 21407 13379
rect 12817 13277 12851 13311
rect 15301 13277 15335 13311
rect 16773 13277 16807 13311
rect 18613 13277 18647 13311
rect 18889 13277 18923 13311
rect 21649 13277 21683 13311
rect 21925 13277 21959 13311
rect 22569 13277 22603 13311
rect 24133 13277 24167 13311
rect 17969 13209 18003 13243
rect 24685 13209 24719 13243
rect 14657 13141 14691 13175
rect 15853 13141 15887 13175
rect 18337 13141 18371 13175
rect 19809 13141 19843 13175
rect 20637 13141 20671 13175
rect 23581 13141 23615 13175
rect 23949 13141 23983 13175
rect 12173 12937 12207 12971
rect 18981 12937 19015 12971
rect 19257 12937 19291 12971
rect 22293 12937 22327 12971
rect 22661 12937 22695 12971
rect 24869 12937 24903 12971
rect 25559 12869 25593 12903
rect 13737 12801 13771 12835
rect 14657 12801 14691 12835
rect 15301 12801 15335 12835
rect 16773 12801 16807 12835
rect 18061 12801 18095 12835
rect 20545 12801 20579 12835
rect 21373 12801 21407 12835
rect 23949 12801 23983 12835
rect 24593 12801 24627 12835
rect 12909 12733 12943 12767
rect 13277 12733 13311 12767
rect 13553 12733 13587 12767
rect 16129 12733 16163 12767
rect 16681 12733 16715 12767
rect 17233 12733 17267 12767
rect 17877 12733 17911 12767
rect 19809 12733 19843 12767
rect 20269 12733 20303 12767
rect 25488 12733 25522 12767
rect 25973 12733 26007 12767
rect 14749 12665 14783 12699
rect 15669 12665 15703 12699
rect 18423 12665 18457 12699
rect 21694 12665 21728 12699
rect 23489 12665 23523 12699
rect 24041 12665 24075 12699
rect 14013 12597 14047 12631
rect 14473 12597 14507 12631
rect 16037 12597 16071 12631
rect 19625 12597 19659 12631
rect 20821 12597 20855 12631
rect 21281 12597 21315 12631
rect 22937 12597 22971 12631
rect 8171 12393 8205 12427
rect 13093 12393 13127 12427
rect 16773 12393 16807 12427
rect 18705 12393 18739 12427
rect 20637 12393 20671 12427
rect 22109 12393 22143 12427
rect 23029 12393 23063 12427
rect 24133 12393 24167 12427
rect 24593 12393 24627 12427
rect 12541 12325 12575 12359
rect 15485 12325 15519 12359
rect 18429 12325 18463 12359
rect 21510 12325 21544 12359
rect 7941 12257 7975 12291
rect 12081 12257 12115 12291
rect 12357 12257 12391 12291
rect 13369 12257 13403 12291
rect 13829 12257 13863 12291
rect 17693 12257 17727 12291
rect 19257 12257 19291 12291
rect 19717 12257 19751 12291
rect 23029 12257 23063 12291
rect 23351 12257 23385 12291
rect 24685 12257 24719 12291
rect 24961 12257 24995 12291
rect 14105 12189 14139 12223
rect 15393 12189 15427 12223
rect 15669 12189 15703 12223
rect 17840 12189 17874 12223
rect 18061 12189 18095 12223
rect 19993 12189 20027 12223
rect 20361 12189 20395 12223
rect 21189 12189 21223 12223
rect 14565 12053 14599 12087
rect 14933 12053 14967 12087
rect 16313 12053 16347 12087
rect 17601 12053 17635 12087
rect 17969 12053 18003 12087
rect 19073 12053 19107 12087
rect 11897 11849 11931 11883
rect 13001 11849 13035 11883
rect 16589 11849 16623 11883
rect 22017 11849 22051 11883
rect 23397 11849 23431 11883
rect 24685 11849 24719 11883
rect 25053 11849 25087 11883
rect 25789 11849 25823 11883
rect 14749 11781 14783 11815
rect 15485 11781 15519 11815
rect 22569 11781 22603 11815
rect 25375 11781 25409 11815
rect 11529 11713 11563 11747
rect 10701 11645 10735 11679
rect 11437 11645 11471 11679
rect 13829 11645 13863 11679
rect 15945 11713 15979 11747
rect 18981 11713 19015 11747
rect 20269 11713 20303 11747
rect 24041 11713 24075 11747
rect 18061 11645 18095 11679
rect 19533 11645 19567 11679
rect 19993 11645 20027 11679
rect 21097 11645 21131 11679
rect 25304 11645 25338 11679
rect 12265 11577 12299 11611
rect 14191 11577 14225 11611
rect 15485 11577 15519 11611
rect 15658 11577 15692 11611
rect 15761 11577 15795 11611
rect 17325 11577 17359 11611
rect 21418 11577 21452 11611
rect 23765 11577 23799 11611
rect 23857 11577 23891 11611
rect 8033 11509 8067 11543
rect 13277 11509 13311 11543
rect 13737 11509 13771 11543
rect 15301 11509 15335 11543
rect 17049 11509 17083 11543
rect 17785 11509 17819 11543
rect 18245 11509 18279 11543
rect 18613 11509 18647 11543
rect 19349 11509 19383 11543
rect 20637 11509 20671 11543
rect 20913 11509 20947 11543
rect 22937 11509 22971 11543
rect 14565 11305 14599 11339
rect 15117 11305 15151 11339
rect 17509 11305 17543 11339
rect 20637 11305 20671 11339
rect 21189 11305 21223 11339
rect 13690 11237 13724 11271
rect 16865 11237 16899 11271
rect 17693 11237 17727 11271
rect 18429 11237 18463 11271
rect 20269 11237 20303 11271
rect 23673 11237 23707 11271
rect 11897 11169 11931 11203
rect 12541 11169 12575 11203
rect 15945 11169 15979 11203
rect 19257 11169 19291 11203
rect 19809 11169 19843 11203
rect 20913 11169 20947 11203
rect 21465 11169 21499 11203
rect 25120 11169 25154 11203
rect 13369 11101 13403 11135
rect 16497 11101 16531 11135
rect 18061 11101 18095 11135
rect 19993 11101 20027 11135
rect 22477 11101 22511 11135
rect 23581 11101 23615 11135
rect 23949 11101 23983 11135
rect 14289 11033 14323 11067
rect 16405 11033 16439 11067
rect 17969 11033 18003 11067
rect 19073 11033 19107 11067
rect 21925 11033 21959 11067
rect 13185 10965 13219 10999
rect 15577 10965 15611 10999
rect 16294 10965 16328 10999
rect 17233 10965 17267 10999
rect 17858 10965 17892 10999
rect 18705 10965 18739 10999
rect 24501 10965 24535 10999
rect 25191 10965 25225 10999
rect 11897 10761 11931 10795
rect 16773 10761 16807 10795
rect 20637 10761 20671 10795
rect 22293 10761 22327 10795
rect 23029 10761 23063 10795
rect 25145 10761 25179 10795
rect 12633 10693 12667 10727
rect 15945 10693 15979 10727
rect 16589 10693 16623 10727
rect 18337 10693 18371 10727
rect 19809 10693 19843 10727
rect 22661 10693 22695 10727
rect 23489 10693 23523 10727
rect 24685 10693 24719 10727
rect 14197 10625 14231 10659
rect 7364 10557 7398 10591
rect 12449 10557 12483 10591
rect 12909 10557 12943 10591
rect 15301 10557 15335 10591
rect 15853 10557 15887 10591
rect 16681 10625 16715 10659
rect 18429 10625 18463 10659
rect 18797 10625 18831 10659
rect 21097 10625 21131 10659
rect 23765 10625 23799 10659
rect 24041 10625 24075 10659
rect 16460 10557 16494 10591
rect 18208 10557 18242 10591
rect 19625 10557 19659 10591
rect 20085 10557 20119 10591
rect 22017 10557 22051 10591
rect 13553 10489 13587 10523
rect 13645 10489 13679 10523
rect 15209 10489 15243 10523
rect 15945 10489 15979 10523
rect 16313 10489 16347 10523
rect 18061 10489 18095 10523
rect 21418 10489 21452 10523
rect 23857 10489 23891 10523
rect 7435 10421 7469 10455
rect 7757 10421 7791 10455
rect 13277 10421 13311 10455
rect 14473 10421 14507 10455
rect 15485 10421 15519 10455
rect 16221 10421 16255 10455
rect 17417 10421 17451 10455
rect 17693 10421 17727 10455
rect 19257 10421 19291 10455
rect 21005 10421 21039 10455
rect 25237 10421 25271 10455
rect 12909 10217 12943 10251
rect 13185 10217 13219 10251
rect 17233 10217 17267 10251
rect 19257 10217 19291 10251
rect 21281 10217 21315 10251
rect 21833 10217 21867 10251
rect 11529 10149 11563 10183
rect 17785 10149 17819 10183
rect 23489 10149 23523 10183
rect 24041 10149 24075 10183
rect 25053 10149 25087 10183
rect 11676 10081 11710 10115
rect 13093 10081 13127 10115
rect 13553 10081 13587 10115
rect 16405 10081 16439 10115
rect 19349 10081 19383 10115
rect 11897 10013 11931 10047
rect 15577 10013 15611 10047
rect 18153 10013 18187 10047
rect 18521 10013 18555 10047
rect 19809 10013 19843 10047
rect 20913 10013 20947 10047
rect 23397 10013 23431 10047
rect 24961 10013 24995 10047
rect 16773 9945 16807 9979
rect 17601 9945 17635 9979
rect 17923 9945 17957 9979
rect 18797 9945 18831 9979
rect 25513 9945 25547 9979
rect 10885 9877 10919 9911
rect 11805 9877 11839 9911
rect 12173 9877 12207 9911
rect 14197 9877 14231 9911
rect 15025 9877 15059 9911
rect 16221 9877 16255 9911
rect 18061 9877 18095 9911
rect 19533 9877 19567 9911
rect 11805 9673 11839 9707
rect 12725 9673 12759 9707
rect 13093 9673 13127 9707
rect 14086 9673 14120 9707
rect 16589 9673 16623 9707
rect 17049 9673 17083 9707
rect 22201 9673 22235 9707
rect 23121 9673 23155 9707
rect 23397 9673 23431 9707
rect 24961 9673 24995 9707
rect 25789 9673 25823 9707
rect 26065 9673 26099 9707
rect 9965 9605 9999 9639
rect 14197 9605 14231 9639
rect 17417 9605 17451 9639
rect 13737 9537 13771 9571
rect 14381 9537 14415 9571
rect 18889 9537 18923 9571
rect 22753 9537 22787 9571
rect 24041 9537 24075 9571
rect 9781 9469 9815 9503
rect 10885 9469 10919 9503
rect 12909 9469 12943 9503
rect 13369 9469 13403 9503
rect 14260 9469 14294 9503
rect 15393 9469 15427 9503
rect 15577 9469 15611 9503
rect 17785 9469 17819 9503
rect 18061 9469 18095 9503
rect 18521 9469 18555 9503
rect 19257 9469 19291 9503
rect 19441 9469 19475 9503
rect 19901 9469 19935 9503
rect 20177 9469 20211 9503
rect 21005 9469 21039 9503
rect 25288 9469 25322 9503
rect 10333 9401 10367 9435
rect 11529 9401 11563 9435
rect 13921 9401 13955 9435
rect 16221 9401 16255 9435
rect 21326 9401 21360 9435
rect 23765 9401 23799 9435
rect 23857 9401 23891 9435
rect 25375 9401 25409 9435
rect 10609 9333 10643 9367
rect 12173 9333 12207 9367
rect 14933 9333 14967 9367
rect 18245 9333 18279 9367
rect 20545 9333 20579 9367
rect 20821 9333 20855 9367
rect 21925 9333 21959 9367
rect 21097 9129 21131 9163
rect 22201 9129 22235 9163
rect 13553 9061 13587 9095
rect 14473 9061 14507 9095
rect 15301 9061 15335 9095
rect 17877 9061 17911 9095
rect 21602 9061 21636 9095
rect 23213 9061 23247 9095
rect 24777 9061 24811 9095
rect 25329 9061 25363 9095
rect 10885 8993 10919 9027
rect 11989 8993 12023 9027
rect 12357 8993 12391 9027
rect 15393 8993 15427 9027
rect 17141 8993 17175 9027
rect 17325 8993 17359 9027
rect 19257 8993 19291 9027
rect 19809 8993 19843 9027
rect 10977 8925 11011 8959
rect 12541 8925 12575 8959
rect 13461 8925 13495 8959
rect 17601 8925 17635 8959
rect 19993 8925 20027 8959
rect 21281 8925 21315 8959
rect 23121 8925 23155 8959
rect 23397 8925 23431 8959
rect 24685 8925 24719 8959
rect 14013 8857 14047 8891
rect 11529 8789 11563 8823
rect 13093 8789 13127 8823
rect 16313 8789 16347 8823
rect 18889 8789 18923 8823
rect 22569 8789 22603 8823
rect 24041 8789 24075 8823
rect 9321 8585 9355 8619
rect 9689 8585 9723 8619
rect 9965 8585 9999 8619
rect 11897 8585 11931 8619
rect 12265 8585 12299 8619
rect 14105 8585 14139 8619
rect 15945 8585 15979 8619
rect 16957 8585 16991 8619
rect 17325 8585 17359 8619
rect 19901 8585 19935 8619
rect 23121 8585 23155 8619
rect 23397 8585 23431 8619
rect 24777 8585 24811 8619
rect 25789 8585 25823 8619
rect 8907 8517 8941 8551
rect 13737 8517 13771 8551
rect 15761 8517 15795 8551
rect 16497 8517 16531 8551
rect 19441 8517 19475 8551
rect 21097 8517 21131 8551
rect 22661 8517 22695 8551
rect 10701 8449 10735 8483
rect 12541 8449 12575 8483
rect 14289 8449 14323 8483
rect 15632 8449 15666 8483
rect 15853 8449 15887 8483
rect 18889 8449 18923 8483
rect 22109 8449 22143 8483
rect 8836 8381 8870 8415
rect 9781 8381 9815 8415
rect 11069 8381 11103 8415
rect 11345 8381 11379 8415
rect 18613 8381 18647 8415
rect 25304 8381 25338 8415
rect 10333 8313 10367 8347
rect 11529 8313 11563 8347
rect 12862 8313 12896 8347
rect 15025 8313 15059 8347
rect 15485 8313 15519 8347
rect 18981 8313 19015 8347
rect 20545 8313 20579 8347
rect 20637 8313 20671 8347
rect 22201 8313 22235 8347
rect 23765 8313 23799 8347
rect 23857 8313 23891 8347
rect 24409 8313 24443 8347
rect 25053 8313 25087 8347
rect 13461 8245 13495 8279
rect 15301 8245 15335 8279
rect 20361 8245 20395 8279
rect 21465 8245 21499 8279
rect 21833 8245 21867 8279
rect 25375 8245 25409 8279
rect 7711 8041 7745 8075
rect 8769 8041 8803 8075
rect 12265 8041 12299 8075
rect 13093 8041 13127 8075
rect 18613 8041 18647 8075
rect 19717 8041 19751 8075
rect 20545 8041 20579 8075
rect 21281 8041 21315 8075
rect 23121 8041 23155 8075
rect 23765 8041 23799 8075
rect 25559 8041 25593 8075
rect 13461 7973 13495 8007
rect 13829 7973 13863 8007
rect 18014 7973 18048 8007
rect 19257 7973 19291 8007
rect 22154 7973 22188 8007
rect 24041 7973 24075 8007
rect 7481 7905 7515 7939
rect 8585 7905 8619 7939
rect 10425 7905 10459 7939
rect 11897 7905 11931 7939
rect 15301 7905 15335 7939
rect 17693 7905 17727 7939
rect 19441 7905 19475 7939
rect 19625 7905 19659 7939
rect 22753 7905 22787 7939
rect 25488 7905 25522 7939
rect 13737 7837 13771 7871
rect 14013 7837 14047 7871
rect 15669 7837 15703 7871
rect 21833 7837 21867 7871
rect 23949 7837 23983 7871
rect 24409 7837 24443 7871
rect 12817 7769 12851 7803
rect 15761 7769 15795 7803
rect 10149 7701 10183 7735
rect 10609 7701 10643 7735
rect 11437 7701 11471 7735
rect 11805 7701 11839 7735
rect 14657 7701 14691 7735
rect 15025 7701 15059 7735
rect 15439 7701 15473 7735
rect 15577 7701 15611 7735
rect 16313 7701 16347 7735
rect 16681 7701 16715 7735
rect 7665 7497 7699 7531
rect 8309 7497 8343 7531
rect 8953 7497 8987 7531
rect 9689 7497 9723 7531
rect 10609 7497 10643 7531
rect 13921 7497 13955 7531
rect 14289 7497 14323 7531
rect 15393 7497 15427 7531
rect 16083 7497 16117 7531
rect 17325 7497 17359 7531
rect 18705 7497 18739 7531
rect 18981 7497 19015 7531
rect 19165 7497 19199 7531
rect 21833 7497 21867 7531
rect 23397 7497 23431 7531
rect 25513 7497 25547 7531
rect 9965 7429 9999 7463
rect 11437 7429 11471 7463
rect 14657 7429 14691 7463
rect 16221 7429 16255 7463
rect 10885 7361 10919 7395
rect 12725 7361 12759 7395
rect 13001 7361 13035 7395
rect 14528 7361 14562 7395
rect 14749 7361 14783 7395
rect 15853 7361 15887 7395
rect 16313 7361 16347 7395
rect 16681 7361 16715 7395
rect 7824 7293 7858 7327
rect 8769 7293 8803 7327
rect 9781 7293 9815 7327
rect 11989 7293 12023 7327
rect 14381 7293 14415 7327
rect 15945 7293 15979 7327
rect 17785 7293 17819 7327
rect 20729 7429 20763 7463
rect 19349 7361 19383 7395
rect 19625 7361 19659 7395
rect 20821 7361 20855 7395
rect 22109 7361 22143 7395
rect 24409 7361 24443 7395
rect 24685 7361 24719 7395
rect 24133 7293 24167 7327
rect 8033 7225 8067 7259
rect 10977 7225 11011 7259
rect 12817 7225 12851 7259
rect 18245 7225 18279 7259
rect 18981 7225 19015 7259
rect 19441 7225 19475 7259
rect 21557 7225 21591 7259
rect 22201 7225 22235 7259
rect 22753 7225 22787 7259
rect 24501 7225 24535 7259
rect 8677 7157 8711 7191
rect 9229 7157 9263 7191
rect 10333 7157 10367 7191
rect 15025 7157 15059 7191
rect 16957 7157 16991 7191
rect 20269 7157 20303 7191
rect 6837 6953 6871 6987
rect 8769 6953 8803 6987
rect 11253 6953 11287 6987
rect 11713 6953 11747 6987
rect 12725 6953 12759 6987
rect 13185 6953 13219 6987
rect 14381 6953 14415 6987
rect 15117 6953 15151 6987
rect 15945 6953 15979 6987
rect 17325 6953 17359 6987
rect 17693 6953 17727 6987
rect 21281 6953 21315 6987
rect 23949 6953 23983 6987
rect 24409 6953 24443 6987
rect 7711 6885 7745 6919
rect 10793 6885 10827 6919
rect 23121 6885 23155 6919
rect 24685 6885 24719 6919
rect 6561 6817 6595 6851
rect 7624 6817 7658 6851
rect 8585 6817 8619 6851
rect 9137 6817 9171 6851
rect 10149 6817 10183 6851
rect 12265 6817 12299 6851
rect 13369 6817 13403 6851
rect 13645 6817 13679 6851
rect 15301 6817 15335 6851
rect 16313 6817 16347 6851
rect 16865 6817 16899 6851
rect 17877 6817 17911 6851
rect 19073 6817 19107 6851
rect 19717 6817 19751 6851
rect 19901 6817 19935 6851
rect 22477 6817 22511 6851
rect 10517 6749 10551 6783
rect 11345 6749 11379 6783
rect 17049 6749 17083 6783
rect 20913 6749 20947 6783
rect 23029 6749 23063 6783
rect 24593 6749 24627 6783
rect 24869 6749 24903 6783
rect 9505 6681 9539 6715
rect 18705 6681 18739 6715
rect 23581 6681 23615 6715
rect 7113 6613 7147 6647
rect 8125 6613 8159 6647
rect 15485 6613 15519 6647
rect 18061 6613 18095 6647
rect 18429 6613 18463 6647
rect 19993 6613 20027 6647
rect 21833 6613 21867 6647
rect 22201 6613 22235 6647
rect 6653 6409 6687 6443
rect 7573 6409 7607 6443
rect 9210 6409 9244 6443
rect 10149 6409 10183 6443
rect 10517 6409 10551 6443
rect 11897 6409 11931 6443
rect 12173 6409 12207 6443
rect 13461 6409 13495 6443
rect 13921 6409 13955 6443
rect 16175 6409 16209 6443
rect 16313 6409 16347 6443
rect 17417 6409 17451 6443
rect 24685 6409 24719 6443
rect 9321 6341 9355 6375
rect 17785 6341 17819 6375
rect 22017 6341 22051 6375
rect 23029 6341 23063 6375
rect 25053 6341 25087 6375
rect 25421 6341 25455 6375
rect 9413 6273 9447 6307
rect 10609 6273 10643 6307
rect 16405 6273 16439 6307
rect 17049 6273 17083 6307
rect 19901 6273 19935 6307
rect 21097 6273 21131 6307
rect 22293 6273 22327 6307
rect 23489 6273 23523 6307
rect 6929 6205 6963 6239
rect 8068 6205 8102 6239
rect 8171 6205 8205 6239
rect 12449 6205 12483 6239
rect 13001 6205 13035 6239
rect 14473 6205 14507 6239
rect 15025 6205 15059 6239
rect 18521 6205 18555 6239
rect 18889 6205 18923 6239
rect 18981 6205 19015 6239
rect 19809 6205 19843 6239
rect 20085 6205 20119 6239
rect 23765 6205 23799 6239
rect 25237 6205 25271 6239
rect 25789 6205 25823 6239
rect 9045 6137 9079 6171
rect 15209 6137 15243 6171
rect 16037 6137 16071 6171
rect 16773 6137 16807 6171
rect 20545 6137 20579 6171
rect 21005 6137 21039 6171
rect 21418 6137 21452 6171
rect 23673 6137 23707 6171
rect 7159 6069 7193 6103
rect 8585 6069 8619 6103
rect 9689 6069 9723 6103
rect 10977 6069 11011 6103
rect 11529 6069 11563 6103
rect 12541 6069 12575 6103
rect 14289 6069 14323 6103
rect 15485 6069 15519 6103
rect 15853 6069 15887 6103
rect 9045 5865 9079 5899
rect 9413 5865 9447 5899
rect 10701 5865 10735 5899
rect 12173 5865 12207 5899
rect 13737 5865 13771 5899
rect 15117 5865 15151 5899
rect 16129 5865 16163 5899
rect 21097 5865 21131 5899
rect 23029 5865 23063 5899
rect 7159 5797 7193 5831
rect 11161 5797 11195 5831
rect 11253 5797 11287 5831
rect 12449 5797 12483 5831
rect 12817 5797 12851 5831
rect 18429 5797 18463 5831
rect 21465 5797 21499 5831
rect 23489 5797 23523 5831
rect 25053 5797 25087 5831
rect 6076 5729 6110 5763
rect 7072 5729 7106 5763
rect 8033 5729 8067 5763
rect 10057 5729 10091 5763
rect 10195 5729 10229 5763
rect 15301 5729 15335 5763
rect 17049 5729 17083 5763
rect 18889 5729 18923 5763
rect 19717 5729 19751 5763
rect 19901 5729 19935 5763
rect 21557 5729 21591 5763
rect 8401 5661 8435 5695
rect 11805 5661 11839 5695
rect 12725 5661 12759 5695
rect 13001 5661 13035 5695
rect 14197 5661 14231 5695
rect 16405 5661 16439 5695
rect 23397 5661 23431 5695
rect 23673 5661 23707 5695
rect 24961 5661 24995 5695
rect 25237 5661 25271 5695
rect 8198 5593 8232 5627
rect 18705 5593 18739 5627
rect 6147 5525 6181 5559
rect 7665 5525 7699 5559
rect 8309 5525 8343 5559
rect 8677 5525 8711 5559
rect 14105 5525 14139 5559
rect 14657 5525 14691 5559
rect 15485 5525 15519 5559
rect 17877 5525 17911 5559
rect 19993 5525 20027 5559
rect 5871 5321 5905 5355
rect 6653 5321 6687 5355
rect 7113 5321 7147 5355
rect 7481 5321 7515 5355
rect 8401 5321 8435 5355
rect 11253 5321 11287 5355
rect 12173 5321 12207 5355
rect 14565 5321 14599 5355
rect 14933 5321 14967 5355
rect 15669 5321 15703 5355
rect 16313 5321 16347 5355
rect 17325 5321 17359 5355
rect 18521 5321 18555 5355
rect 18889 5321 18923 5355
rect 21281 5321 21315 5355
rect 21557 5321 21591 5355
rect 23121 5321 23155 5355
rect 24961 5321 24995 5355
rect 10057 5253 10091 5287
rect 11621 5253 11655 5287
rect 10241 5185 10275 5219
rect 10885 5185 10919 5219
rect 13001 5185 13035 5219
rect 14804 5185 14838 5219
rect 15025 5185 15059 5219
rect 21741 5185 21775 5219
rect 4788 5117 4822 5151
rect 5800 5117 5834 5151
rect 7640 5117 7674 5151
rect 8861 5117 8895 5151
rect 9137 5117 9171 5151
rect 13185 5117 13219 5151
rect 13553 5117 13587 5151
rect 16221 5117 16255 5151
rect 16773 5117 16807 5151
rect 19073 5117 19107 5151
rect 19901 5117 19935 5151
rect 20085 5117 20119 5151
rect 20821 5117 20855 5151
rect 25237 5117 25271 5151
rect 25789 5117 25823 5151
rect 9321 5049 9355 5083
rect 10333 5049 10367 5083
rect 14657 5049 14691 5083
rect 20453 5049 20487 5083
rect 22062 5049 22096 5083
rect 23765 5049 23799 5083
rect 23857 5049 23891 5083
rect 24409 5049 24443 5083
rect 4859 4981 4893 5015
rect 5273 4981 5307 5015
rect 6285 4981 6319 5015
rect 7711 4981 7745 5015
rect 8125 4981 8159 5015
rect 9689 4981 9723 5015
rect 13185 4981 13219 5015
rect 14197 4981 14231 5015
rect 15301 4981 15335 5015
rect 16037 4981 16071 5015
rect 18061 4981 18095 5015
rect 20177 4981 20211 5015
rect 22661 4981 22695 5015
rect 23489 4981 23523 5015
rect 25421 4981 25455 5015
rect 4767 4777 4801 4811
rect 5779 4777 5813 4811
rect 7941 4777 7975 4811
rect 9045 4777 9079 4811
rect 9321 4777 9355 4811
rect 9505 4777 9539 4811
rect 10885 4777 10919 4811
rect 13461 4777 13495 4811
rect 13737 4777 13771 4811
rect 14657 4777 14691 4811
rect 16681 4777 16715 4811
rect 18521 4777 18555 4811
rect 18889 4777 18923 4811
rect 21741 4777 21775 4811
rect 23397 4777 23431 4811
rect 23765 4777 23799 4811
rect 24961 4777 24995 4811
rect 4696 4641 4730 4675
rect 5708 4641 5742 4675
rect 7088 4641 7122 4675
rect 8309 4641 8343 4675
rect 8585 4641 8619 4675
rect 8769 4573 8803 4607
rect 9873 4709 9907 4743
rect 11621 4709 11655 4743
rect 19257 4709 19291 4743
rect 22338 4709 22372 4743
rect 24133 4709 24167 4743
rect 24685 4709 24719 4743
rect 10517 4641 10551 4675
rect 13645 4641 13679 4675
rect 14197 4641 14231 4675
rect 15301 4641 15335 4675
rect 15531 4641 15565 4675
rect 17509 4641 17543 4675
rect 20913 4641 20947 4675
rect 11529 4573 11563 4607
rect 11805 4573 11839 4607
rect 13093 4573 13127 4607
rect 15669 4573 15703 4607
rect 17785 4573 17819 4607
rect 18061 4573 18095 4607
rect 19165 4573 19199 4607
rect 19441 4573 19475 4607
rect 22017 4573 22051 4607
rect 24041 4573 24075 4607
rect 15117 4505 15151 4539
rect 16313 4505 16347 4539
rect 16957 4505 16991 4539
rect 21097 4505 21131 4539
rect 22937 4505 22971 4539
rect 7159 4437 7193 4471
rect 9321 4437 9355 4471
rect 12725 4437 12759 4471
rect 15439 4437 15473 4471
rect 15945 4437 15979 4471
rect 1547 4233 1581 4267
rect 3985 4233 4019 4267
rect 4859 4233 4893 4267
rect 13645 4233 13679 4267
rect 16773 4233 16807 4267
rect 17141 4233 17175 4267
rect 17785 4233 17819 4267
rect 18981 4233 19015 4267
rect 19257 4233 19291 4267
rect 22385 4233 22419 4267
rect 23397 4233 23431 4267
rect 2973 4165 3007 4199
rect 4077 4165 4111 4199
rect 8769 4165 8803 4199
rect 10333 4165 10367 4199
rect 11805 4165 11839 4199
rect 23029 4165 23063 4199
rect 7573 4097 7607 4131
rect 12173 4097 12207 4131
rect 12541 4097 12575 4131
rect 18061 4097 18095 4131
rect 22569 4097 22603 4131
rect 1444 4029 1478 4063
rect 2764 4029 2798 4063
rect 3776 4029 3810 4063
rect 4788 4029 4822 4063
rect 5800 4029 5834 4063
rect 6561 4029 6595 4063
rect 8125 4029 8159 4063
rect 9137 4029 9171 4063
rect 9321 4029 9355 4063
rect 10701 4029 10735 4063
rect 11345 4029 11379 4063
rect 11529 4029 11563 4063
rect 13093 4029 13127 4063
rect 15761 4029 15795 4063
rect 16221 4029 16255 4063
rect 20269 4029 20303 4063
rect 20821 4029 20855 4063
rect 23949 4029 23983 4063
rect 24593 4029 24627 4063
rect 25513 4029 25547 4063
rect 26065 4029 26099 4063
rect 5641 3961 5675 3995
rect 13369 3961 13403 3995
rect 14289 3961 14323 3995
rect 14381 3961 14415 3995
rect 14933 3961 14967 3995
rect 15393 3961 15427 3995
rect 18382 3961 18416 3995
rect 21142 3961 21176 3995
rect 22017 3961 22051 3995
rect 1869 3893 1903 3927
rect 3249 3893 3283 3927
rect 3847 3893 3881 3927
rect 4261 3893 4295 3927
rect 5181 3893 5215 3927
rect 5871 3893 5905 3927
rect 6193 3893 6227 3927
rect 7113 3893 7147 3927
rect 8493 3893 8527 3927
rect 9689 3893 9723 3927
rect 14013 3893 14047 3927
rect 15853 3893 15887 3927
rect 19625 3893 19659 3927
rect 19809 3893 19843 3927
rect 20729 3893 20763 3927
rect 21741 3893 21775 3927
rect 25697 3893 25731 3927
rect 6745 3689 6779 3723
rect 9827 3689 9861 3723
rect 11345 3689 11379 3723
rect 12173 3689 12207 3723
rect 14013 3689 14047 3723
rect 15025 3689 15059 3723
rect 15485 3689 15519 3723
rect 17141 3689 17175 3723
rect 17877 3689 17911 3723
rect 23581 3689 23615 3723
rect 24409 3689 24443 3723
rect 5273 3621 5307 3655
rect 12541 3621 12575 3655
rect 13087 3621 13121 3655
rect 15761 3621 15795 3655
rect 15945 3621 15979 3655
rect 16037 3621 16071 3655
rect 19441 3621 19475 3655
rect 21234 3621 21268 3655
rect 24961 3621 24995 3655
rect 25053 3621 25087 3655
rect 2881 3553 2915 3587
rect 4512 3553 4546 3587
rect 6653 3553 6687 3587
rect 8677 3553 8711 3587
rect 9756 3553 9790 3587
rect 5457 3485 5491 3519
rect 8769 3485 8803 3519
rect 10977 3485 11011 3519
rect 4583 3417 4617 3451
rect 10793 3417 10827 3451
rect 14289 3417 14323 3451
rect 19073 3553 19107 3587
rect 23489 3553 23523 3587
rect 17509 3485 17543 3519
rect 18705 3485 18739 3519
rect 19349 3485 19383 3519
rect 19625 3485 19659 3519
rect 20913 3485 20947 3519
rect 25237 3485 25271 3519
rect 16497 3417 16531 3451
rect 3111 3349 3145 3383
rect 7757 3349 7791 3383
rect 11897 3349 11931 3383
rect 13645 3349 13679 3383
rect 14657 3349 14691 3383
rect 15761 3349 15795 3383
rect 18429 3349 18463 3383
rect 20269 3349 20303 3383
rect 20637 3349 20671 3383
rect 21833 3349 21867 3383
rect 2421 3145 2455 3179
rect 3065 3145 3099 3179
rect 3295 3145 3329 3179
rect 9321 3145 9355 3179
rect 19349 3145 19383 3179
rect 19901 3145 19935 3179
rect 22477 3145 22511 3179
rect 23121 3145 23155 3179
rect 3709 3077 3743 3111
rect 8677 3077 8711 3111
rect 10609 3077 10643 3111
rect 11897 3077 11931 3111
rect 13461 3077 13495 3111
rect 13921 3077 13955 3111
rect 25421 3077 25455 3111
rect 9045 3009 9079 3043
rect 10885 3009 10919 3043
rect 11529 3009 11563 3043
rect 12541 3009 12575 3043
rect 12817 3009 12851 3043
rect 15577 3009 15611 3043
rect 15669 3009 15703 3043
rect 15853 3009 15887 3043
rect 17233 3009 17267 3043
rect 18153 3009 18187 3043
rect 18429 3009 18463 3043
rect 21189 3009 21223 3043
rect 23765 3009 23799 3043
rect 24041 3009 24075 3043
rect 2212 2941 2246 2975
rect 3224 2941 3258 2975
rect 4204 2941 4238 2975
rect 5365 2941 5399 2975
rect 7573 2941 7607 2975
rect 8309 2941 8343 2975
rect 9505 2941 9539 2975
rect 9781 2941 9815 2975
rect 14105 2941 14139 2975
rect 16773 2941 16807 2975
rect 19625 2941 19659 2975
rect 19809 2941 19843 2975
rect 21833 2941 21867 2975
rect 25237 2941 25271 2975
rect 25789 2941 25823 2975
rect 2697 2873 2731 2907
rect 4629 2873 4663 2907
rect 5917 2873 5951 2907
rect 8401 2873 8435 2907
rect 10977 2873 11011 2907
rect 12173 2873 12207 2907
rect 12633 2873 12667 2907
rect 14467 2873 14501 2907
rect 15577 2873 15611 2907
rect 16174 2873 16208 2907
rect 17509 2873 17543 2907
rect 18245 2873 18279 2907
rect 20453 2873 20487 2907
rect 21281 2873 21315 2907
rect 22109 2873 22143 2907
rect 23857 2873 23891 2907
rect 4307 2805 4341 2839
rect 5089 2805 5123 2839
rect 6561 2805 6595 2839
rect 10241 2805 10275 2839
rect 15025 2805 15059 2839
rect 15301 2805 15335 2839
rect 20913 2805 20947 2839
rect 23397 2805 23431 2839
rect 24869 2805 24903 2839
rect 1547 2601 1581 2635
rect 2559 2601 2593 2635
rect 4399 2601 4433 2635
rect 7251 2601 7285 2635
rect 9321 2601 9355 2635
rect 9965 2601 9999 2635
rect 11161 2601 11195 2635
rect 11989 2601 12023 2635
rect 14105 2601 14139 2635
rect 16497 2601 16531 2635
rect 16957 2601 16991 2635
rect 17325 2601 17359 2635
rect 23765 2601 23799 2635
rect 10241 2533 10275 2567
rect 10333 2533 10367 2567
rect 10885 2533 10919 2567
rect 12817 2533 12851 2567
rect 15669 2533 15703 2567
rect 16221 2533 16255 2567
rect 18797 2533 18831 2567
rect 19349 2533 19383 2567
rect 21373 2533 21407 2567
rect 24133 2533 24167 2567
rect 24225 2533 24259 2567
rect 24777 2533 24811 2567
rect 1444 2465 1478 2499
rect 1869 2465 1903 2499
rect 2488 2465 2522 2499
rect 4328 2465 4362 2499
rect 5181 2465 5215 2499
rect 5917 2465 5951 2499
rect 7180 2465 7214 2499
rect 8033 2465 8067 2499
rect 8769 2465 8803 2499
rect 8861 2465 8895 2499
rect 13737 2465 13771 2499
rect 14289 2465 14323 2499
rect 17141 2465 17175 2499
rect 19625 2465 19659 2499
rect 22753 2465 22787 2499
rect 23489 2465 23523 2499
rect 25053 2465 25087 2499
rect 6009 2397 6043 2431
rect 11529 2397 11563 2431
rect 12725 2397 12759 2431
rect 13001 2397 13035 2431
rect 15209 2397 15243 2431
rect 15577 2397 15611 2431
rect 18705 2397 18739 2431
rect 19993 2397 20027 2431
rect 21281 2397 21315 2431
rect 21557 2397 21591 2431
rect 25605 2397 25639 2431
rect 7665 2329 7699 2363
rect 12357 2329 12391 2363
rect 14933 2329 14967 2363
rect 20545 2329 20579 2363
rect 2881 2261 2915 2295
rect 4813 2261 4847 2295
rect 14473 2261 14507 2295
rect 17693 2261 17727 2295
rect 18061 2261 18095 2295
rect 20913 2261 20947 2295
rect 22569 2261 22603 2295
rect 22937 2261 22971 2295
rect 25421 2261 25455 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 24762 24392 24768 24404
rect 24723 24364 24768 24392
rect 24762 24352 24768 24364
rect 24820 24352 24826 24404
rect 24581 24259 24639 24265
rect 24581 24225 24593 24259
rect 24627 24256 24639 24259
rect 25130 24256 25136 24268
rect 24627 24228 25136 24256
rect 24627 24225 24639 24228
rect 24581 24219 24639 24225
rect 25130 24216 25136 24228
rect 25188 24216 25194 24268
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 24765 23851 24823 23857
rect 24765 23817 24777 23851
rect 24811 23848 24823 23851
rect 24946 23848 24952 23860
rect 24811 23820 24952 23848
rect 24811 23817 24823 23820
rect 24765 23811 24823 23817
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 25130 23848 25136 23860
rect 25091 23820 25136 23848
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 24412 23616 24593 23644
rect 23658 23468 23664 23520
rect 23716 23508 23722 23520
rect 24412 23517 24440 23616
rect 24581 23613 24593 23616
rect 24627 23613 24639 23647
rect 24581 23607 24639 23613
rect 24397 23511 24455 23517
rect 24397 23508 24409 23511
rect 23716 23480 24409 23508
rect 23716 23468 23722 23480
rect 24397 23477 24409 23480
rect 24443 23477 24455 23511
rect 24397 23471 24455 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 24765 23307 24823 23313
rect 24765 23273 24777 23307
rect 24811 23304 24823 23307
rect 27614 23304 27620 23316
rect 24811 23276 27620 23304
rect 24811 23273 24823 23276
rect 24765 23267 24823 23273
rect 27614 23264 27620 23276
rect 27672 23264 27678 23316
rect 15562 23128 15568 23180
rect 15620 23168 15626 23180
rect 15692 23171 15750 23177
rect 15692 23168 15704 23171
rect 15620 23140 15704 23168
rect 15620 23128 15626 23140
rect 15692 23137 15704 23140
rect 15738 23137 15750 23171
rect 18966 23168 18972 23180
rect 18927 23140 18972 23168
rect 15692 23131 15750 23137
rect 18966 23128 18972 23140
rect 19024 23128 19030 23180
rect 24581 23171 24639 23177
rect 24581 23137 24593 23171
rect 24627 23168 24639 23171
rect 24670 23168 24676 23180
rect 24627 23140 24676 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 19199 23103 19257 23109
rect 19199 23069 19211 23103
rect 19245 23100 19257 23103
rect 20898 23100 20904 23112
rect 19245 23072 20904 23100
rect 19245 23069 19257 23072
rect 19199 23063 19257 23069
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 15795 22967 15853 22973
rect 15795 22933 15807 22967
rect 15841 22964 15853 22967
rect 23290 22964 23296 22976
rect 15841 22936 23296 22964
rect 15841 22933 15853 22936
rect 15795 22927 15853 22933
rect 23290 22924 23296 22936
rect 23348 22924 23354 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 15562 22380 15568 22432
rect 15620 22420 15626 22432
rect 15657 22423 15715 22429
rect 15657 22420 15669 22423
rect 15620 22392 15669 22420
rect 15620 22380 15626 22392
rect 15657 22389 15669 22392
rect 15703 22389 15715 22423
rect 15657 22383 15715 22389
rect 18322 22380 18328 22432
rect 18380 22420 18386 22432
rect 18966 22420 18972 22432
rect 18380 22392 18972 22420
rect 18380 22380 18386 22392
rect 18966 22380 18972 22392
rect 19024 22420 19030 22432
rect 19061 22423 19119 22429
rect 19061 22420 19073 22423
rect 19024 22392 19073 22420
rect 19024 22380 19030 22392
rect 19061 22389 19073 22392
rect 19107 22389 19119 22423
rect 24578 22420 24584 22432
rect 24539 22392 24584 22420
rect 19061 22383 19119 22389
rect 24578 22380 24584 22392
rect 24636 22380 24642 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 24765 21675 24823 21681
rect 24765 21641 24777 21675
rect 24811 21672 24823 21675
rect 24854 21672 24860 21684
rect 24811 21644 24860 21672
rect 24811 21641 24823 21644
rect 24765 21635 24823 21641
rect 24854 21632 24860 21644
rect 24912 21632 24918 21684
rect 24581 21471 24639 21477
rect 24581 21437 24593 21471
rect 24627 21468 24639 21471
rect 24627 21440 25268 21468
rect 24627 21437 24639 21440
rect 24581 21431 24639 21437
rect 25240 21341 25268 21440
rect 25225 21335 25283 21341
rect 25225 21301 25237 21335
rect 25271 21332 25283 21335
rect 25314 21332 25320 21344
rect 25271 21304 25320 21332
rect 25271 21301 25283 21304
rect 25225 21295 25283 21301
rect 25314 21292 25320 21304
rect 25372 21292 25378 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 24762 21128 24768 21140
rect 24723 21100 24768 21128
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 24581 20995 24639 21001
rect 24581 20961 24593 20995
rect 24627 20992 24639 20995
rect 24670 20992 24676 21004
rect 24627 20964 24676 20992
rect 24627 20961 24639 20964
rect 24581 20955 24639 20961
rect 24670 20952 24676 20964
rect 24728 20952 24734 21004
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 24351 20519 24409 20525
rect 24351 20485 24363 20519
rect 24397 20516 24409 20519
rect 24670 20516 24676 20528
rect 24397 20488 24676 20516
rect 24397 20485 24409 20488
rect 24351 20479 24409 20485
rect 24670 20476 24676 20488
rect 24728 20516 24734 20528
rect 25041 20519 25099 20525
rect 25041 20516 25053 20519
rect 24728 20488 25053 20516
rect 24728 20476 24734 20488
rect 25041 20485 25053 20488
rect 25087 20485 25099 20519
rect 25041 20479 25099 20485
rect 24280 20383 24338 20389
rect 24280 20349 24292 20383
rect 24326 20380 24338 20383
rect 24326 20352 24808 20380
rect 24326 20349 24338 20352
rect 24280 20343 24338 20349
rect 24780 20253 24808 20352
rect 24765 20247 24823 20253
rect 24765 20213 24777 20247
rect 24811 20244 24823 20247
rect 24946 20244 24952 20256
rect 24811 20216 24952 20244
rect 24811 20213 24823 20216
rect 24765 20207 24823 20213
rect 24946 20204 24952 20216
rect 25004 20204 25010 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 24762 20040 24768 20052
rect 24723 20012 24768 20040
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 24581 19907 24639 19913
rect 24581 19873 24593 19907
rect 24627 19904 24639 19907
rect 24670 19904 24676 19916
rect 24627 19876 24676 19904
rect 24627 19873 24639 19876
rect 24581 19867 24639 19873
rect 24670 19864 24676 19876
rect 24728 19864 24734 19916
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 24535 19431 24593 19437
rect 24535 19397 24547 19431
rect 24581 19428 24593 19431
rect 24670 19428 24676 19440
rect 24581 19400 24676 19428
rect 24581 19397 24593 19400
rect 24535 19391 24593 19397
rect 24670 19388 24676 19400
rect 24728 19428 24734 19440
rect 25225 19431 25283 19437
rect 25225 19428 25237 19431
rect 24728 19400 25237 19428
rect 24728 19388 24734 19400
rect 25225 19397 25237 19400
rect 25271 19397 25283 19431
rect 25225 19391 25283 19397
rect 24464 19295 24522 19301
rect 24464 19261 24476 19295
rect 24510 19292 24522 19295
rect 24510 19264 24900 19292
rect 24510 19261 24522 19264
rect 24464 19255 24522 19261
rect 24872 19168 24900 19264
rect 24854 19156 24860 19168
rect 24815 19128 24860 19156
rect 24854 19116 24860 19128
rect 24912 19116 24918 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 24762 18952 24768 18964
rect 24723 18924 24768 18952
rect 24762 18912 24768 18924
rect 24820 18912 24826 18964
rect 23566 18816 23572 18828
rect 23527 18788 23572 18816
rect 23566 18776 23572 18788
rect 23624 18776 23630 18828
rect 24581 18819 24639 18825
rect 24581 18785 24593 18819
rect 24627 18816 24639 18819
rect 24670 18816 24676 18828
rect 24627 18788 24676 18816
rect 24627 18785 24639 18788
rect 24581 18779 24639 18785
rect 24670 18776 24676 18788
rect 24728 18776 24734 18828
rect 22557 18751 22615 18757
rect 22557 18717 22569 18751
rect 22603 18748 22615 18751
rect 23750 18748 23756 18760
rect 22603 18720 23756 18748
rect 22603 18717 22615 18720
rect 22557 18711 22615 18717
rect 23750 18708 23756 18720
rect 23808 18708 23814 18760
rect 23707 18615 23765 18621
rect 23707 18581 23719 18615
rect 23753 18612 23765 18615
rect 25222 18612 25228 18624
rect 23753 18584 25228 18612
rect 23753 18581 23765 18584
rect 23707 18575 23765 18581
rect 25222 18572 25228 18584
rect 25280 18572 25286 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 24489 18411 24547 18417
rect 24489 18408 24501 18411
rect 23446 18380 24501 18408
rect 22695 18343 22753 18349
rect 22695 18309 22707 18343
rect 22741 18340 22753 18343
rect 23446 18340 23474 18380
rect 24489 18377 24501 18380
rect 24535 18408 24547 18411
rect 24670 18408 24676 18420
rect 24535 18380 24676 18408
rect 24535 18377 24547 18380
rect 24489 18371 24547 18377
rect 24670 18368 24676 18380
rect 24728 18368 24734 18420
rect 22741 18312 23474 18340
rect 22741 18309 22753 18312
rect 22695 18303 22753 18309
rect 24118 18300 24124 18352
rect 24176 18340 24182 18352
rect 24765 18343 24823 18349
rect 24765 18340 24777 18343
rect 24176 18312 24777 18340
rect 24176 18300 24182 18312
rect 24765 18309 24777 18312
rect 24811 18309 24823 18343
rect 24765 18303 24823 18309
rect 22624 18207 22682 18213
rect 22624 18173 22636 18207
rect 22670 18204 22682 18207
rect 23109 18207 23167 18213
rect 23109 18204 23121 18207
rect 22670 18176 23121 18204
rect 22670 18173 22682 18176
rect 22624 18167 22682 18173
rect 23109 18173 23121 18176
rect 23155 18204 23167 18207
rect 23934 18204 23940 18216
rect 23155 18176 23940 18204
rect 23155 18173 23167 18176
rect 23109 18167 23167 18173
rect 23934 18164 23940 18176
rect 23992 18164 23998 18216
rect 24210 18164 24216 18216
rect 24268 18204 24274 18216
rect 24581 18207 24639 18213
rect 24581 18204 24593 18207
rect 24268 18176 24593 18204
rect 24268 18164 24274 18176
rect 24581 18173 24593 18176
rect 24627 18204 24639 18207
rect 25133 18207 25191 18213
rect 25133 18204 25145 18207
rect 24627 18176 25145 18204
rect 24627 18173 24639 18176
rect 24581 18167 24639 18173
rect 25133 18173 25145 18176
rect 25179 18173 25191 18207
rect 25133 18167 25191 18173
rect 21545 18071 21603 18077
rect 21545 18037 21557 18071
rect 21591 18068 21603 18071
rect 22094 18068 22100 18080
rect 21591 18040 22100 18068
rect 21591 18037 21603 18040
rect 21545 18031 21603 18037
rect 22094 18028 22100 18040
rect 22152 18028 22158 18080
rect 23566 18028 23572 18080
rect 23624 18068 23630 18080
rect 23937 18071 23995 18077
rect 23937 18068 23949 18071
rect 23624 18040 23949 18068
rect 23624 18028 23630 18040
rect 23937 18037 23949 18040
rect 23983 18068 23995 18071
rect 25498 18068 25504 18080
rect 23983 18040 25504 18068
rect 23983 18037 23995 18040
rect 23937 18031 23995 18037
rect 25498 18028 25504 18040
rect 25556 18028 25562 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 16390 17864 16396 17876
rect 16351 17836 16396 17864
rect 16390 17824 16396 17836
rect 16448 17824 16454 17876
rect 16114 17728 16120 17740
rect 16075 17700 16120 17728
rect 16114 17688 16120 17700
rect 16172 17688 16178 17740
rect 17770 17728 17776 17740
rect 17731 17700 17776 17728
rect 17770 17688 17776 17700
rect 17828 17688 17834 17740
rect 21542 17728 21548 17740
rect 21503 17700 21548 17728
rect 21542 17688 21548 17700
rect 21600 17688 21606 17740
rect 22830 17728 22836 17740
rect 22791 17700 22836 17728
rect 22830 17688 22836 17700
rect 22888 17688 22894 17740
rect 24857 17731 24915 17737
rect 24857 17697 24869 17731
rect 24903 17728 24915 17731
rect 25038 17728 25044 17740
rect 24903 17700 25044 17728
rect 24903 17697 24915 17700
rect 24857 17691 24915 17697
rect 25038 17688 25044 17700
rect 25096 17688 25102 17740
rect 21818 17660 21824 17672
rect 21779 17632 21824 17660
rect 21818 17620 21824 17632
rect 21876 17620 21882 17672
rect 23842 17620 23848 17672
rect 23900 17660 23906 17672
rect 24213 17663 24271 17669
rect 24213 17660 24225 17663
rect 23900 17632 24225 17660
rect 23900 17620 23906 17632
rect 24213 17629 24225 17632
rect 24259 17629 24271 17663
rect 24213 17623 24271 17629
rect 18138 17524 18144 17536
rect 18099 17496 18144 17524
rect 18138 17484 18144 17496
rect 18196 17484 18202 17536
rect 23109 17527 23167 17533
rect 23109 17493 23121 17527
rect 23155 17524 23167 17527
rect 23290 17524 23296 17536
rect 23155 17496 23296 17524
rect 23155 17493 23167 17496
rect 23109 17487 23167 17493
rect 23290 17484 23296 17496
rect 23348 17484 23354 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 15933 17323 15991 17329
rect 15933 17289 15945 17323
rect 15979 17320 15991 17323
rect 16114 17320 16120 17332
rect 15979 17292 16120 17320
rect 15979 17289 15991 17292
rect 15933 17283 15991 17289
rect 16114 17280 16120 17292
rect 16172 17280 16178 17332
rect 17770 17320 17776 17332
rect 17731 17292 17776 17320
rect 17770 17280 17776 17292
rect 17828 17280 17834 17332
rect 21542 17320 21548 17332
rect 21503 17292 21548 17320
rect 21542 17280 21548 17292
rect 21600 17320 21606 17332
rect 21910 17320 21916 17332
rect 21600 17292 21916 17320
rect 21600 17280 21606 17292
rect 21910 17280 21916 17292
rect 21968 17280 21974 17332
rect 24765 17323 24823 17329
rect 24765 17289 24777 17323
rect 24811 17320 24823 17323
rect 25038 17320 25044 17332
rect 24811 17292 25044 17320
rect 24811 17289 24823 17292
rect 24765 17283 24823 17289
rect 25038 17280 25044 17292
rect 25096 17280 25102 17332
rect 25406 17320 25412 17332
rect 25367 17292 25412 17320
rect 25406 17280 25412 17292
rect 25464 17280 25470 17332
rect 14737 17119 14795 17125
rect 14737 17085 14749 17119
rect 14783 17116 14795 17119
rect 14921 17119 14979 17125
rect 14921 17116 14933 17119
rect 14783 17088 14933 17116
rect 14783 17085 14795 17088
rect 14737 17079 14795 17085
rect 14921 17085 14933 17088
rect 14967 17116 14979 17119
rect 15470 17116 15476 17128
rect 14967 17088 15476 17116
rect 14967 17085 14979 17088
rect 14921 17079 14979 17085
rect 15470 17076 15476 17088
rect 15528 17076 15534 17128
rect 16301 17119 16359 17125
rect 16301 17085 16313 17119
rect 16347 17116 16359 17119
rect 16485 17119 16543 17125
rect 16485 17116 16497 17119
rect 16347 17088 16497 17116
rect 16347 17085 16359 17088
rect 16301 17079 16359 17085
rect 16485 17085 16497 17088
rect 16531 17116 16543 17119
rect 17034 17116 17040 17128
rect 16531 17088 17040 17116
rect 16531 17085 16543 17088
rect 16485 17079 16543 17085
rect 17034 17076 17040 17088
rect 17092 17076 17098 17128
rect 18693 17119 18751 17125
rect 18693 17085 18705 17119
rect 18739 17116 18751 17119
rect 18877 17119 18935 17125
rect 18877 17116 18889 17119
rect 18739 17088 18889 17116
rect 18739 17085 18751 17088
rect 18693 17079 18751 17085
rect 18877 17085 18889 17088
rect 18923 17116 18935 17119
rect 18966 17116 18972 17128
rect 18923 17088 18972 17116
rect 18923 17085 18935 17088
rect 18877 17079 18935 17085
rect 18966 17076 18972 17088
rect 19024 17076 19030 17128
rect 20349 17119 20407 17125
rect 20349 17085 20361 17119
rect 20395 17116 20407 17119
rect 20533 17119 20591 17125
rect 20533 17116 20545 17119
rect 20395 17088 20545 17116
rect 20395 17085 20407 17088
rect 20349 17079 20407 17085
rect 20533 17085 20545 17088
rect 20579 17116 20591 17119
rect 20806 17116 20812 17128
rect 20579 17088 20812 17116
rect 20579 17085 20591 17088
rect 20533 17079 20591 17085
rect 20806 17076 20812 17088
rect 20864 17076 20870 17128
rect 21913 17119 21971 17125
rect 21913 17085 21925 17119
rect 21959 17116 21971 17119
rect 22002 17116 22008 17128
rect 21959 17088 22008 17116
rect 21959 17085 21971 17088
rect 21913 17079 21971 17085
rect 22002 17076 22008 17088
rect 22060 17116 22066 17128
rect 22097 17119 22155 17125
rect 22097 17116 22109 17119
rect 22060 17088 22109 17116
rect 22060 17076 22066 17088
rect 22097 17085 22109 17088
rect 22143 17085 22155 17119
rect 22097 17079 22155 17085
rect 23198 17076 23204 17128
rect 23256 17116 23262 17128
rect 23385 17119 23443 17125
rect 23385 17116 23397 17119
rect 23256 17088 23397 17116
rect 23256 17076 23262 17088
rect 23385 17085 23397 17088
rect 23431 17116 23443 17119
rect 23753 17119 23811 17125
rect 23753 17116 23765 17119
rect 23431 17088 23765 17116
rect 23431 17085 23443 17088
rect 23385 17079 23443 17085
rect 23753 17085 23765 17088
rect 23799 17085 23811 17119
rect 25222 17116 25228 17128
rect 25183 17088 25228 17116
rect 23753 17079 23811 17085
rect 25222 17076 25228 17088
rect 25280 17116 25286 17128
rect 25777 17119 25835 17125
rect 25777 17116 25789 17119
rect 25280 17088 25789 17116
rect 25280 17076 25286 17088
rect 25777 17085 25789 17088
rect 25823 17085 25835 17119
rect 25777 17079 25835 17085
rect 16390 17048 16396 17060
rect 16351 17020 16396 17048
rect 16390 17008 16396 17020
rect 16448 17008 16454 17060
rect 22738 17048 22744 17060
rect 22699 17020 22744 17048
rect 22738 17008 22744 17020
rect 22796 17008 22802 17060
rect 23474 17008 23480 17060
rect 23532 17048 23538 17060
rect 23661 17051 23719 17057
rect 23661 17048 23673 17051
rect 23532 17020 23673 17048
rect 23532 17008 23538 17020
rect 23661 17017 23673 17020
rect 23707 17017 23719 17051
rect 23661 17011 23719 17017
rect 15286 16980 15292 16992
rect 15247 16952 15292 16980
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 19058 16980 19064 16992
rect 19019 16952 19064 16980
rect 19058 16940 19064 16952
rect 19116 16940 19122 16992
rect 20714 16980 20720 16992
rect 20675 16952 20720 16980
rect 20714 16940 20720 16952
rect 20772 16940 20778 16992
rect 22186 16940 22192 16992
rect 22244 16980 22250 16992
rect 22830 16980 22836 16992
rect 22244 16952 22836 16980
rect 22244 16940 22250 16952
rect 22830 16940 22836 16952
rect 22888 16980 22894 16992
rect 23017 16983 23075 16989
rect 23017 16980 23029 16983
rect 22888 16952 23029 16980
rect 22888 16940 22894 16952
rect 23017 16949 23029 16952
rect 23063 16949 23075 16983
rect 23017 16943 23075 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 19935 16779 19993 16785
rect 19935 16745 19947 16779
rect 19981 16776 19993 16779
rect 24210 16776 24216 16788
rect 19981 16748 24216 16776
rect 19981 16745 19993 16748
rect 19935 16739 19993 16745
rect 24210 16736 24216 16748
rect 24268 16736 24274 16788
rect 15473 16711 15531 16717
rect 15473 16677 15485 16711
rect 15519 16708 15531 16711
rect 16206 16708 16212 16720
rect 15519 16680 16212 16708
rect 15519 16677 15531 16680
rect 15473 16671 15531 16677
rect 16206 16668 16212 16680
rect 16264 16668 16270 16720
rect 18138 16668 18144 16720
rect 18196 16708 18202 16720
rect 18233 16711 18291 16717
rect 18233 16708 18245 16711
rect 18196 16680 18245 16708
rect 18196 16668 18202 16680
rect 18233 16677 18245 16680
rect 18279 16677 18291 16711
rect 18233 16671 18291 16677
rect 19518 16600 19524 16652
rect 19576 16640 19582 16652
rect 19832 16643 19890 16649
rect 19832 16640 19844 16643
rect 19576 16612 19844 16640
rect 19576 16600 19582 16612
rect 19832 16609 19844 16612
rect 19878 16609 19890 16643
rect 21634 16640 21640 16652
rect 21595 16612 21640 16640
rect 19832 16603 19890 16609
rect 21634 16600 21640 16612
rect 21692 16600 21698 16652
rect 22554 16600 22560 16652
rect 22612 16640 22618 16652
rect 23109 16643 23167 16649
rect 23109 16640 23121 16643
rect 22612 16612 23121 16640
rect 22612 16600 22618 16612
rect 23109 16609 23121 16612
rect 23155 16609 23167 16643
rect 23382 16640 23388 16652
rect 23343 16612 23388 16640
rect 23109 16603 23167 16609
rect 23382 16600 23388 16612
rect 23440 16600 23446 16652
rect 25038 16640 25044 16652
rect 24999 16612 25044 16640
rect 25038 16600 25044 16612
rect 25096 16600 25102 16652
rect 15381 16575 15439 16581
rect 15381 16541 15393 16575
rect 15427 16541 15439 16575
rect 15654 16572 15660 16584
rect 15615 16544 15660 16572
rect 15381 16535 15439 16541
rect 15396 16504 15424 16535
rect 15654 16532 15660 16544
rect 15712 16532 15718 16584
rect 18138 16572 18144 16584
rect 18099 16544 18144 16572
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 18322 16532 18328 16584
rect 18380 16572 18386 16584
rect 18417 16575 18475 16581
rect 18417 16572 18429 16575
rect 18380 16544 18429 16572
rect 18380 16532 18386 16544
rect 18417 16541 18429 16544
rect 18463 16541 18475 16575
rect 18417 16535 18475 16541
rect 22281 16575 22339 16581
rect 22281 16541 22293 16575
rect 22327 16572 22339 16575
rect 22646 16572 22652 16584
rect 22327 16544 22652 16572
rect 22327 16541 22339 16544
rect 22281 16535 22339 16541
rect 22646 16532 22652 16544
rect 22704 16532 22710 16584
rect 24118 16532 24124 16584
rect 24176 16572 24182 16584
rect 24673 16575 24731 16581
rect 24673 16572 24685 16575
rect 24176 16544 24685 16572
rect 24176 16532 24182 16544
rect 24673 16541 24685 16544
rect 24719 16541 24731 16575
rect 24673 16535 24731 16541
rect 16666 16504 16672 16516
rect 15396 16476 16672 16504
rect 16666 16464 16672 16476
rect 16724 16464 16730 16516
rect 19242 16436 19248 16448
rect 19203 16408 19248 16436
rect 19242 16396 19248 16408
rect 19300 16396 19306 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 15105 16235 15163 16241
rect 15105 16201 15117 16235
rect 15151 16232 15163 16235
rect 15286 16232 15292 16244
rect 15151 16204 15292 16232
rect 15151 16201 15163 16204
rect 15105 16195 15163 16201
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 18230 16192 18236 16244
rect 18288 16232 18294 16244
rect 18509 16235 18567 16241
rect 18509 16232 18521 16235
rect 18288 16204 18521 16232
rect 18288 16192 18294 16204
rect 18509 16201 18521 16204
rect 18555 16201 18567 16235
rect 19058 16232 19064 16244
rect 19019 16204 19064 16232
rect 18509 16195 18567 16201
rect 19058 16192 19064 16204
rect 19116 16192 19122 16244
rect 21542 16232 21548 16244
rect 21503 16204 21548 16232
rect 21542 16192 21548 16204
rect 21600 16192 21606 16244
rect 21818 16232 21824 16244
rect 21779 16204 21824 16232
rect 21818 16192 21824 16204
rect 21876 16192 21882 16244
rect 25314 16192 25320 16244
rect 25372 16232 25378 16244
rect 25731 16235 25789 16241
rect 25731 16232 25743 16235
rect 25372 16204 25743 16232
rect 25372 16192 25378 16204
rect 25731 16201 25743 16204
rect 25777 16201 25789 16235
rect 25731 16195 25789 16201
rect 23017 16167 23075 16173
rect 23017 16164 23029 16167
rect 22112 16136 23029 16164
rect 22112 16108 22140 16136
rect 23017 16133 23029 16136
rect 23063 16133 23075 16167
rect 23017 16127 23075 16133
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16096 15991 16099
rect 16114 16096 16120 16108
rect 15979 16068 16120 16096
rect 15979 16065 15991 16068
rect 15933 16059 15991 16065
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 17865 16099 17923 16105
rect 17865 16065 17877 16099
rect 17911 16096 17923 16099
rect 18049 16099 18107 16105
rect 18049 16096 18061 16099
rect 17911 16068 18061 16096
rect 17911 16065 17923 16068
rect 17865 16059 17923 16065
rect 18049 16065 18061 16068
rect 18095 16096 18107 16099
rect 18138 16096 18144 16108
rect 18095 16068 18144 16096
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 18138 16056 18144 16068
rect 18196 16056 18202 16108
rect 19242 16096 19248 16108
rect 19203 16068 19248 16096
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 19518 16096 19524 16108
rect 19479 16068 19524 16096
rect 19518 16056 19524 16068
rect 19576 16096 19582 16108
rect 20165 16099 20223 16105
rect 20165 16096 20177 16099
rect 19576 16068 20177 16096
rect 19576 16056 19582 16068
rect 20165 16065 20177 16068
rect 20211 16065 20223 16099
rect 22094 16096 22100 16108
rect 22055 16068 22100 16096
rect 20165 16059 20223 16065
rect 22094 16056 22100 16068
rect 22152 16056 22158 16108
rect 22462 16096 22468 16108
rect 22423 16068 22468 16096
rect 22462 16056 22468 16068
rect 22520 16096 22526 16108
rect 22520 16068 25671 16096
rect 22520 16056 22526 16068
rect 21060 16031 21118 16037
rect 21060 15997 21072 16031
rect 21106 16028 21118 16031
rect 21542 16028 21548 16040
rect 21106 16000 21548 16028
rect 21106 15997 21118 16000
rect 21060 15991 21118 15997
rect 21542 15988 21548 16000
rect 21600 15988 21606 16040
rect 25643 16037 25671 16068
rect 23937 16031 23995 16037
rect 23937 16028 23949 16031
rect 23446 16000 23949 16028
rect 14185 15963 14243 15969
rect 14185 15929 14197 15963
rect 14231 15960 14243 15963
rect 14737 15963 14795 15969
rect 14737 15960 14749 15963
rect 14231 15932 14749 15960
rect 14231 15929 14243 15932
rect 14185 15923 14243 15929
rect 14737 15929 14749 15932
rect 14783 15960 14795 15963
rect 15289 15963 15347 15969
rect 15289 15960 15301 15963
rect 14783 15932 15301 15960
rect 14783 15929 14795 15932
rect 14737 15923 14795 15929
rect 15289 15929 15301 15932
rect 15335 15929 15347 15963
rect 15289 15923 15347 15929
rect 15378 15920 15384 15972
rect 15436 15960 15442 15972
rect 19337 15963 19395 15969
rect 15436 15932 15481 15960
rect 15436 15920 15442 15932
rect 19337 15929 19349 15963
rect 19383 15929 19395 15963
rect 19337 15923 19395 15929
rect 22189 15963 22247 15969
rect 22189 15929 22201 15963
rect 22235 15929 22247 15963
rect 22189 15923 22247 15929
rect 16206 15892 16212 15904
rect 16167 15864 16212 15892
rect 16206 15852 16212 15864
rect 16264 15852 16270 15904
rect 16666 15892 16672 15904
rect 16627 15864 16672 15892
rect 16666 15852 16672 15864
rect 16724 15852 16730 15904
rect 19058 15852 19064 15904
rect 19116 15892 19122 15904
rect 19352 15892 19380 15923
rect 19116 15864 19380 15892
rect 19116 15852 19122 15864
rect 19426 15852 19432 15904
rect 19484 15892 19490 15904
rect 21131 15895 21189 15901
rect 21131 15892 21143 15895
rect 19484 15864 21143 15892
rect 19484 15852 19490 15864
rect 21131 15861 21143 15864
rect 21177 15861 21189 15895
rect 21131 15855 21189 15861
rect 21818 15852 21824 15904
rect 21876 15892 21882 15904
rect 22204 15892 22232 15923
rect 22922 15920 22928 15972
rect 22980 15960 22986 15972
rect 23446 15960 23474 16000
rect 23937 15997 23949 16000
rect 23983 16028 23995 16031
rect 24121 16031 24179 16037
rect 24121 16028 24133 16031
rect 23983 16000 24133 16028
rect 23983 15997 23995 16000
rect 23937 15991 23995 15997
rect 24121 15997 24133 16000
rect 24167 15997 24179 16031
rect 24121 15991 24179 15997
rect 25628 16031 25686 16037
rect 25628 15997 25640 16031
rect 25674 16028 25686 16031
rect 26053 16031 26111 16037
rect 26053 16028 26065 16031
rect 25674 16000 26065 16028
rect 25674 15997 25686 16000
rect 25628 15991 25686 15997
rect 26053 15997 26065 16000
rect 26099 15997 26111 16031
rect 26053 15991 26111 15997
rect 22980 15932 23474 15960
rect 24765 15963 24823 15969
rect 22980 15920 22986 15932
rect 24765 15929 24777 15963
rect 24811 15960 24823 15963
rect 24946 15960 24952 15972
rect 24811 15932 24952 15960
rect 24811 15929 24823 15932
rect 24765 15923 24823 15929
rect 24946 15920 24952 15932
rect 25004 15920 25010 15972
rect 21876 15864 22232 15892
rect 21876 15852 21882 15864
rect 22278 15852 22284 15904
rect 22336 15892 22342 15904
rect 23382 15892 23388 15904
rect 22336 15864 23388 15892
rect 22336 15852 22342 15864
rect 23382 15852 23388 15864
rect 23440 15852 23446 15904
rect 25038 15892 25044 15904
rect 24999 15864 25044 15892
rect 25038 15852 25044 15864
rect 25096 15852 25102 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 18138 15648 18144 15700
rect 18196 15688 18202 15700
rect 18417 15691 18475 15697
rect 18417 15688 18429 15691
rect 18196 15660 18429 15688
rect 18196 15648 18202 15660
rect 18417 15657 18429 15660
rect 18463 15688 18475 15691
rect 19426 15688 19432 15700
rect 18463 15660 19432 15688
rect 18463 15657 18475 15660
rect 18417 15651 18475 15657
rect 19426 15648 19432 15660
rect 19484 15648 19490 15700
rect 21634 15688 21640 15700
rect 21595 15660 21640 15688
rect 21634 15648 21640 15660
rect 21692 15648 21698 15700
rect 13814 15580 13820 15632
rect 13872 15620 13878 15632
rect 15470 15620 15476 15632
rect 13872 15592 13917 15620
rect 15431 15592 15476 15620
rect 13872 15580 13878 15592
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 16025 15623 16083 15629
rect 16025 15589 16037 15623
rect 16071 15620 16083 15623
rect 16114 15620 16120 15632
rect 16071 15592 16120 15620
rect 16071 15589 16083 15592
rect 16025 15583 16083 15589
rect 16114 15580 16120 15592
rect 16172 15580 16178 15632
rect 17497 15623 17555 15629
rect 17497 15589 17509 15623
rect 17543 15620 17555 15623
rect 17770 15620 17776 15632
rect 17543 15592 17776 15620
rect 17543 15589 17555 15592
rect 17497 15583 17555 15589
rect 17770 15580 17776 15592
rect 17828 15580 17834 15632
rect 18049 15623 18107 15629
rect 18049 15589 18061 15623
rect 18095 15620 18107 15623
rect 18322 15620 18328 15632
rect 18095 15592 18328 15620
rect 18095 15589 18107 15592
rect 18049 15583 18107 15589
rect 18322 15580 18328 15592
rect 18380 15580 18386 15632
rect 18966 15580 18972 15632
rect 19024 15620 19030 15632
rect 19061 15623 19119 15629
rect 19061 15620 19073 15623
rect 19024 15592 19073 15620
rect 19024 15580 19030 15592
rect 19061 15589 19073 15592
rect 19107 15589 19119 15623
rect 21910 15620 21916 15632
rect 21871 15592 21916 15620
rect 19061 15583 19119 15589
rect 21910 15580 21916 15592
rect 21968 15580 21974 15632
rect 22462 15620 22468 15632
rect 22423 15592 22468 15620
rect 22462 15580 22468 15592
rect 22520 15580 22526 15632
rect 24210 15552 24216 15564
rect 24171 15524 24216 15552
rect 24210 15512 24216 15524
rect 24268 15512 24274 15564
rect 13722 15484 13728 15496
rect 13683 15456 13728 15484
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 14369 15487 14427 15493
rect 14369 15453 14381 15487
rect 14415 15484 14427 15487
rect 15381 15487 15439 15493
rect 15381 15484 15393 15487
rect 14415 15456 15393 15484
rect 14415 15453 14427 15456
rect 14369 15447 14427 15453
rect 15381 15453 15393 15456
rect 15427 15484 15439 15487
rect 15654 15484 15660 15496
rect 15427 15456 15660 15484
rect 15427 15453 15439 15456
rect 15381 15447 15439 15453
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 17402 15484 17408 15496
rect 17363 15456 17408 15484
rect 17402 15444 17408 15456
rect 17460 15444 17466 15496
rect 18969 15487 19027 15493
rect 18969 15453 18981 15487
rect 19015 15484 19027 15487
rect 19426 15484 19432 15496
rect 19015 15456 19432 15484
rect 19015 15453 19027 15456
rect 18969 15447 19027 15453
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 21818 15484 21824 15496
rect 21779 15456 21824 15484
rect 21818 15444 21824 15456
rect 21876 15444 21882 15496
rect 24762 15484 24768 15496
rect 24723 15456 24768 15484
rect 24762 15444 24768 15456
rect 24820 15444 24826 15496
rect 19518 15416 19524 15428
rect 19479 15388 19524 15416
rect 19518 15376 19524 15388
rect 19576 15376 19582 15428
rect 16482 15348 16488 15360
rect 16443 15320 16488 15348
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 13814 15144 13820 15156
rect 13786 15104 13820 15144
rect 13872 15144 13878 15156
rect 15289 15147 15347 15153
rect 13872 15116 13917 15144
rect 13872 15104 13878 15116
rect 15289 15113 15301 15147
rect 15335 15144 15347 15147
rect 15470 15144 15476 15156
rect 15335 15116 15476 15144
rect 15335 15113 15347 15116
rect 15289 15107 15347 15113
rect 15470 15104 15476 15116
rect 15528 15144 15534 15156
rect 15565 15147 15623 15153
rect 15565 15144 15577 15147
rect 15528 15116 15577 15144
rect 15528 15104 15534 15116
rect 15565 15113 15577 15116
rect 15611 15113 15623 15147
rect 15565 15107 15623 15113
rect 16301 15147 16359 15153
rect 16301 15113 16313 15147
rect 16347 15144 16359 15147
rect 16390 15144 16396 15156
rect 16347 15116 16396 15144
rect 16347 15113 16359 15116
rect 16301 15107 16359 15113
rect 16390 15104 16396 15116
rect 16448 15104 16454 15156
rect 17497 15147 17555 15153
rect 17497 15113 17509 15147
rect 17543 15144 17555 15147
rect 17770 15144 17776 15156
rect 17543 15116 17776 15144
rect 17543 15113 17555 15116
rect 17497 15107 17555 15113
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 18966 15104 18972 15156
rect 19024 15144 19030 15156
rect 19061 15147 19119 15153
rect 19061 15144 19073 15147
rect 19024 15116 19073 15144
rect 19024 15104 19030 15116
rect 19061 15113 19073 15116
rect 19107 15113 19119 15147
rect 19061 15107 19119 15113
rect 20625 15147 20683 15153
rect 20625 15113 20637 15147
rect 20671 15144 20683 15147
rect 20714 15144 20720 15156
rect 20671 15116 20720 15144
rect 20671 15113 20683 15116
rect 20625 15107 20683 15113
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 21821 15147 21879 15153
rect 21821 15113 21833 15147
rect 21867 15144 21879 15147
rect 21910 15144 21916 15156
rect 21867 15116 21916 15144
rect 21867 15113 21879 15116
rect 21821 15107 21879 15113
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 23106 15144 23112 15156
rect 23067 15116 23112 15144
rect 23106 15104 23112 15116
rect 23164 15104 23170 15156
rect 23658 15104 23664 15156
rect 23716 15144 23722 15156
rect 24210 15144 24216 15156
rect 23716 15116 24216 15144
rect 23716 15104 23722 15116
rect 24210 15104 24216 15116
rect 24268 15144 24274 15156
rect 24673 15147 24731 15153
rect 24673 15144 24685 15147
rect 24268 15116 24685 15144
rect 24268 15104 24274 15116
rect 24673 15113 24685 15116
rect 24719 15113 24731 15147
rect 25774 15144 25780 15156
rect 25735 15116 25780 15144
rect 24673 15107 24731 15113
rect 25774 15104 25780 15116
rect 25832 15104 25838 15156
rect 13541 15011 13599 15017
rect 13541 14977 13553 15011
rect 13587 15008 13599 15011
rect 13786 15008 13814 15104
rect 24302 15036 24308 15088
rect 24360 15076 24366 15088
rect 25363 15079 25421 15085
rect 25363 15076 25375 15079
rect 24360 15048 25375 15076
rect 24360 15036 24366 15048
rect 25363 15045 25375 15048
rect 25409 15045 25421 15079
rect 25363 15039 25421 15045
rect 13587 14980 13814 15008
rect 17129 15011 17187 15017
rect 13587 14977 13599 14980
rect 13541 14971 13599 14977
rect 17129 14977 17141 15011
rect 17175 15008 17187 15011
rect 17402 15008 17408 15020
rect 17175 14980 17408 15008
rect 17175 14977 17187 14980
rect 17129 14971 17187 14977
rect 17402 14968 17408 14980
rect 17460 15008 17466 15020
rect 18417 15011 18475 15017
rect 18417 15008 18429 15011
rect 17460 14980 18429 15008
rect 17460 14968 17466 14980
rect 18417 14977 18429 14980
rect 18463 14977 18475 15011
rect 18417 14971 18475 14977
rect 19242 14968 19248 15020
rect 19300 15008 19306 15020
rect 19613 15011 19671 15017
rect 19613 15008 19625 15011
rect 19300 14980 19625 15008
rect 19300 14968 19306 14980
rect 19613 14977 19625 14980
rect 19659 14977 19671 15011
rect 23750 15008 23756 15020
rect 23711 14980 23756 15008
rect 19613 14971 19671 14977
rect 23750 14968 23756 14980
rect 23808 14968 23814 15020
rect 12713 14943 12771 14949
rect 12713 14909 12725 14943
rect 12759 14940 12771 14943
rect 13446 14940 13452 14952
rect 12759 14912 13452 14940
rect 12759 14909 12771 14912
rect 12713 14903 12771 14909
rect 13446 14900 13452 14912
rect 13504 14900 13510 14952
rect 14366 14940 14372 14952
rect 14327 14912 14372 14940
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 22624 14943 22682 14949
rect 22624 14909 22636 14943
rect 22670 14940 22682 14943
rect 23106 14940 23112 14952
rect 22670 14912 23112 14940
rect 22670 14909 22682 14912
rect 22624 14903 22682 14909
rect 23106 14900 23112 14912
rect 23164 14900 23170 14952
rect 25292 14943 25350 14949
rect 25292 14909 25304 14943
rect 25338 14940 25350 14943
rect 25774 14940 25780 14952
rect 25338 14912 25780 14940
rect 25338 14909 25350 14912
rect 25292 14903 25350 14909
rect 25774 14900 25780 14912
rect 25832 14900 25838 14952
rect 14690 14875 14748 14881
rect 14690 14872 14702 14875
rect 14292 14844 14702 14872
rect 14292 14816 14320 14844
rect 14690 14841 14702 14844
rect 14736 14841 14748 14875
rect 16482 14872 16488 14884
rect 16443 14844 16488 14872
rect 14690 14835 14748 14841
rect 16482 14832 16488 14844
rect 16540 14832 16546 14884
rect 16577 14875 16635 14881
rect 16577 14841 16589 14875
rect 16623 14841 16635 14875
rect 18138 14872 18144 14884
rect 18099 14844 18144 14872
rect 16577 14835 16635 14841
rect 14274 14804 14280 14816
rect 14235 14776 14280 14804
rect 14274 14764 14280 14776
rect 14332 14764 14338 14816
rect 16390 14764 16396 14816
rect 16448 14804 16454 14816
rect 16592 14804 16620 14835
rect 18138 14832 18144 14844
rect 18196 14832 18202 14884
rect 18233 14875 18291 14881
rect 18233 14841 18245 14875
rect 18279 14841 18291 14875
rect 20809 14875 20867 14881
rect 20809 14872 20821 14875
rect 18233 14835 18291 14841
rect 20180 14844 20821 14872
rect 16448 14776 16620 14804
rect 16448 14764 16454 14776
rect 17034 14764 17040 14816
rect 17092 14804 17098 14816
rect 17773 14807 17831 14813
rect 17773 14804 17785 14807
rect 17092 14776 17785 14804
rect 17092 14764 17098 14776
rect 17773 14773 17785 14776
rect 17819 14804 17831 14807
rect 18248 14804 18276 14835
rect 20180 14816 20208 14844
rect 20809 14841 20821 14844
rect 20855 14841 20867 14875
rect 20809 14835 20867 14841
rect 20901 14875 20959 14881
rect 20901 14841 20913 14875
rect 20947 14841 20959 14875
rect 20901 14835 20959 14841
rect 21453 14875 21511 14881
rect 21453 14841 21465 14875
rect 21499 14872 21511 14875
rect 21818 14872 21824 14884
rect 21499 14844 21824 14872
rect 21499 14841 21511 14844
rect 21453 14835 21511 14841
rect 19426 14804 19432 14816
rect 17819 14776 18276 14804
rect 19387 14776 19432 14804
rect 17819 14773 17831 14776
rect 17773 14767 17831 14773
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 20162 14804 20168 14816
rect 20123 14776 20168 14804
rect 20162 14764 20168 14776
rect 20220 14764 20226 14816
rect 20714 14764 20720 14816
rect 20772 14804 20778 14816
rect 20916 14804 20944 14835
rect 21818 14832 21824 14844
rect 21876 14872 21882 14884
rect 22189 14875 22247 14881
rect 22189 14872 22201 14875
rect 21876 14844 22201 14872
rect 21876 14832 21882 14844
rect 22189 14841 22201 14844
rect 22235 14872 22247 14875
rect 23382 14872 23388 14884
rect 22235 14844 23388 14872
rect 22235 14841 22247 14844
rect 22189 14835 22247 14841
rect 23382 14832 23388 14844
rect 23440 14832 23446 14884
rect 23842 14832 23848 14884
rect 23900 14872 23906 14884
rect 24397 14875 24455 14881
rect 23900 14844 23945 14872
rect 23900 14832 23906 14844
rect 24397 14841 24409 14875
rect 24443 14872 24455 14875
rect 24578 14872 24584 14884
rect 24443 14844 24584 14872
rect 24443 14841 24455 14844
rect 24397 14835 24455 14841
rect 24578 14832 24584 14844
rect 24636 14872 24642 14884
rect 24854 14872 24860 14884
rect 24636 14844 24860 14872
rect 24636 14832 24642 14844
rect 24854 14832 24860 14844
rect 24912 14832 24918 14884
rect 20772 14776 20944 14804
rect 20772 14764 20778 14776
rect 20990 14764 20996 14816
rect 21048 14804 21054 14816
rect 22695 14807 22753 14813
rect 22695 14804 22707 14807
rect 21048 14776 22707 14804
rect 21048 14764 21054 14776
rect 22695 14773 22707 14776
rect 22741 14773 22753 14807
rect 22695 14767 22753 14773
rect 23477 14807 23535 14813
rect 23477 14773 23489 14807
rect 23523 14804 23535 14807
rect 23860 14804 23888 14832
rect 23523 14776 23888 14804
rect 23523 14773 23535 14776
rect 23477 14767 23535 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 12759 14603 12817 14609
rect 12759 14569 12771 14603
rect 12805 14600 12817 14603
rect 13541 14603 13599 14609
rect 13541 14600 13553 14603
rect 12805 14572 13553 14600
rect 12805 14569 12817 14572
rect 12759 14563 12817 14569
rect 13541 14569 13553 14572
rect 13587 14600 13599 14603
rect 13722 14600 13728 14612
rect 13587 14572 13728 14600
rect 13587 14569 13599 14572
rect 13541 14563 13599 14569
rect 13722 14560 13728 14572
rect 13780 14560 13786 14612
rect 15565 14603 15623 14609
rect 15565 14569 15577 14603
rect 15611 14600 15623 14603
rect 15654 14600 15660 14612
rect 15611 14572 15660 14600
rect 15611 14569 15623 14572
rect 15565 14563 15623 14569
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 17034 14600 17040 14612
rect 16995 14572 17040 14600
rect 17034 14560 17040 14572
rect 17092 14560 17098 14612
rect 17402 14600 17408 14612
rect 17363 14572 17408 14600
rect 17402 14560 17408 14572
rect 17460 14560 17466 14612
rect 18785 14603 18843 14609
rect 18785 14569 18797 14603
rect 18831 14600 18843 14603
rect 18966 14600 18972 14612
rect 18831 14572 18972 14600
rect 18831 14569 18843 14572
rect 18785 14563 18843 14569
rect 18966 14560 18972 14572
rect 19024 14560 19030 14612
rect 21269 14603 21327 14609
rect 21269 14600 21281 14603
rect 19996 14572 21281 14600
rect 14274 14492 14280 14544
rect 14332 14532 14338 14544
rect 16438 14535 16496 14541
rect 16438 14532 16450 14535
rect 14332 14504 16450 14532
rect 14332 14492 14338 14504
rect 16438 14501 16450 14504
rect 16484 14532 16496 14535
rect 16850 14532 16856 14544
rect 16484 14504 16856 14532
rect 16484 14501 16496 14504
rect 16438 14495 16496 14501
rect 16850 14492 16856 14504
rect 16908 14532 16914 14544
rect 18186 14535 18244 14541
rect 18186 14532 18198 14535
rect 16908 14504 18198 14532
rect 16908 14492 16914 14504
rect 18186 14501 18198 14504
rect 18232 14532 18244 14535
rect 19996 14532 20024 14572
rect 21269 14569 21281 14572
rect 21315 14569 21327 14603
rect 21269 14563 21327 14569
rect 21821 14603 21879 14609
rect 21821 14569 21833 14603
rect 21867 14600 21879 14603
rect 21910 14600 21916 14612
rect 21867 14572 21916 14600
rect 21867 14569 21879 14572
rect 21821 14563 21879 14569
rect 21910 14560 21916 14572
rect 21968 14560 21974 14612
rect 23750 14600 23756 14612
rect 23711 14572 23756 14600
rect 23750 14560 23756 14572
rect 23808 14560 23814 14612
rect 22830 14532 22836 14544
rect 18232 14504 20024 14532
rect 22204 14504 22836 14532
rect 18232 14501 18244 14504
rect 18186 14495 18244 14501
rect 6362 14464 6368 14476
rect 6323 14436 6368 14464
rect 6362 14424 6368 14436
rect 6420 14424 6426 14476
rect 12688 14467 12746 14473
rect 12688 14433 12700 14467
rect 12734 14464 12746 14467
rect 13078 14464 13084 14476
rect 12734 14436 13084 14464
rect 12734 14433 12746 14436
rect 12688 14427 12746 14433
rect 13078 14424 13084 14436
rect 13136 14424 13142 14476
rect 13354 14424 13360 14476
rect 13412 14464 13418 14476
rect 13633 14467 13691 14473
rect 13633 14464 13645 14467
rect 13412 14436 13645 14464
rect 13412 14424 13418 14436
rect 13633 14433 13645 14436
rect 13679 14433 13691 14467
rect 14090 14464 14096 14476
rect 14051 14436 14096 14464
rect 13633 14427 13691 14433
rect 14090 14424 14096 14436
rect 14148 14424 14154 14476
rect 20806 14424 20812 14476
rect 20864 14464 20870 14476
rect 22204 14464 22232 14504
rect 22830 14492 22836 14504
rect 22888 14492 22894 14544
rect 23382 14532 23388 14544
rect 23343 14504 23388 14532
rect 23382 14492 23388 14504
rect 23440 14492 23446 14544
rect 24397 14535 24455 14541
rect 24397 14501 24409 14535
rect 24443 14532 24455 14535
rect 25130 14532 25136 14544
rect 24443 14504 25136 14532
rect 24443 14501 24455 14504
rect 24397 14495 24455 14501
rect 25130 14492 25136 14504
rect 25188 14492 25194 14544
rect 20864 14436 22232 14464
rect 20864 14424 20870 14436
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14396 14427 14399
rect 15930 14396 15936 14408
rect 14415 14368 15936 14396
rect 14415 14365 14427 14368
rect 14369 14359 14427 14365
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 16114 14396 16120 14408
rect 16075 14368 16120 14396
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 17862 14396 17868 14408
rect 17823 14368 17868 14396
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 19797 14399 19855 14405
rect 19797 14365 19809 14399
rect 19843 14396 19855 14399
rect 20714 14396 20720 14408
rect 19843 14368 20720 14396
rect 19843 14365 19855 14368
rect 19797 14359 19855 14365
rect 20714 14356 20720 14368
rect 20772 14356 20778 14408
rect 20898 14396 20904 14408
rect 20859 14368 20904 14396
rect 20898 14356 20904 14368
rect 20956 14356 20962 14408
rect 22741 14399 22799 14405
rect 22741 14365 22753 14399
rect 22787 14396 22799 14399
rect 23566 14396 23572 14408
rect 22787 14368 23572 14396
rect 22787 14365 22799 14368
rect 22741 14359 22799 14365
rect 23566 14356 23572 14368
rect 23624 14356 23630 14408
rect 24026 14356 24032 14408
rect 24084 14396 24090 14408
rect 24305 14399 24363 14405
rect 24305 14396 24317 14399
rect 24084 14368 24317 14396
rect 24084 14356 24090 14368
rect 24305 14365 24317 14368
rect 24351 14365 24363 14399
rect 24578 14396 24584 14408
rect 24539 14368 24584 14396
rect 24305 14359 24363 14365
rect 24578 14356 24584 14368
rect 24636 14356 24642 14408
rect 6595 14331 6653 14337
rect 6595 14297 6607 14331
rect 6641 14328 6653 14331
rect 12618 14328 12624 14340
rect 6641 14300 12624 14328
rect 6641 14297 6653 14300
rect 6595 14291 6653 14297
rect 12618 14288 12624 14300
rect 12676 14288 12682 14340
rect 14366 14220 14372 14272
rect 14424 14260 14430 14272
rect 14645 14263 14703 14269
rect 14645 14260 14657 14263
rect 14424 14232 14657 14260
rect 14424 14220 14430 14232
rect 14645 14229 14657 14232
rect 14691 14229 14703 14263
rect 14645 14223 14703 14229
rect 18874 14220 18880 14272
rect 18932 14260 18938 14272
rect 19061 14263 19119 14269
rect 19061 14260 19073 14263
rect 18932 14232 19073 14260
rect 18932 14220 18938 14232
rect 19061 14229 19073 14232
rect 19107 14229 19119 14263
rect 19061 14223 19119 14229
rect 21910 14220 21916 14272
rect 21968 14260 21974 14272
rect 22097 14263 22155 14269
rect 22097 14260 22109 14263
rect 21968 14232 22109 14260
rect 21968 14220 21974 14232
rect 22097 14229 22109 14232
rect 22143 14229 22155 14263
rect 22097 14223 22155 14229
rect 23750 14220 23756 14272
rect 23808 14260 23814 14272
rect 24029 14263 24087 14269
rect 24029 14260 24041 14263
rect 23808 14232 24041 14260
rect 23808 14220 23814 14232
rect 24029 14229 24041 14232
rect 24075 14229 24087 14263
rect 24029 14223 24087 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 14090 14056 14096 14068
rect 13188 14028 14096 14056
rect 12713 13991 12771 13997
rect 12713 13957 12725 13991
rect 12759 13988 12771 13991
rect 13078 13988 13084 14000
rect 12759 13960 13084 13988
rect 12759 13957 12771 13960
rect 12713 13951 12771 13957
rect 13078 13948 13084 13960
rect 13136 13948 13142 14000
rect 13188 13920 13216 14028
rect 14090 14016 14096 14028
rect 14148 14016 14154 14068
rect 15930 14016 15936 14068
rect 15988 14056 15994 14068
rect 17405 14059 17463 14065
rect 17405 14056 17417 14059
rect 15988 14028 17417 14056
rect 15988 14016 15994 14028
rect 17405 14025 17417 14028
rect 17451 14056 17463 14059
rect 17862 14056 17868 14068
rect 17451 14028 17868 14056
rect 17451 14025 17463 14028
rect 17405 14019 17463 14025
rect 17862 14016 17868 14028
rect 17920 14016 17926 14068
rect 19794 14016 19800 14068
rect 19852 14056 19858 14068
rect 19889 14059 19947 14065
rect 19889 14056 19901 14059
rect 19852 14028 19901 14056
rect 19852 14016 19858 14028
rect 19889 14025 19901 14028
rect 19935 14025 19947 14059
rect 19889 14019 19947 14025
rect 20806 14016 20812 14068
rect 20864 14056 20870 14068
rect 20901 14059 20959 14065
rect 20901 14056 20913 14059
rect 20864 14028 20913 14056
rect 20864 14016 20870 14028
rect 20901 14025 20913 14028
rect 20947 14025 20959 14059
rect 20901 14019 20959 14025
rect 22649 14059 22707 14065
rect 22649 14025 22661 14059
rect 22695 14056 22707 14059
rect 24765 14059 24823 14065
rect 24765 14056 24777 14059
rect 22695 14028 24777 14056
rect 22695 14025 22707 14028
rect 22649 14019 22707 14025
rect 24765 14025 24777 14028
rect 24811 14056 24823 14059
rect 25130 14056 25136 14068
rect 24811 14028 25136 14056
rect 24811 14025 24823 14028
rect 24765 14019 24823 14025
rect 25130 14016 25136 14028
rect 25188 14016 25194 14068
rect 25774 14056 25780 14068
rect 25735 14028 25780 14056
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 13446 13948 13452 14000
rect 13504 13988 13510 14000
rect 14921 13991 14979 13997
rect 14921 13988 14933 13991
rect 13504 13960 14933 13988
rect 13504 13948 13510 13960
rect 14921 13957 14933 13960
rect 14967 13988 14979 13991
rect 16206 13988 16212 14000
rect 14967 13960 16212 13988
rect 14967 13957 14979 13960
rect 14921 13951 14979 13957
rect 16206 13948 16212 13960
rect 16264 13948 16270 14000
rect 16850 13988 16856 14000
rect 16811 13960 16856 13988
rect 16850 13948 16856 13960
rect 16908 13988 16914 14000
rect 17773 13991 17831 13997
rect 17773 13988 17785 13991
rect 16908 13960 17785 13988
rect 16908 13948 16914 13960
rect 17773 13957 17785 13960
rect 17819 13957 17831 13991
rect 17773 13951 17831 13957
rect 18782 13948 18788 14000
rect 18840 13988 18846 14000
rect 18969 13991 19027 13997
rect 18969 13988 18981 13991
rect 18840 13960 18981 13988
rect 18840 13948 18846 13960
rect 18969 13957 18981 13960
rect 19015 13988 19027 13991
rect 19426 13988 19432 14000
rect 19015 13960 19432 13988
rect 19015 13957 19027 13960
rect 18969 13951 19027 13957
rect 19426 13948 19432 13960
rect 19484 13948 19490 14000
rect 20530 13948 20536 14000
rect 20588 13988 20594 14000
rect 21910 13988 21916 14000
rect 20588 13960 21916 13988
rect 20588 13948 20594 13960
rect 21910 13948 21916 13960
rect 21968 13948 21974 14000
rect 22830 13948 22836 14000
rect 22888 13988 22894 14000
rect 22925 13991 22983 13997
rect 22925 13988 22937 13991
rect 22888 13960 22937 13988
rect 22888 13948 22894 13960
rect 22925 13957 22937 13960
rect 22971 13957 22983 13991
rect 22925 13951 22983 13957
rect 15657 13923 15715 13929
rect 15657 13920 15669 13923
rect 13096 13892 13216 13920
rect 14108 13892 15669 13920
rect 12342 13812 12348 13864
rect 12400 13852 12406 13864
rect 13096 13861 13124 13892
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 12400 13824 13093 13852
rect 12400 13812 12406 13824
rect 13081 13821 13093 13824
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 13722 13812 13728 13864
rect 13780 13852 13786 13864
rect 14001 13855 14059 13861
rect 14001 13852 14013 13855
rect 13780 13824 14013 13852
rect 13780 13812 13786 13824
rect 14001 13821 14013 13824
rect 14047 13821 14059 13855
rect 14001 13815 14059 13821
rect 13262 13744 13268 13796
rect 13320 13784 13326 13796
rect 14108 13784 14136 13892
rect 15657 13889 15669 13892
rect 15703 13920 15715 13923
rect 18417 13923 18475 13929
rect 15703 13892 15884 13920
rect 15703 13889 15715 13892
rect 15657 13883 15715 13889
rect 14274 13852 14280 13864
rect 14187 13824 14280 13852
rect 13320 13756 14136 13784
rect 13320 13744 13326 13756
rect 6362 13676 6368 13728
rect 6420 13716 6426 13728
rect 6457 13719 6515 13725
rect 6457 13716 6469 13719
rect 6420 13688 6469 13716
rect 6420 13676 6426 13688
rect 6457 13685 6469 13688
rect 6503 13685 6515 13719
rect 6457 13679 6515 13685
rect 13354 13676 13360 13728
rect 13412 13716 13418 13728
rect 13449 13719 13507 13725
rect 13449 13716 13461 13719
rect 13412 13688 13461 13716
rect 13412 13676 13418 13688
rect 13449 13685 13461 13688
rect 13495 13685 13507 13719
rect 13814 13716 13820 13728
rect 13775 13688 13820 13716
rect 13449 13679 13507 13685
rect 13814 13676 13820 13688
rect 13872 13716 13878 13728
rect 14200 13716 14228 13824
rect 14274 13812 14280 13824
rect 14332 13852 14338 13864
rect 15856 13861 15884 13892
rect 18417 13889 18429 13923
rect 18463 13920 18475 13923
rect 18874 13920 18880 13932
rect 18463 13892 18880 13920
rect 18463 13889 18475 13892
rect 18417 13883 18475 13889
rect 18874 13880 18880 13892
rect 18932 13920 18938 13932
rect 19150 13920 19156 13932
rect 18932 13892 19156 13920
rect 18932 13880 18938 13892
rect 19150 13880 19156 13892
rect 19208 13880 19214 13932
rect 19521 13923 19579 13929
rect 19521 13889 19533 13923
rect 19567 13920 19579 13923
rect 19981 13923 20039 13929
rect 19981 13920 19993 13923
rect 19567 13892 19993 13920
rect 19567 13889 19579 13892
rect 19521 13883 19579 13889
rect 19981 13889 19993 13892
rect 20027 13920 20039 13923
rect 21818 13920 21824 13932
rect 20027 13892 21824 13920
rect 20027 13889 20039 13892
rect 19981 13883 20039 13889
rect 21818 13880 21824 13892
rect 21876 13880 21882 13932
rect 22002 13880 22008 13932
rect 22060 13920 22066 13932
rect 22060 13892 23152 13920
rect 22060 13880 22066 13892
rect 15841 13855 15899 13861
rect 14332 13824 14412 13852
rect 14332 13812 14338 13824
rect 14384 13793 14412 13824
rect 15841 13821 15853 13855
rect 15887 13821 15899 13855
rect 15841 13815 15899 13821
rect 15930 13812 15936 13864
rect 15988 13852 15994 13864
rect 16301 13855 16359 13861
rect 16301 13852 16313 13855
rect 15988 13824 16313 13852
rect 15988 13812 15994 13824
rect 16301 13821 16313 13824
rect 16347 13821 16359 13855
rect 16301 13815 16359 13821
rect 21729 13855 21787 13861
rect 21729 13821 21741 13855
rect 21775 13852 21787 13855
rect 21910 13852 21916 13864
rect 21775 13824 21916 13852
rect 21775 13821 21787 13824
rect 21729 13815 21787 13821
rect 21910 13812 21916 13824
rect 21968 13812 21974 13864
rect 23124 13814 23152 13892
rect 23198 13880 23204 13932
rect 23256 13920 23262 13932
rect 24026 13920 24032 13932
rect 23256 13892 24032 13920
rect 23256 13880 23262 13892
rect 24026 13880 24032 13892
rect 24084 13920 24090 13932
rect 25041 13923 25099 13929
rect 25041 13920 25053 13923
rect 24084 13892 25053 13920
rect 24084 13880 24090 13892
rect 25041 13889 25053 13892
rect 25087 13889 25099 13923
rect 25041 13883 25099 13889
rect 23385 13855 23443 13861
rect 23385 13852 23397 13855
rect 23216 13824 23397 13852
rect 23216 13814 23244 13824
rect 23385 13821 23397 13824
rect 23431 13821 23443 13855
rect 23385 13815 23443 13821
rect 25292 13855 25350 13861
rect 25292 13821 25304 13855
rect 25338 13852 25350 13855
rect 25774 13852 25780 13864
rect 25338 13824 25780 13852
rect 25338 13821 25350 13824
rect 25292 13815 25350 13821
rect 14363 13787 14421 13793
rect 14363 13753 14375 13787
rect 14409 13753 14421 13787
rect 14363 13747 14421 13753
rect 18509 13787 18567 13793
rect 18509 13753 18521 13787
rect 18555 13753 18567 13787
rect 18509 13747 18567 13753
rect 16114 13716 16120 13728
rect 13872 13688 14228 13716
rect 16075 13688 16120 13716
rect 13872 13676 13878 13688
rect 16114 13676 16120 13688
rect 16172 13676 16178 13728
rect 18322 13676 18328 13728
rect 18380 13716 18386 13728
rect 18524 13716 18552 13747
rect 19794 13744 19800 13796
rect 19852 13784 19858 13796
rect 20343 13787 20401 13793
rect 20343 13784 20355 13787
rect 19852 13756 20355 13784
rect 19852 13744 19858 13756
rect 20343 13753 20355 13756
rect 20389 13784 20401 13787
rect 22050 13787 22108 13793
rect 20389 13756 21312 13784
rect 20389 13753 20401 13756
rect 20343 13747 20401 13753
rect 21284 13728 21312 13756
rect 22050 13753 22062 13787
rect 22096 13753 22108 13787
rect 23124 13786 23244 13814
rect 22050 13747 22108 13753
rect 21266 13716 21272 13728
rect 18380 13688 18552 13716
rect 21227 13688 21272 13716
rect 18380 13676 18386 13688
rect 21266 13676 21272 13688
rect 21324 13716 21330 13728
rect 21545 13719 21603 13725
rect 21545 13716 21557 13719
rect 21324 13688 21557 13716
rect 21324 13676 21330 13688
rect 21545 13685 21557 13688
rect 21591 13716 21603 13719
rect 22065 13716 22093 13747
rect 21591 13688 22093 13716
rect 23400 13716 23428 13815
rect 25774 13812 25780 13824
rect 25832 13812 25838 13864
rect 23750 13784 23756 13796
rect 23711 13756 23756 13784
rect 23750 13744 23756 13756
rect 23808 13744 23814 13796
rect 23845 13787 23903 13793
rect 23845 13753 23857 13787
rect 23891 13753 23903 13787
rect 23845 13747 23903 13753
rect 23860 13716 23888 13747
rect 23400 13688 23888 13716
rect 21591 13685 21603 13688
rect 21545 13679 21603 13685
rect 24302 13676 24308 13728
rect 24360 13716 24366 13728
rect 25363 13719 25421 13725
rect 25363 13716 25375 13719
rect 24360 13688 25375 13716
rect 24360 13676 24366 13688
rect 25363 13685 25375 13688
rect 25409 13685 25421 13719
rect 25363 13679 25421 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 16114 13472 16120 13524
rect 16172 13512 16178 13524
rect 16209 13515 16267 13521
rect 16209 13512 16221 13515
rect 16172 13484 16221 13512
rect 16172 13472 16178 13484
rect 16209 13481 16221 13484
rect 16255 13481 16267 13515
rect 16209 13475 16267 13481
rect 17681 13515 17739 13521
rect 17681 13481 17693 13515
rect 17727 13512 17739 13515
rect 17770 13512 17776 13524
rect 17727 13484 17776 13512
rect 17727 13481 17739 13484
rect 17681 13475 17739 13481
rect 17770 13472 17776 13484
rect 17828 13472 17834 13524
rect 14366 13444 14372 13456
rect 14327 13416 14372 13444
rect 14366 13404 14372 13416
rect 14424 13404 14430 13456
rect 16850 13404 16856 13456
rect 16908 13444 16914 13456
rect 17082 13447 17140 13453
rect 17082 13444 17094 13447
rect 16908 13416 17094 13444
rect 16908 13404 16914 13416
rect 17082 13413 17094 13416
rect 17128 13413 17140 13447
rect 18693 13447 18751 13453
rect 18693 13444 18705 13447
rect 17082 13407 17140 13413
rect 17236 13416 18705 13444
rect 12618 13376 12624 13388
rect 12579 13348 12624 13376
rect 12618 13336 12624 13348
rect 12676 13336 12682 13388
rect 13906 13376 13912 13388
rect 13867 13348 13912 13376
rect 13906 13336 13912 13348
rect 13964 13336 13970 13388
rect 14185 13379 14243 13385
rect 14185 13345 14197 13379
rect 14231 13376 14243 13379
rect 14458 13376 14464 13388
rect 14231 13348 14464 13376
rect 14231 13345 14243 13348
rect 14185 13339 14243 13345
rect 14458 13336 14464 13348
rect 14516 13336 14522 13388
rect 17236 13376 17264 13416
rect 18693 13413 18705 13416
rect 18739 13444 18751 13447
rect 19242 13444 19248 13456
rect 18739 13416 19248 13444
rect 18739 13413 18751 13416
rect 18693 13407 18751 13413
rect 19242 13404 19248 13416
rect 19300 13404 19306 13456
rect 22649 13447 22707 13453
rect 22649 13413 22661 13447
rect 22695 13444 22707 13447
rect 22738 13444 22744 13456
rect 22695 13416 22744 13444
rect 22695 13413 22707 13416
rect 22649 13407 22707 13413
rect 22738 13404 22744 13416
rect 22796 13404 22802 13456
rect 23198 13444 23204 13456
rect 23159 13416 23204 13444
rect 23198 13404 23204 13416
rect 23256 13404 23262 13456
rect 24210 13444 24216 13456
rect 24123 13416 24216 13444
rect 24210 13404 24216 13416
rect 24268 13444 24274 13456
rect 24854 13444 24860 13456
rect 24268 13416 24860 13444
rect 24268 13404 24274 13416
rect 24854 13404 24860 13416
rect 24912 13404 24918 13456
rect 15212 13348 17264 13376
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13308 12863 13311
rect 15212 13308 15240 13348
rect 20806 13336 20812 13388
rect 20864 13376 20870 13388
rect 20901 13379 20959 13385
rect 20901 13376 20913 13379
rect 20864 13348 20913 13376
rect 20864 13336 20870 13348
rect 20901 13345 20913 13348
rect 20947 13345 20959 13379
rect 20901 13339 20959 13345
rect 21361 13379 21419 13385
rect 21361 13345 21373 13379
rect 21407 13345 21419 13379
rect 21361 13339 21419 13345
rect 12851 13280 15240 13308
rect 15289 13311 15347 13317
rect 12851 13277 12863 13280
rect 12805 13271 12863 13277
rect 15289 13277 15301 13311
rect 15335 13308 15347 13311
rect 15378 13308 15384 13320
rect 15335 13280 15384 13308
rect 15335 13277 15347 13280
rect 15289 13271 15347 13277
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 16758 13308 16764 13320
rect 16719 13280 16764 13308
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 18601 13311 18659 13317
rect 18601 13308 18613 13311
rect 17972 13280 18613 13308
rect 14550 13200 14556 13252
rect 14608 13240 14614 13252
rect 17972 13249 18000 13280
rect 18601 13277 18613 13280
rect 18647 13277 18659 13311
rect 18601 13271 18659 13277
rect 18782 13268 18788 13320
rect 18840 13308 18846 13320
rect 18877 13311 18935 13317
rect 18877 13308 18889 13311
rect 18840 13280 18889 13308
rect 18840 13268 18846 13280
rect 18877 13277 18889 13280
rect 18923 13277 18935 13311
rect 21376 13308 21404 13339
rect 21634 13308 21640 13320
rect 18877 13271 18935 13277
rect 20272 13280 21404 13308
rect 21547 13280 21640 13308
rect 17957 13243 18015 13249
rect 17957 13240 17969 13243
rect 14608 13212 17969 13240
rect 14608 13200 14614 13212
rect 17957 13209 17969 13212
rect 18003 13209 18015 13243
rect 17957 13203 18015 13209
rect 20272 13184 20300 13280
rect 21634 13268 21640 13280
rect 21692 13308 21698 13320
rect 21913 13311 21971 13317
rect 21913 13308 21925 13311
rect 21692 13280 21925 13308
rect 21692 13268 21698 13280
rect 21913 13277 21925 13280
rect 21959 13277 21971 13311
rect 21913 13271 21971 13277
rect 22557 13311 22615 13317
rect 22557 13277 22569 13311
rect 22603 13308 22615 13311
rect 22830 13308 22836 13320
rect 22603 13280 22836 13308
rect 22603 13277 22615 13280
rect 22557 13271 22615 13277
rect 22830 13268 22836 13280
rect 22888 13268 22894 13320
rect 24118 13308 24124 13320
rect 23446 13280 24124 13308
rect 20714 13200 20720 13252
rect 20772 13240 20778 13252
rect 23446 13240 23474 13280
rect 24118 13268 24124 13280
rect 24176 13268 24182 13320
rect 24670 13240 24676 13252
rect 20772 13212 23474 13240
rect 24631 13212 24676 13240
rect 20772 13200 20778 13212
rect 24670 13200 24676 13212
rect 24728 13200 24734 13252
rect 13722 13132 13728 13184
rect 13780 13172 13786 13184
rect 14645 13175 14703 13181
rect 14645 13172 14657 13175
rect 13780 13144 14657 13172
rect 13780 13132 13786 13144
rect 14645 13141 14657 13144
rect 14691 13141 14703 13175
rect 15838 13172 15844 13184
rect 15799 13144 15844 13172
rect 14645 13135 14703 13141
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 18322 13172 18328 13184
rect 18283 13144 18328 13172
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 18414 13132 18420 13184
rect 18472 13172 18478 13184
rect 19797 13175 19855 13181
rect 19797 13172 19809 13175
rect 18472 13144 19809 13172
rect 18472 13132 18478 13144
rect 19797 13141 19809 13144
rect 19843 13172 19855 13175
rect 20254 13172 20260 13184
rect 19843 13144 20260 13172
rect 19843 13141 19855 13144
rect 19797 13135 19855 13141
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 20625 13175 20683 13181
rect 20625 13141 20637 13175
rect 20671 13172 20683 13175
rect 20898 13172 20904 13184
rect 20671 13144 20904 13172
rect 20671 13141 20683 13144
rect 20625 13135 20683 13141
rect 20898 13132 20904 13144
rect 20956 13172 20962 13184
rect 23014 13172 23020 13184
rect 20956 13144 23020 13172
rect 20956 13132 20962 13144
rect 23014 13132 23020 13144
rect 23072 13132 23078 13184
rect 23566 13172 23572 13184
rect 23527 13144 23572 13172
rect 23566 13132 23572 13144
rect 23624 13132 23630 13184
rect 23934 13172 23940 13184
rect 23895 13144 23940 13172
rect 23934 13132 23940 13144
rect 23992 13132 23998 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 12161 12971 12219 12977
rect 12161 12937 12173 12971
rect 12207 12968 12219 12971
rect 12618 12968 12624 12980
rect 12207 12940 12624 12968
rect 12207 12937 12219 12940
rect 12161 12931 12219 12937
rect 12618 12928 12624 12940
rect 12676 12968 12682 12980
rect 18322 12968 18328 12980
rect 12676 12940 18328 12968
rect 12676 12928 12682 12940
rect 18322 12928 18328 12940
rect 18380 12968 18386 12980
rect 18969 12971 19027 12977
rect 18969 12968 18981 12971
rect 18380 12940 18981 12968
rect 18380 12928 18386 12940
rect 18969 12937 18981 12940
rect 19015 12937 19027 12971
rect 19242 12968 19248 12980
rect 19203 12940 19248 12968
rect 18969 12931 19027 12937
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 22002 12928 22008 12980
rect 22060 12968 22066 12980
rect 22281 12971 22339 12977
rect 22281 12968 22293 12971
rect 22060 12940 22293 12968
rect 22060 12928 22066 12940
rect 22281 12937 22293 12940
rect 22327 12937 22339 12971
rect 22281 12931 22339 12937
rect 22649 12971 22707 12977
rect 22649 12937 22661 12971
rect 22695 12968 22707 12971
rect 22738 12968 22744 12980
rect 22695 12940 22744 12968
rect 22695 12937 22707 12940
rect 22649 12931 22707 12937
rect 22738 12928 22744 12940
rect 22796 12928 22802 12980
rect 24854 12968 24860 12980
rect 24815 12940 24860 12968
rect 24854 12928 24860 12940
rect 24912 12928 24918 12980
rect 12526 12860 12532 12912
rect 12584 12900 12590 12912
rect 12584 12872 18092 12900
rect 12584 12860 12590 12872
rect 13722 12832 13728 12844
rect 13683 12804 13728 12832
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 14645 12835 14703 12841
rect 14645 12801 14657 12835
rect 14691 12832 14703 12835
rect 14826 12832 14832 12844
rect 14691 12804 14832 12832
rect 14691 12801 14703 12804
rect 14645 12795 14703 12801
rect 14826 12792 14832 12804
rect 14884 12792 14890 12844
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12832 15347 12835
rect 15562 12832 15568 12844
rect 15335 12804 15568 12832
rect 15335 12801 15347 12804
rect 15289 12795 15347 12801
rect 15562 12792 15568 12804
rect 15620 12792 15626 12844
rect 16758 12832 16764 12844
rect 16719 12804 16764 12832
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 18064 12841 18092 12872
rect 23750 12860 23756 12912
rect 23808 12900 23814 12912
rect 25547 12903 25605 12909
rect 25547 12900 25559 12903
rect 23808 12872 25559 12900
rect 23808 12860 23814 12872
rect 25547 12869 25559 12872
rect 25593 12869 25605 12903
rect 25547 12863 25605 12869
rect 18049 12835 18107 12841
rect 18049 12801 18061 12835
rect 18095 12832 18107 12835
rect 18690 12832 18696 12844
rect 18095 12804 18696 12832
rect 18095 12801 18107 12804
rect 18049 12795 18107 12801
rect 18690 12792 18696 12804
rect 18748 12792 18754 12844
rect 20530 12832 20536 12844
rect 19536 12804 20392 12832
rect 20491 12804 20536 12832
rect 12710 12724 12716 12776
rect 12768 12764 12774 12776
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12768 12736 12909 12764
rect 12768 12724 12774 12736
rect 12897 12733 12909 12736
rect 12943 12764 12955 12767
rect 13262 12764 13268 12776
rect 12943 12736 13268 12764
rect 12943 12733 12955 12736
rect 12897 12727 12955 12733
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 13538 12764 13544 12776
rect 13451 12736 13544 12764
rect 13538 12724 13544 12736
rect 13596 12764 13602 12776
rect 14458 12764 14464 12776
rect 13596 12736 14464 12764
rect 13596 12724 13602 12736
rect 14458 12724 14464 12736
rect 14516 12724 14522 12776
rect 16022 12724 16028 12776
rect 16080 12764 16086 12776
rect 16117 12767 16175 12773
rect 16117 12764 16129 12767
rect 16080 12736 16129 12764
rect 16080 12724 16086 12736
rect 16117 12733 16129 12736
rect 16163 12733 16175 12767
rect 16666 12764 16672 12776
rect 16627 12736 16672 12764
rect 16117 12727 16175 12733
rect 16666 12724 16672 12736
rect 16724 12724 16730 12776
rect 17221 12767 17279 12773
rect 17221 12733 17233 12767
rect 17267 12764 17279 12767
rect 17865 12767 17923 12773
rect 17865 12764 17877 12767
rect 17267 12736 17877 12764
rect 17267 12733 17279 12736
rect 17221 12727 17279 12733
rect 17865 12733 17877 12736
rect 17911 12764 17923 12767
rect 19536 12764 19564 12804
rect 19797 12767 19855 12773
rect 19797 12764 19809 12767
rect 17911 12736 19564 12764
rect 19628 12736 19809 12764
rect 17911 12733 17923 12736
rect 17865 12727 17923 12733
rect 14734 12656 14740 12708
rect 14792 12696 14798 12708
rect 15657 12699 15715 12705
rect 14792 12668 14837 12696
rect 14792 12656 14798 12668
rect 15657 12665 15669 12699
rect 15703 12696 15715 12699
rect 15838 12696 15844 12708
rect 15703 12668 15844 12696
rect 15703 12665 15715 12668
rect 15657 12659 15715 12665
rect 15838 12656 15844 12668
rect 15896 12696 15902 12708
rect 16684 12696 16712 12724
rect 18426 12705 18454 12736
rect 18411 12699 18469 12705
rect 18411 12696 18423 12699
rect 15896 12668 16712 12696
rect 18389 12668 18423 12696
rect 15896 12656 15902 12668
rect 18411 12665 18423 12668
rect 18457 12665 18469 12699
rect 18411 12659 18469 12665
rect 13262 12588 13268 12640
rect 13320 12628 13326 12640
rect 13906 12628 13912 12640
rect 13320 12600 13912 12628
rect 13320 12588 13326 12600
rect 13906 12588 13912 12600
rect 13964 12628 13970 12640
rect 14001 12631 14059 12637
rect 14001 12628 14013 12631
rect 13964 12600 14013 12628
rect 13964 12588 13970 12600
rect 14001 12597 14013 12600
rect 14047 12597 14059 12631
rect 14458 12628 14464 12640
rect 14419 12600 14464 12628
rect 14001 12591 14059 12597
rect 14458 12588 14464 12600
rect 14516 12588 14522 12640
rect 16022 12628 16028 12640
rect 15983 12600 16028 12628
rect 16022 12588 16028 12600
rect 16080 12588 16086 12640
rect 19518 12588 19524 12640
rect 19576 12628 19582 12640
rect 19628 12637 19656 12736
rect 19797 12733 19809 12736
rect 19843 12733 19855 12767
rect 20254 12764 20260 12776
rect 20215 12736 20260 12764
rect 19797 12727 19855 12733
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 20364 12764 20392 12804
rect 20530 12792 20536 12804
rect 20588 12792 20594 12844
rect 21361 12835 21419 12841
rect 21361 12801 21373 12835
rect 21407 12832 21419 12835
rect 21634 12832 21640 12844
rect 21407 12804 21640 12832
rect 21407 12801 21419 12804
rect 21361 12795 21419 12801
rect 21634 12792 21640 12804
rect 21692 12792 21698 12844
rect 23934 12832 23940 12844
rect 23895 12804 23940 12832
rect 23934 12792 23940 12804
rect 23992 12792 23998 12844
rect 24581 12835 24639 12841
rect 24581 12801 24593 12835
rect 24627 12832 24639 12835
rect 24670 12832 24676 12844
rect 24627 12804 24676 12832
rect 24627 12801 24639 12804
rect 24581 12795 24639 12801
rect 24670 12792 24676 12804
rect 24728 12792 24734 12844
rect 25476 12767 25534 12773
rect 20364 12736 21312 12764
rect 21284 12696 21312 12736
rect 25476 12733 25488 12767
rect 25522 12764 25534 12767
rect 25961 12767 26019 12773
rect 25961 12764 25973 12767
rect 25522 12736 25973 12764
rect 25522 12733 25534 12736
rect 25476 12727 25534 12733
rect 25961 12733 25973 12736
rect 26007 12764 26019 12767
rect 27614 12764 27620 12776
rect 26007 12736 27620 12764
rect 26007 12733 26019 12736
rect 25961 12727 26019 12733
rect 27614 12724 27620 12736
rect 27672 12724 27678 12776
rect 21682 12699 21740 12705
rect 21682 12696 21694 12699
rect 21284 12668 21694 12696
rect 21284 12640 21312 12668
rect 21682 12665 21694 12668
rect 21728 12665 21740 12699
rect 21682 12659 21740 12665
rect 22094 12656 22100 12708
rect 22152 12696 22158 12708
rect 23477 12699 23535 12705
rect 23477 12696 23489 12699
rect 22152 12668 23489 12696
rect 22152 12656 22158 12668
rect 23477 12665 23489 12668
rect 23523 12696 23535 12699
rect 24029 12699 24087 12705
rect 24029 12696 24041 12699
rect 23523 12668 24041 12696
rect 23523 12665 23535 12668
rect 23477 12659 23535 12665
rect 24029 12665 24041 12668
rect 24075 12696 24087 12699
rect 25038 12696 25044 12708
rect 24075 12668 25044 12696
rect 24075 12665 24087 12668
rect 24029 12659 24087 12665
rect 25038 12656 25044 12668
rect 25096 12656 25102 12708
rect 19613 12631 19671 12637
rect 19613 12628 19625 12631
rect 19576 12600 19625 12628
rect 19576 12588 19582 12600
rect 19613 12597 19625 12600
rect 19659 12597 19671 12631
rect 20806 12628 20812 12640
rect 20767 12600 20812 12628
rect 19613 12591 19671 12597
rect 20806 12588 20812 12600
rect 20864 12588 20870 12640
rect 21266 12628 21272 12640
rect 21227 12600 21272 12628
rect 21266 12588 21272 12600
rect 21324 12588 21330 12640
rect 22830 12588 22836 12640
rect 22888 12628 22894 12640
rect 22925 12631 22983 12637
rect 22925 12628 22937 12631
rect 22888 12600 22937 12628
rect 22888 12588 22894 12600
rect 22925 12597 22937 12600
rect 22971 12597 22983 12631
rect 22925 12591 22983 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 8159 12427 8217 12433
rect 8159 12393 8171 12427
rect 8205 12424 8217 12427
rect 8294 12424 8300 12436
rect 8205 12396 8300 12424
rect 8205 12393 8217 12396
rect 8159 12387 8217 12393
rect 8294 12384 8300 12396
rect 8352 12384 8358 12436
rect 13081 12427 13139 12433
rect 13081 12393 13093 12427
rect 13127 12424 13139 12427
rect 13538 12424 13544 12436
rect 13127 12396 13544 12424
rect 13127 12393 13139 12396
rect 13081 12387 13139 12393
rect 13538 12384 13544 12396
rect 13596 12384 13602 12436
rect 15286 12384 15292 12436
rect 15344 12424 15350 12436
rect 16758 12424 16764 12436
rect 15344 12396 15516 12424
rect 16719 12396 16764 12424
rect 15344 12384 15350 12396
rect 12526 12356 12532 12368
rect 12487 12328 12532 12356
rect 12526 12316 12532 12328
rect 12584 12316 12590 12368
rect 15488 12365 15516 12396
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 18690 12424 18696 12436
rect 18651 12396 18696 12424
rect 18690 12384 18696 12396
rect 18748 12384 18754 12436
rect 20254 12384 20260 12436
rect 20312 12424 20318 12436
rect 20625 12427 20683 12433
rect 20625 12424 20637 12427
rect 20312 12396 20637 12424
rect 20312 12384 20318 12396
rect 20625 12393 20637 12396
rect 20671 12393 20683 12427
rect 22094 12424 22100 12436
rect 22055 12396 22100 12424
rect 20625 12387 20683 12393
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 23014 12424 23020 12436
rect 22975 12396 23020 12424
rect 23014 12384 23020 12396
rect 23072 12384 23078 12436
rect 24118 12424 24124 12436
rect 24079 12396 24124 12424
rect 24118 12384 24124 12396
rect 24176 12384 24182 12436
rect 24581 12427 24639 12433
rect 24581 12393 24593 12427
rect 24627 12393 24639 12427
rect 24581 12387 24639 12393
rect 15473 12359 15531 12365
rect 15473 12325 15485 12359
rect 15519 12325 15531 12359
rect 18414 12356 18420 12368
rect 18375 12328 18420 12356
rect 15473 12319 15531 12325
rect 18414 12316 18420 12328
rect 18472 12316 18478 12368
rect 20806 12356 20812 12368
rect 19260 12328 20812 12356
rect 7926 12288 7932 12300
rect 7887 12260 7932 12288
rect 7926 12248 7932 12260
rect 7984 12248 7990 12300
rect 12069 12291 12127 12297
rect 12069 12257 12081 12291
rect 12115 12257 12127 12291
rect 12342 12288 12348 12300
rect 12303 12260 12348 12288
rect 12069 12251 12127 12257
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 12084 12220 12112 12251
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 13262 12248 13268 12300
rect 13320 12288 13326 12300
rect 13357 12291 13415 12297
rect 13357 12288 13369 12291
rect 13320 12260 13369 12288
rect 13320 12248 13326 12260
rect 13357 12257 13369 12260
rect 13403 12257 13415 12291
rect 13357 12251 13415 12257
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 13872 12260 13917 12288
rect 13872 12248 13878 12260
rect 17218 12248 17224 12300
rect 17276 12288 17282 12300
rect 19260 12297 19288 12328
rect 20806 12316 20812 12328
rect 20864 12316 20870 12368
rect 21266 12316 21272 12368
rect 21324 12356 21330 12368
rect 21498 12359 21556 12365
rect 21498 12356 21510 12359
rect 21324 12328 21510 12356
rect 21324 12316 21330 12328
rect 21498 12325 21510 12328
rect 21544 12325 21556 12359
rect 21498 12319 21556 12325
rect 21818 12316 21824 12368
rect 21876 12356 21882 12368
rect 24596 12356 24624 12387
rect 21876 12328 24624 12356
rect 21876 12316 21882 12328
rect 17681 12291 17739 12297
rect 17681 12288 17693 12291
rect 17276 12260 17693 12288
rect 17276 12248 17282 12260
rect 17681 12257 17693 12260
rect 17727 12257 17739 12291
rect 19245 12291 19303 12297
rect 19245 12288 19257 12291
rect 17681 12251 17739 12257
rect 18984 12260 19257 12288
rect 12618 12220 12624 12232
rect 11940 12192 12624 12220
rect 11940 12180 11946 12192
rect 12618 12180 12624 12192
rect 12676 12220 12682 12232
rect 14090 12220 14096 12232
rect 12676 12192 13814 12220
rect 14051 12192 14096 12220
rect 12676 12180 12682 12192
rect 13786 12152 13814 12192
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 15378 12220 15384 12232
rect 15339 12192 15384 12220
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 15562 12180 15568 12232
rect 15620 12220 15626 12232
rect 17862 12229 17868 12232
rect 15657 12223 15715 12229
rect 15657 12220 15669 12223
rect 15620 12192 15669 12220
rect 15620 12180 15626 12192
rect 15657 12189 15669 12192
rect 15703 12189 15715 12223
rect 15657 12183 15715 12189
rect 17828 12223 17868 12229
rect 17828 12189 17840 12223
rect 17828 12183 17868 12189
rect 17862 12180 17868 12183
rect 17920 12180 17926 12232
rect 18046 12220 18052 12232
rect 18007 12192 18052 12220
rect 18046 12180 18052 12192
rect 18104 12180 18110 12232
rect 18984 12164 19012 12260
rect 19245 12257 19257 12260
rect 19291 12257 19303 12291
rect 19245 12251 19303 12257
rect 19705 12291 19763 12297
rect 19705 12257 19717 12291
rect 19751 12257 19763 12291
rect 23014 12288 23020 12300
rect 22975 12260 23020 12288
rect 19705 12251 19763 12257
rect 19720 12220 19748 12251
rect 23014 12248 23020 12260
rect 23072 12248 23078 12300
rect 23198 12248 23204 12300
rect 23256 12288 23262 12300
rect 23339 12291 23397 12297
rect 23339 12288 23351 12291
rect 23256 12260 23351 12288
rect 23256 12248 23262 12260
rect 23339 12257 23351 12260
rect 23385 12257 23397 12291
rect 24670 12288 24676 12300
rect 24631 12260 24676 12288
rect 23339 12251 23397 12257
rect 24670 12248 24676 12260
rect 24728 12248 24734 12300
rect 24949 12291 25007 12297
rect 24949 12257 24961 12291
rect 24995 12257 25007 12291
rect 24949 12251 25007 12257
rect 19978 12220 19984 12232
rect 19076 12192 19748 12220
rect 19939 12192 19984 12220
rect 18966 12152 18972 12164
rect 13786 12124 18972 12152
rect 18966 12112 18972 12124
rect 19024 12112 19030 12164
rect 19076 12096 19104 12192
rect 19978 12180 19984 12192
rect 20036 12180 20042 12232
rect 20254 12180 20260 12232
rect 20312 12220 20318 12232
rect 20349 12223 20407 12229
rect 20349 12220 20361 12223
rect 20312 12192 20361 12220
rect 20312 12180 20318 12192
rect 20349 12189 20361 12192
rect 20395 12220 20407 12223
rect 21177 12223 21235 12229
rect 21177 12220 21189 12223
rect 20395 12192 21189 12220
rect 20395 12189 20407 12192
rect 20349 12183 20407 12189
rect 21177 12189 21189 12192
rect 21223 12189 21235 12223
rect 21177 12183 21235 12189
rect 20806 12112 20812 12164
rect 20864 12152 20870 12164
rect 24670 12152 24676 12164
rect 20864 12124 24676 12152
rect 20864 12112 20870 12124
rect 24670 12112 24676 12124
rect 24728 12112 24734 12164
rect 14550 12084 14556 12096
rect 14511 12056 14556 12084
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 14826 12044 14832 12096
rect 14884 12084 14890 12096
rect 14921 12087 14979 12093
rect 14921 12084 14933 12087
rect 14884 12056 14933 12084
rect 14884 12044 14890 12056
rect 14921 12053 14933 12056
rect 14967 12053 14979 12087
rect 14921 12047 14979 12053
rect 15746 12044 15752 12096
rect 15804 12084 15810 12096
rect 16301 12087 16359 12093
rect 16301 12084 16313 12087
rect 15804 12056 16313 12084
rect 15804 12044 15810 12056
rect 16301 12053 16313 12056
rect 16347 12053 16359 12087
rect 16301 12047 16359 12053
rect 17589 12087 17647 12093
rect 17589 12053 17601 12087
rect 17635 12084 17647 12087
rect 17954 12084 17960 12096
rect 17635 12056 17960 12084
rect 17635 12053 17647 12056
rect 17589 12047 17647 12053
rect 17954 12044 17960 12056
rect 18012 12044 18018 12096
rect 19058 12084 19064 12096
rect 19019 12056 19064 12084
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 23198 12044 23204 12096
rect 23256 12084 23262 12096
rect 24964 12084 24992 12251
rect 25038 12084 25044 12096
rect 23256 12056 25044 12084
rect 23256 12044 23262 12056
rect 25038 12044 25044 12056
rect 25096 12044 25102 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 11882 11880 11888 11892
rect 11843 11852 11888 11880
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 12989 11883 13047 11889
rect 12989 11849 13001 11883
rect 13035 11880 13047 11883
rect 13814 11880 13820 11892
rect 13035 11852 13820 11880
rect 13035 11849 13047 11852
rect 12989 11843 13047 11849
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 15378 11840 15384 11892
rect 15436 11880 15442 11892
rect 16577 11883 16635 11889
rect 16577 11880 16589 11883
rect 15436 11852 16589 11880
rect 15436 11840 15442 11852
rect 16577 11849 16589 11852
rect 16623 11849 16635 11883
rect 20990 11880 20996 11892
rect 16577 11843 16635 11849
rect 16684 11852 20996 11880
rect 11974 11772 11980 11824
rect 12032 11812 12038 11824
rect 14550 11812 14556 11824
rect 12032 11784 14556 11812
rect 12032 11772 12038 11784
rect 14550 11772 14556 11784
rect 14608 11812 14614 11824
rect 14737 11815 14795 11821
rect 14737 11812 14749 11815
rect 14608 11784 14749 11812
rect 14608 11772 14614 11784
rect 14737 11781 14749 11784
rect 14783 11781 14795 11815
rect 14737 11775 14795 11781
rect 15473 11815 15531 11821
rect 15473 11781 15485 11815
rect 15519 11812 15531 11815
rect 16684 11812 16712 11852
rect 20990 11840 20996 11852
rect 21048 11840 21054 11892
rect 22002 11880 22008 11892
rect 21963 11852 22008 11880
rect 22002 11840 22008 11852
rect 22060 11840 22066 11892
rect 23382 11880 23388 11892
rect 23343 11852 23388 11880
rect 23382 11840 23388 11852
rect 23440 11840 23446 11892
rect 24670 11880 24676 11892
rect 24631 11852 24676 11880
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 25038 11880 25044 11892
rect 24999 11852 25044 11880
rect 25038 11840 25044 11852
rect 25096 11840 25102 11892
rect 25774 11880 25780 11892
rect 25735 11852 25780 11880
rect 25774 11840 25780 11852
rect 25832 11840 25838 11892
rect 15519 11784 16712 11812
rect 15519 11781 15531 11784
rect 15473 11775 15531 11781
rect 16850 11772 16856 11824
rect 16908 11812 16914 11824
rect 22557 11815 22615 11821
rect 22557 11812 22569 11815
rect 16908 11784 22569 11812
rect 16908 11772 16914 11784
rect 22557 11781 22569 11784
rect 22603 11812 22615 11815
rect 23198 11812 23204 11824
rect 22603 11784 23204 11812
rect 22603 11781 22615 11784
rect 22557 11775 22615 11781
rect 23198 11772 23204 11784
rect 23256 11772 23262 11824
rect 23566 11772 23572 11824
rect 23624 11812 23630 11824
rect 25363 11815 25421 11821
rect 25363 11812 25375 11815
rect 23624 11784 25375 11812
rect 23624 11772 23630 11784
rect 25363 11781 25375 11784
rect 25409 11781 25421 11815
rect 25363 11775 25421 11781
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11744 11575 11747
rect 13630 11744 13636 11756
rect 11563 11716 13636 11744
rect 11563 11713 11575 11716
rect 11517 11707 11575 11713
rect 13630 11704 13636 11716
rect 13688 11704 13694 11756
rect 14826 11704 14832 11756
rect 14884 11744 14890 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 14884 11716 15945 11744
rect 14884 11704 14890 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 18966 11744 18972 11756
rect 18927 11716 18972 11744
rect 15933 11707 15991 11713
rect 18966 11704 18972 11716
rect 19024 11704 19030 11756
rect 20254 11744 20260 11756
rect 20215 11716 20260 11744
rect 20254 11704 20260 11716
rect 20312 11704 20318 11756
rect 23934 11704 23940 11756
rect 23992 11744 23998 11756
rect 24029 11747 24087 11753
rect 24029 11744 24041 11747
rect 23992 11716 24041 11744
rect 23992 11704 23998 11716
rect 24029 11713 24041 11716
rect 24075 11713 24087 11747
rect 24029 11707 24087 11713
rect 10689 11679 10747 11685
rect 10689 11645 10701 11679
rect 10735 11676 10747 11679
rect 11425 11679 11483 11685
rect 11425 11676 11437 11679
rect 10735 11648 11437 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 11425 11645 11437 11648
rect 11471 11676 11483 11679
rect 13446 11676 13452 11688
rect 11471 11648 13452 11676
rect 11471 11645 11483 11648
rect 11425 11639 11483 11645
rect 13446 11636 13452 11648
rect 13504 11636 13510 11688
rect 13817 11679 13875 11685
rect 13817 11645 13829 11679
rect 13863 11676 13875 11679
rect 14090 11676 14096 11688
rect 13863 11648 14096 11676
rect 13863 11645 13875 11648
rect 13817 11639 13875 11645
rect 14090 11636 14096 11648
rect 14148 11676 14154 11688
rect 14550 11676 14556 11688
rect 14148 11648 14556 11676
rect 14148 11636 14154 11648
rect 14550 11636 14556 11648
rect 14608 11636 14614 11688
rect 18049 11679 18107 11685
rect 18049 11645 18061 11679
rect 18095 11676 18107 11679
rect 18095 11648 18644 11676
rect 18095 11645 18107 11648
rect 18049 11639 18107 11645
rect 12253 11611 12311 11617
rect 12253 11577 12265 11611
rect 12299 11608 12311 11611
rect 12342 11608 12348 11620
rect 12299 11580 12348 11608
rect 12299 11577 12311 11580
rect 12253 11571 12311 11577
rect 12342 11568 12348 11580
rect 12400 11608 12406 11620
rect 13538 11608 13544 11620
rect 12400 11580 13544 11608
rect 12400 11568 12406 11580
rect 13538 11568 13544 11580
rect 13596 11568 13602 11620
rect 14179 11611 14237 11617
rect 14179 11608 14191 11611
rect 13740 11580 14191 11608
rect 13740 11552 13768 11580
rect 14179 11577 14191 11580
rect 14225 11577 14237 11611
rect 14179 11571 14237 11577
rect 15102 11568 15108 11620
rect 15160 11608 15166 11620
rect 15473 11611 15531 11617
rect 15473 11608 15485 11611
rect 15160 11580 15485 11608
rect 15160 11568 15166 11580
rect 15473 11577 15485 11580
rect 15519 11608 15531 11611
rect 15646 11611 15704 11617
rect 15646 11608 15658 11611
rect 15519 11580 15658 11608
rect 15519 11577 15531 11580
rect 15473 11571 15531 11577
rect 15646 11577 15658 11580
rect 15692 11577 15704 11611
rect 15646 11571 15704 11577
rect 15746 11568 15752 11620
rect 15804 11608 15810 11620
rect 17313 11611 17371 11617
rect 15804 11580 15849 11608
rect 15804 11568 15810 11580
rect 17313 11577 17325 11611
rect 17359 11608 17371 11611
rect 17862 11608 17868 11620
rect 17359 11580 17868 11608
rect 17359 11577 17371 11580
rect 17313 11571 17371 11577
rect 17862 11568 17868 11580
rect 17920 11608 17926 11620
rect 17920 11580 18276 11608
rect 17920 11568 17926 11580
rect 6914 11500 6920 11552
rect 6972 11540 6978 11552
rect 7926 11540 7932 11552
rect 6972 11512 7932 11540
rect 6972 11500 6978 11512
rect 7926 11500 7932 11512
rect 7984 11540 7990 11552
rect 8021 11543 8079 11549
rect 8021 11540 8033 11543
rect 7984 11512 8033 11540
rect 7984 11500 7990 11512
rect 8021 11509 8033 11512
rect 8067 11509 8079 11543
rect 13262 11540 13268 11552
rect 13223 11512 13268 11540
rect 8021 11503 8079 11509
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 13722 11540 13728 11552
rect 13683 11512 13728 11540
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 15286 11540 15292 11552
rect 15247 11512 15292 11540
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 17037 11543 17095 11549
rect 17037 11509 17049 11543
rect 17083 11540 17095 11543
rect 17218 11540 17224 11552
rect 17083 11512 17224 11540
rect 17083 11509 17095 11512
rect 17037 11503 17095 11509
rect 17218 11500 17224 11512
rect 17276 11500 17282 11552
rect 17773 11543 17831 11549
rect 17773 11509 17785 11543
rect 17819 11540 17831 11543
rect 18046 11540 18052 11552
rect 17819 11512 18052 11540
rect 17819 11509 17831 11512
rect 17773 11503 17831 11509
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 18248 11549 18276 11580
rect 18616 11549 18644 11648
rect 19150 11636 19156 11688
rect 19208 11676 19214 11688
rect 19518 11676 19524 11688
rect 19208 11648 19524 11676
rect 19208 11636 19214 11648
rect 19518 11636 19524 11648
rect 19576 11636 19582 11688
rect 19981 11679 20039 11685
rect 19981 11645 19993 11679
rect 20027 11645 20039 11679
rect 21082 11676 21088 11688
rect 21043 11648 21088 11676
rect 19981 11639 20039 11645
rect 19058 11568 19064 11620
rect 19116 11608 19122 11620
rect 19996 11608 20024 11639
rect 21082 11636 21088 11648
rect 21140 11636 21146 11688
rect 25292 11679 25350 11685
rect 25292 11645 25304 11679
rect 25338 11676 25350 11679
rect 25774 11676 25780 11688
rect 25338 11648 25780 11676
rect 25338 11645 25350 11648
rect 25292 11639 25350 11645
rect 25774 11636 25780 11648
rect 25832 11636 25838 11688
rect 19116 11580 20024 11608
rect 20088 11580 21036 11608
rect 19116 11568 19122 11580
rect 18233 11543 18291 11549
rect 18233 11509 18245 11543
rect 18279 11509 18291 11543
rect 18233 11503 18291 11509
rect 18601 11543 18659 11549
rect 18601 11509 18613 11543
rect 18647 11540 18659 11543
rect 18782 11540 18788 11552
rect 18647 11512 18788 11540
rect 18647 11509 18659 11512
rect 18601 11503 18659 11509
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 19150 11500 19156 11552
rect 19208 11540 19214 11552
rect 19337 11543 19395 11549
rect 19337 11540 19349 11543
rect 19208 11512 19349 11540
rect 19208 11500 19214 11512
rect 19337 11509 19349 11512
rect 19383 11540 19395 11543
rect 20088 11540 20116 11580
rect 20622 11540 20628 11552
rect 19383 11512 20116 11540
rect 20583 11512 20628 11540
rect 19383 11509 19395 11512
rect 19337 11503 19395 11509
rect 20622 11500 20628 11512
rect 20680 11540 20686 11552
rect 20901 11543 20959 11549
rect 20901 11540 20913 11543
rect 20680 11512 20913 11540
rect 20680 11500 20686 11512
rect 20901 11509 20913 11512
rect 20947 11509 20959 11543
rect 21008 11540 21036 11580
rect 21266 11568 21272 11620
rect 21324 11608 21330 11620
rect 21406 11611 21464 11617
rect 21406 11608 21418 11611
rect 21324 11580 21418 11608
rect 21324 11568 21330 11580
rect 21406 11577 21418 11580
rect 21452 11577 21464 11611
rect 23750 11608 23756 11620
rect 23711 11580 23756 11608
rect 21406 11571 21464 11577
rect 23750 11568 23756 11580
rect 23808 11568 23814 11620
rect 23845 11611 23903 11617
rect 23845 11577 23857 11611
rect 23891 11577 23903 11611
rect 23845 11571 23903 11577
rect 22925 11543 22983 11549
rect 22925 11540 22937 11543
rect 21008 11512 22937 11540
rect 20901 11503 20959 11509
rect 22925 11509 22937 11512
rect 22971 11540 22983 11543
rect 23014 11540 23020 11552
rect 22971 11512 23020 11540
rect 22971 11509 22983 11512
rect 22925 11503 22983 11509
rect 23014 11500 23020 11512
rect 23072 11500 23078 11552
rect 23382 11500 23388 11552
rect 23440 11540 23446 11552
rect 23860 11540 23888 11571
rect 23440 11512 23888 11540
rect 23440 11500 23446 11512
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 14550 11336 14556 11348
rect 12124 11308 14365 11336
rect 14511 11308 14556 11336
rect 12124 11296 12130 11308
rect 12802 11228 12808 11280
rect 12860 11268 12866 11280
rect 13722 11277 13728 11280
rect 13678 11271 13728 11277
rect 13678 11268 13690 11271
rect 12860 11240 13690 11268
rect 12860 11228 12866 11240
rect 13678 11237 13690 11240
rect 13724 11237 13728 11271
rect 13678 11231 13728 11237
rect 13722 11228 13728 11231
rect 13780 11228 13786 11280
rect 14337 11268 14365 11308
rect 14550 11296 14556 11308
rect 14608 11296 14614 11348
rect 15102 11336 15108 11348
rect 15063 11308 15108 11336
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 17034 11336 17040 11348
rect 15580 11308 17040 11336
rect 15580 11268 15608 11308
rect 17034 11296 17040 11308
rect 17092 11336 17098 11348
rect 17497 11339 17555 11345
rect 17497 11336 17509 11339
rect 17092 11308 17509 11336
rect 17092 11296 17098 11308
rect 17497 11305 17509 11308
rect 17543 11336 17555 11339
rect 17543 11308 17724 11336
rect 17543 11305 17555 11308
rect 17497 11299 17555 11305
rect 16850 11268 16856 11280
rect 14337 11240 15608 11268
rect 16811 11240 16856 11268
rect 11882 11200 11888 11212
rect 11843 11172 11888 11200
rect 11882 11160 11888 11172
rect 11940 11160 11946 11212
rect 12529 11203 12587 11209
rect 12529 11169 12541 11203
rect 12575 11200 12587 11203
rect 15286 11200 15292 11212
rect 12575 11172 15292 11200
rect 12575 11169 12587 11172
rect 12529 11163 12587 11169
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 15580 11200 15608 11240
rect 16850 11228 16856 11240
rect 16908 11228 16914 11280
rect 17696 11277 17724 11308
rect 19978 11296 19984 11348
rect 20036 11336 20042 11348
rect 20625 11339 20683 11345
rect 20625 11336 20637 11339
rect 20036 11308 20637 11336
rect 20036 11296 20042 11308
rect 20625 11305 20637 11308
rect 20671 11336 20683 11339
rect 21082 11336 21088 11348
rect 20671 11308 21088 11336
rect 20671 11305 20683 11308
rect 20625 11299 20683 11305
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 21174 11296 21180 11348
rect 21232 11336 21238 11348
rect 21232 11308 21277 11336
rect 21232 11296 21238 11308
rect 17681 11271 17739 11277
rect 17681 11237 17693 11271
rect 17727 11237 17739 11271
rect 17681 11231 17739 11237
rect 18417 11271 18475 11277
rect 18417 11237 18429 11271
rect 18463 11268 18475 11271
rect 19058 11268 19064 11280
rect 18463 11240 19064 11268
rect 18463 11237 18475 11240
rect 18417 11231 18475 11237
rect 19058 11228 19064 11240
rect 19116 11268 19122 11280
rect 20257 11271 20315 11277
rect 20257 11268 20269 11271
rect 19116 11240 20269 11268
rect 19116 11228 19122 11240
rect 20257 11237 20269 11240
rect 20303 11237 20315 11271
rect 20257 11231 20315 11237
rect 20364 11240 21496 11268
rect 15933 11203 15991 11209
rect 15933 11200 15945 11203
rect 15580 11172 15945 11200
rect 15933 11169 15945 11172
rect 15979 11169 15991 11203
rect 15933 11163 15991 11169
rect 19150 11160 19156 11212
rect 19208 11200 19214 11212
rect 19245 11203 19303 11209
rect 19245 11200 19257 11203
rect 19208 11172 19257 11200
rect 19208 11160 19214 11172
rect 19245 11169 19257 11172
rect 19291 11169 19303 11203
rect 19245 11163 19303 11169
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 19797 11203 19855 11209
rect 19797 11200 19809 11203
rect 19392 11172 19809 11200
rect 19392 11160 19398 11172
rect 19797 11169 19809 11172
rect 19843 11200 19855 11203
rect 20364 11200 20392 11240
rect 21468 11212 21496 11240
rect 22002 11228 22008 11280
rect 22060 11268 22066 11280
rect 23661 11271 23719 11277
rect 23661 11268 23673 11271
rect 22060 11240 23673 11268
rect 22060 11228 22066 11240
rect 23661 11237 23673 11240
rect 23707 11237 23719 11271
rect 25314 11268 25320 11280
rect 23661 11231 23719 11237
rect 25123 11240 25320 11268
rect 19843 11172 20392 11200
rect 19843 11169 19855 11172
rect 19797 11163 19855 11169
rect 20806 11160 20812 11212
rect 20864 11200 20870 11212
rect 20901 11203 20959 11209
rect 20901 11200 20913 11203
rect 20864 11172 20913 11200
rect 20864 11160 20870 11172
rect 20901 11169 20913 11172
rect 20947 11169 20959 11203
rect 21450 11200 21456 11212
rect 21411 11172 21456 11200
rect 20901 11163 20959 11169
rect 21450 11160 21456 11172
rect 21508 11160 21514 11212
rect 25123 11209 25151 11240
rect 25314 11228 25320 11240
rect 25372 11228 25378 11280
rect 25108 11203 25166 11209
rect 25108 11169 25120 11203
rect 25154 11169 25166 11203
rect 25108 11163 25166 11169
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 13170 10996 13176 11008
rect 13131 10968 13176 10996
rect 13170 10956 13176 10968
rect 13228 10996 13234 11008
rect 13372 10996 13400 11095
rect 16206 11092 16212 11144
rect 16264 11132 16270 11144
rect 16485 11135 16543 11141
rect 16264 11104 16436 11132
rect 16264 11092 16270 11104
rect 13446 11024 13452 11076
rect 13504 11064 13510 11076
rect 14277 11067 14335 11073
rect 14277 11064 14289 11067
rect 13504 11036 14289 11064
rect 13504 11024 13510 11036
rect 14277 11033 14289 11036
rect 14323 11064 14335 11067
rect 15746 11064 15752 11076
rect 14323 11036 15752 11064
rect 14323 11033 14335 11036
rect 14277 11027 14335 11033
rect 15746 11024 15752 11036
rect 15804 11024 15810 11076
rect 16408 11073 16436 11104
rect 16485 11101 16497 11135
rect 16531 11132 16543 11135
rect 16574 11132 16580 11144
rect 16531 11104 16580 11132
rect 16531 11101 16543 11104
rect 16485 11095 16543 11101
rect 16574 11092 16580 11104
rect 16632 11092 16638 11144
rect 18046 11132 18052 11144
rect 18007 11104 18052 11132
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 19981 11135 20039 11141
rect 19981 11101 19993 11135
rect 20027 11132 20039 11135
rect 21082 11132 21088 11144
rect 20027 11104 21088 11132
rect 20027 11101 20039 11104
rect 19981 11095 20039 11101
rect 21082 11092 21088 11104
rect 21140 11092 21146 11144
rect 22465 11135 22523 11141
rect 22465 11101 22477 11135
rect 22511 11132 22523 11135
rect 23014 11132 23020 11144
rect 22511 11104 23020 11132
rect 22511 11101 22523 11104
rect 22465 11095 22523 11101
rect 23014 11092 23020 11104
rect 23072 11092 23078 11144
rect 23566 11132 23572 11144
rect 23527 11104 23572 11132
rect 23566 11092 23572 11104
rect 23624 11092 23630 11144
rect 23934 11132 23940 11144
rect 23895 11104 23940 11132
rect 23934 11092 23940 11104
rect 23992 11092 23998 11144
rect 16393 11067 16451 11073
rect 16393 11033 16405 11067
rect 16439 11033 16451 11067
rect 17954 11064 17960 11076
rect 17867 11036 17960 11064
rect 16393 11027 16451 11033
rect 17954 11024 17960 11036
rect 18012 11064 18018 11076
rect 19061 11067 19119 11073
rect 19061 11064 19073 11067
rect 18012 11036 19073 11064
rect 18012 11024 18018 11036
rect 19061 11033 19073 11036
rect 19107 11033 19119 11067
rect 21100 11064 21128 11092
rect 21913 11067 21971 11073
rect 21913 11064 21925 11067
rect 21100 11036 21925 11064
rect 19061 11027 19119 11033
rect 21913 11033 21925 11036
rect 21959 11033 21971 11067
rect 21913 11027 21971 11033
rect 15562 10996 15568 11008
rect 13228 10968 13400 10996
rect 15523 10968 15568 10996
rect 13228 10956 13234 10968
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 16298 11005 16304 11008
rect 16282 10999 16304 11005
rect 16282 10965 16294 10999
rect 16282 10959 16304 10965
rect 16298 10956 16304 10959
rect 16356 10956 16362 11008
rect 17218 10996 17224 11008
rect 17179 10968 17224 10996
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 17862 11005 17868 11008
rect 17846 10999 17868 11005
rect 17846 10965 17858 10999
rect 17846 10959 17868 10965
rect 17862 10956 17868 10959
rect 17920 10956 17926 11008
rect 18322 10956 18328 11008
rect 18380 10996 18386 11008
rect 18693 10999 18751 11005
rect 18693 10996 18705 10999
rect 18380 10968 18705 10996
rect 18380 10956 18386 10968
rect 18693 10965 18705 10968
rect 18739 10965 18751 10999
rect 18693 10959 18751 10965
rect 23750 10956 23756 11008
rect 23808 10996 23814 11008
rect 24489 10999 24547 11005
rect 24489 10996 24501 10999
rect 23808 10968 24501 10996
rect 23808 10956 23814 10968
rect 24489 10965 24501 10968
rect 24535 10965 24547 10999
rect 24489 10959 24547 10965
rect 24670 10956 24676 11008
rect 24728 10996 24734 11008
rect 25179 10999 25237 11005
rect 25179 10996 25191 10999
rect 24728 10968 25191 10996
rect 24728 10956 24734 10968
rect 25179 10965 25191 10968
rect 25225 10965 25237 10999
rect 25179 10959 25237 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 11882 10792 11888 10804
rect 11843 10764 11888 10792
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 12526 10752 12532 10804
rect 12584 10792 12590 10804
rect 12584 10764 15884 10792
rect 12584 10752 12590 10764
rect 12618 10724 12624 10736
rect 12579 10696 12624 10724
rect 12618 10684 12624 10696
rect 12676 10684 12682 10736
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10656 14243 10659
rect 14826 10656 14832 10668
rect 14231 10628 14832 10656
rect 14231 10625 14243 10628
rect 14185 10619 14243 10625
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 7352 10591 7410 10597
rect 7352 10557 7364 10591
rect 7398 10588 7410 10591
rect 12437 10591 12495 10597
rect 7398 10560 7788 10588
rect 7398 10557 7410 10560
rect 7352 10551 7410 10557
rect 7760 10464 7788 10560
rect 12437 10557 12449 10591
rect 12483 10588 12495 10591
rect 12894 10588 12900 10600
rect 12483 10560 12900 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 12894 10548 12900 10560
rect 12952 10548 12958 10600
rect 15286 10588 15292 10600
rect 15247 10560 15292 10588
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 15856 10597 15884 10764
rect 16666 10752 16672 10804
rect 16724 10792 16730 10804
rect 16761 10795 16819 10801
rect 16761 10792 16773 10795
rect 16724 10764 16773 10792
rect 16724 10752 16730 10764
rect 16761 10761 16773 10764
rect 16807 10761 16819 10795
rect 16761 10755 16819 10761
rect 20625 10795 20683 10801
rect 20625 10761 20637 10795
rect 20671 10792 20683 10795
rect 20806 10792 20812 10804
rect 20671 10764 20812 10792
rect 20671 10761 20683 10764
rect 20625 10755 20683 10761
rect 20806 10752 20812 10764
rect 20864 10752 20870 10804
rect 21450 10752 21456 10804
rect 21508 10792 21514 10804
rect 22281 10795 22339 10801
rect 22281 10792 22293 10795
rect 21508 10764 22293 10792
rect 21508 10752 21514 10764
rect 22281 10761 22293 10764
rect 22327 10761 22339 10795
rect 23014 10792 23020 10804
rect 22975 10764 23020 10792
rect 22281 10755 22339 10761
rect 23014 10752 23020 10764
rect 23072 10752 23078 10804
rect 25133 10795 25191 10801
rect 25133 10761 25145 10795
rect 25179 10792 25191 10795
rect 25314 10792 25320 10804
rect 25179 10764 25320 10792
rect 25179 10761 25191 10764
rect 25133 10755 25191 10761
rect 25314 10752 25320 10764
rect 25372 10752 25378 10804
rect 15933 10727 15991 10733
rect 15933 10693 15945 10727
rect 15979 10724 15991 10727
rect 16577 10727 16635 10733
rect 16577 10724 16589 10727
rect 15979 10696 16589 10724
rect 15979 10693 15991 10696
rect 15933 10687 15991 10693
rect 16577 10693 16589 10696
rect 16623 10724 16635 10727
rect 17954 10724 17960 10736
rect 16623 10696 17960 10724
rect 16623 10693 16635 10696
rect 16577 10687 16635 10693
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 18322 10724 18328 10736
rect 18283 10696 18328 10724
rect 18322 10684 18328 10696
rect 18380 10684 18386 10736
rect 19797 10727 19855 10733
rect 19797 10724 19809 10727
rect 18432 10696 19809 10724
rect 16666 10656 16672 10668
rect 16627 10628 16672 10656
rect 16666 10616 16672 10628
rect 16724 10616 16730 10668
rect 17678 10616 17684 10668
rect 17736 10656 17742 10668
rect 18046 10656 18052 10668
rect 17736 10628 18052 10656
rect 17736 10616 17742 10628
rect 18046 10616 18052 10628
rect 18104 10656 18110 10668
rect 18432 10665 18460 10696
rect 19797 10693 19809 10696
rect 19843 10693 19855 10727
rect 19797 10687 19855 10693
rect 22002 10684 22008 10736
rect 22060 10724 22066 10736
rect 22649 10727 22707 10733
rect 22649 10724 22661 10727
rect 22060 10696 22661 10724
rect 22060 10684 22066 10696
rect 22649 10693 22661 10696
rect 22695 10693 22707 10727
rect 22649 10687 22707 10693
rect 18417 10659 18475 10665
rect 18417 10656 18429 10659
rect 18104 10628 18429 10656
rect 18104 10616 18110 10628
rect 18417 10625 18429 10628
rect 18463 10625 18475 10659
rect 18417 10619 18475 10625
rect 18785 10659 18843 10665
rect 18785 10625 18797 10659
rect 18831 10656 18843 10659
rect 19334 10656 19340 10668
rect 18831 10628 19340 10656
rect 18831 10625 18843 10628
rect 18785 10619 18843 10625
rect 19334 10616 19340 10628
rect 19392 10616 19398 10668
rect 21082 10656 21088 10668
rect 21043 10628 21088 10656
rect 21082 10616 21088 10628
rect 21140 10616 21146 10668
rect 23032 10656 23060 10752
rect 23474 10724 23480 10736
rect 23435 10696 23480 10724
rect 23474 10684 23480 10696
rect 23532 10684 23538 10736
rect 23566 10684 23572 10736
rect 23624 10724 23630 10736
rect 24670 10724 24676 10736
rect 23624 10696 24676 10724
rect 23624 10684 23630 10696
rect 24670 10684 24676 10696
rect 24728 10684 24734 10736
rect 23753 10659 23811 10665
rect 23753 10656 23765 10659
rect 23032 10628 23765 10656
rect 23753 10625 23765 10628
rect 23799 10625 23811 10659
rect 24026 10656 24032 10668
rect 23987 10628 24032 10656
rect 23753 10619 23811 10625
rect 24026 10616 24032 10628
rect 24084 10616 24090 10668
rect 15841 10591 15899 10597
rect 15841 10557 15853 10591
rect 15887 10588 15899 10591
rect 16448 10591 16506 10597
rect 16448 10588 16460 10591
rect 15887 10560 16460 10588
rect 15887 10557 15899 10560
rect 15841 10551 15899 10557
rect 16448 10557 16460 10560
rect 16494 10588 16506 10591
rect 16494 10560 17080 10588
rect 16494 10557 16506 10560
rect 16448 10551 16506 10557
rect 12986 10480 12992 10532
rect 13044 10520 13050 10532
rect 13541 10523 13599 10529
rect 13541 10520 13553 10523
rect 13044 10492 13553 10520
rect 13044 10480 13050 10492
rect 13541 10489 13553 10492
rect 13587 10489 13599 10523
rect 13541 10483 13599 10489
rect 13630 10480 13636 10532
rect 13688 10520 13694 10532
rect 15197 10523 15255 10529
rect 13688 10492 13814 10520
rect 13688 10480 13694 10492
rect 7423 10455 7481 10461
rect 7423 10421 7435 10455
rect 7469 10452 7481 10455
rect 7558 10452 7564 10464
rect 7469 10424 7564 10452
rect 7469 10421 7481 10424
rect 7423 10415 7481 10421
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 7742 10452 7748 10464
rect 7703 10424 7748 10452
rect 7742 10412 7748 10424
rect 7800 10412 7806 10464
rect 12250 10412 12256 10464
rect 12308 10452 12314 10464
rect 12802 10452 12808 10464
rect 12308 10424 12808 10452
rect 12308 10412 12314 10424
rect 12802 10412 12808 10424
rect 12860 10452 12866 10464
rect 13265 10455 13323 10461
rect 13265 10452 13277 10455
rect 12860 10424 13277 10452
rect 12860 10412 12866 10424
rect 13265 10421 13277 10424
rect 13311 10421 13323 10455
rect 13786 10452 13814 10492
rect 15197 10489 15209 10523
rect 15243 10520 15255 10523
rect 15930 10520 15936 10532
rect 15243 10492 15936 10520
rect 15243 10489 15255 10492
rect 15197 10483 15255 10489
rect 15930 10480 15936 10492
rect 15988 10480 15994 10532
rect 16301 10523 16359 10529
rect 16301 10489 16313 10523
rect 16347 10489 16359 10523
rect 17052 10520 17080 10560
rect 17862 10548 17868 10600
rect 17920 10588 17926 10600
rect 18196 10591 18254 10597
rect 18196 10588 18208 10591
rect 17920 10560 18208 10588
rect 17920 10548 17926 10560
rect 18196 10557 18208 10560
rect 18242 10557 18254 10591
rect 18196 10551 18254 10557
rect 18690 10548 18696 10600
rect 18748 10588 18754 10600
rect 19613 10591 19671 10597
rect 19613 10588 19625 10591
rect 18748 10560 19625 10588
rect 18748 10548 18754 10560
rect 19613 10557 19625 10560
rect 19659 10588 19671 10591
rect 20073 10591 20131 10597
rect 20073 10588 20085 10591
rect 19659 10560 20085 10588
rect 19659 10557 19671 10560
rect 19613 10551 19671 10557
rect 20073 10557 20085 10560
rect 20119 10557 20131 10591
rect 20073 10551 20131 10557
rect 22005 10591 22063 10597
rect 22005 10557 22017 10591
rect 22051 10588 22063 10591
rect 23290 10588 23296 10600
rect 22051 10560 23296 10588
rect 22051 10557 22063 10560
rect 22005 10551 22063 10557
rect 23290 10548 23296 10560
rect 23348 10548 23354 10600
rect 18046 10520 18052 10532
rect 17052 10492 17816 10520
rect 17959 10492 18052 10520
rect 16301 10483 16359 10489
rect 14461 10455 14519 10461
rect 14461 10452 14473 10455
rect 13786 10424 14473 10452
rect 13265 10415 13323 10421
rect 14461 10421 14473 10424
rect 14507 10421 14519 10455
rect 15470 10452 15476 10464
rect 15431 10424 15476 10452
rect 14461 10415 14519 10421
rect 15470 10412 15476 10424
rect 15528 10412 15534 10464
rect 16206 10452 16212 10464
rect 16167 10424 16212 10452
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 16316 10452 16344 10483
rect 17218 10452 17224 10464
rect 16316 10424 17224 10452
rect 17218 10412 17224 10424
rect 17276 10412 17282 10464
rect 17405 10455 17463 10461
rect 17405 10421 17417 10455
rect 17451 10452 17463 10455
rect 17678 10452 17684 10464
rect 17451 10424 17684 10452
rect 17451 10421 17463 10424
rect 17405 10415 17463 10421
rect 17678 10412 17684 10424
rect 17736 10412 17742 10464
rect 17788 10452 17816 10492
rect 18046 10480 18052 10492
rect 18104 10520 18110 10532
rect 19058 10520 19064 10532
rect 18104 10492 19064 10520
rect 18104 10480 18110 10492
rect 19058 10480 19064 10492
rect 19116 10480 19122 10532
rect 21406 10523 21464 10529
rect 21406 10520 21418 10523
rect 21284 10492 21418 10520
rect 21284 10464 21312 10492
rect 21406 10489 21418 10492
rect 21452 10489 21464 10523
rect 21406 10483 21464 10489
rect 23474 10480 23480 10532
rect 23532 10520 23538 10532
rect 23845 10523 23903 10529
rect 23845 10520 23857 10523
rect 23532 10492 23857 10520
rect 23532 10480 23538 10492
rect 23845 10489 23857 10492
rect 23891 10489 23903 10523
rect 23845 10483 23903 10489
rect 18782 10452 18788 10464
rect 17788 10424 18788 10452
rect 18782 10412 18788 10424
rect 18840 10412 18846 10464
rect 19150 10412 19156 10464
rect 19208 10452 19214 10464
rect 19245 10455 19303 10461
rect 19245 10452 19257 10455
rect 19208 10424 19257 10452
rect 19208 10412 19214 10424
rect 19245 10421 19257 10424
rect 19291 10421 19303 10455
rect 19245 10415 19303 10421
rect 20622 10412 20628 10464
rect 20680 10452 20686 10464
rect 20993 10455 21051 10461
rect 20993 10452 21005 10455
rect 20680 10424 21005 10452
rect 20680 10412 20686 10424
rect 20993 10421 21005 10424
rect 21039 10452 21051 10455
rect 21266 10452 21272 10464
rect 21039 10424 21272 10452
rect 21039 10421 21051 10424
rect 20993 10415 21051 10421
rect 21266 10412 21272 10424
rect 21324 10412 21330 10464
rect 25222 10452 25228 10464
rect 25183 10424 25228 10452
rect 25222 10412 25228 10424
rect 25280 10412 25286 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 7558 10208 7564 10260
rect 7616 10248 7622 10260
rect 12897 10251 12955 10257
rect 12897 10248 12909 10251
rect 7616 10220 12909 10248
rect 7616 10208 7622 10220
rect 12897 10217 12909 10220
rect 12943 10248 12955 10251
rect 12986 10248 12992 10260
rect 12943 10220 12992 10248
rect 12943 10217 12955 10220
rect 12897 10211 12955 10217
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 13170 10248 13176 10260
rect 13131 10220 13176 10248
rect 13170 10208 13176 10220
rect 13228 10208 13234 10260
rect 14734 10208 14740 10260
rect 14792 10248 14798 10260
rect 17218 10248 17224 10260
rect 14792 10220 17224 10248
rect 14792 10208 14798 10220
rect 17218 10208 17224 10220
rect 17276 10248 17282 10260
rect 18046 10248 18052 10260
rect 17276 10220 18052 10248
rect 17276 10208 17282 10220
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 19245 10251 19303 10257
rect 19245 10217 19257 10251
rect 19291 10248 19303 10251
rect 19334 10248 19340 10260
rect 19291 10220 19340 10248
rect 19291 10217 19303 10220
rect 19245 10211 19303 10217
rect 19334 10208 19340 10220
rect 19392 10208 19398 10260
rect 21266 10248 21272 10260
rect 21227 10220 21272 10248
rect 21266 10208 21272 10220
rect 21324 10208 21330 10260
rect 21726 10208 21732 10260
rect 21784 10248 21790 10260
rect 21821 10251 21879 10257
rect 21821 10248 21833 10251
rect 21784 10220 21833 10248
rect 21784 10208 21790 10220
rect 21821 10217 21833 10220
rect 21867 10217 21879 10251
rect 21821 10211 21879 10217
rect 23290 10208 23296 10260
rect 23348 10248 23354 10260
rect 23348 10220 23520 10248
rect 23348 10208 23354 10220
rect 11517 10183 11575 10189
rect 11517 10149 11529 10183
rect 11563 10180 11575 10183
rect 12066 10180 12072 10192
rect 11563 10152 12072 10180
rect 11563 10149 11575 10152
rect 11517 10143 11575 10149
rect 12066 10140 12072 10152
rect 12124 10140 12130 10192
rect 12710 10140 12716 10192
rect 12768 10180 12774 10192
rect 12768 10152 13124 10180
rect 12768 10140 12774 10152
rect 11664 10115 11722 10121
rect 11664 10081 11676 10115
rect 11710 10112 11722 10115
rect 11790 10112 11796 10124
rect 11710 10084 11796 10112
rect 11710 10081 11722 10084
rect 11664 10075 11722 10081
rect 11790 10072 11796 10084
rect 11848 10112 11854 10124
rect 12526 10112 12532 10124
rect 11848 10084 12532 10112
rect 11848 10072 11854 10084
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 12802 10112 12808 10124
rect 12636 10084 12808 10112
rect 11882 10044 11888 10056
rect 11843 10016 11888 10044
rect 11882 10004 11888 10016
rect 11940 10044 11946 10056
rect 12636 10044 12664 10084
rect 12802 10072 12808 10084
rect 12860 10072 12866 10124
rect 13096 10121 13124 10152
rect 13262 10140 13268 10192
rect 13320 10180 13326 10192
rect 16022 10180 16028 10192
rect 13320 10152 16028 10180
rect 13320 10140 13326 10152
rect 16022 10140 16028 10152
rect 16080 10180 16086 10192
rect 16482 10180 16488 10192
rect 16080 10152 16488 10180
rect 16080 10140 16086 10152
rect 16482 10140 16488 10152
rect 16540 10140 16546 10192
rect 17034 10140 17040 10192
rect 17092 10180 17098 10192
rect 23492 10189 23520 10220
rect 17773 10183 17831 10189
rect 17773 10180 17785 10183
rect 17092 10152 17785 10180
rect 17092 10140 17098 10152
rect 17773 10149 17785 10152
rect 17819 10149 17831 10183
rect 17773 10143 17831 10149
rect 23477 10183 23535 10189
rect 23477 10149 23489 10183
rect 23523 10149 23535 10183
rect 24026 10180 24032 10192
rect 23987 10152 24032 10180
rect 23477 10143 23535 10149
rect 24026 10140 24032 10152
rect 24084 10140 24090 10192
rect 24946 10140 24952 10192
rect 25004 10180 25010 10192
rect 25041 10183 25099 10189
rect 25041 10180 25053 10183
rect 25004 10152 25053 10180
rect 25004 10140 25010 10152
rect 25041 10149 25053 10152
rect 25087 10149 25099 10183
rect 25041 10143 25099 10149
rect 13081 10115 13139 10121
rect 13081 10081 13093 10115
rect 13127 10112 13139 10115
rect 13446 10112 13452 10124
rect 13127 10084 13452 10112
rect 13127 10081 13139 10084
rect 13081 10075 13139 10081
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 13541 10115 13599 10121
rect 13541 10081 13553 10115
rect 13587 10112 13599 10115
rect 13814 10112 13820 10124
rect 13587 10084 13820 10112
rect 13587 10081 13599 10084
rect 13541 10075 13599 10081
rect 13556 10044 13584 10075
rect 13814 10072 13820 10084
rect 13872 10072 13878 10124
rect 16393 10115 16451 10121
rect 16393 10081 16405 10115
rect 16439 10112 16451 10115
rect 16574 10112 16580 10124
rect 16439 10084 16580 10112
rect 16439 10081 16451 10084
rect 16393 10075 16451 10081
rect 16574 10072 16580 10084
rect 16632 10112 16638 10124
rect 18690 10112 18696 10124
rect 16632 10084 18696 10112
rect 16632 10072 16638 10084
rect 18690 10072 18696 10084
rect 18748 10072 18754 10124
rect 19334 10112 19340 10124
rect 19295 10084 19340 10112
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 14826 10044 14832 10056
rect 11940 10016 12664 10044
rect 12728 10016 13584 10044
rect 13786 10016 14832 10044
rect 11940 10004 11946 10016
rect 12728 9920 12756 10016
rect 12802 9936 12808 9988
rect 12860 9976 12866 9988
rect 13786 9976 13814 10016
rect 14826 10004 14832 10016
rect 14884 10044 14890 10056
rect 15562 10044 15568 10056
rect 14884 10016 15568 10044
rect 14884 10004 14890 10016
rect 15562 10004 15568 10016
rect 15620 10044 15626 10056
rect 16666 10044 16672 10056
rect 15620 10016 16672 10044
rect 15620 10004 15626 10016
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 17678 10004 17684 10056
rect 17736 10044 17742 10056
rect 18141 10047 18199 10053
rect 18141 10044 18153 10047
rect 17736 10016 18153 10044
rect 17736 10004 17742 10016
rect 18141 10013 18153 10016
rect 18187 10013 18199 10047
rect 18141 10007 18199 10013
rect 18509 10047 18567 10053
rect 18509 10013 18521 10047
rect 18555 10044 18567 10047
rect 19797 10047 19855 10053
rect 19797 10044 19809 10047
rect 18555 10016 19809 10044
rect 18555 10013 18567 10016
rect 18509 10007 18567 10013
rect 19797 10013 19809 10016
rect 19843 10044 19855 10047
rect 19886 10044 19892 10056
rect 19843 10016 19892 10044
rect 19843 10013 19855 10016
rect 19797 10007 19855 10013
rect 19886 10004 19892 10016
rect 19944 10004 19950 10056
rect 20901 10047 20959 10053
rect 20901 10013 20913 10047
rect 20947 10044 20959 10047
rect 21174 10044 21180 10056
rect 20947 10016 21180 10044
rect 20947 10013 20959 10016
rect 20901 10007 20959 10013
rect 21174 10004 21180 10016
rect 21232 10004 21238 10056
rect 23382 10044 23388 10056
rect 23343 10016 23388 10044
rect 23382 10004 23388 10016
rect 23440 10004 23446 10056
rect 24949 10047 25007 10053
rect 24949 10013 24961 10047
rect 24995 10044 25007 10047
rect 25222 10044 25228 10056
rect 24995 10016 25228 10044
rect 24995 10013 25007 10016
rect 24949 10007 25007 10013
rect 25222 10004 25228 10016
rect 25280 10044 25286 10056
rect 26050 10044 26056 10056
rect 25280 10016 26056 10044
rect 25280 10004 25286 10016
rect 26050 10004 26056 10016
rect 26108 10004 26114 10056
rect 16298 9976 16304 9988
rect 12860 9948 13814 9976
rect 14292 9948 16304 9976
rect 12860 9936 12866 9948
rect 14292 9920 14320 9948
rect 16298 9936 16304 9948
rect 16356 9976 16362 9988
rect 16761 9979 16819 9985
rect 16761 9976 16773 9979
rect 16356 9948 16773 9976
rect 16356 9936 16362 9948
rect 16761 9945 16773 9948
rect 16807 9976 16819 9979
rect 17589 9979 17647 9985
rect 17589 9976 17601 9979
rect 16807 9948 17601 9976
rect 16807 9945 16819 9948
rect 16761 9939 16819 9945
rect 17589 9945 17601 9948
rect 17635 9976 17647 9979
rect 17862 9976 17868 9988
rect 17635 9948 17868 9976
rect 17635 9945 17647 9948
rect 17589 9939 17647 9945
rect 17862 9936 17868 9948
rect 17920 9985 17926 9988
rect 17920 9979 17969 9985
rect 17920 9945 17923 9979
rect 17957 9976 17969 9979
rect 18785 9979 18843 9985
rect 18785 9976 18797 9979
rect 17957 9948 18797 9976
rect 17957 9945 17969 9948
rect 17920 9939 17969 9945
rect 18785 9945 18797 9948
rect 18831 9945 18843 9979
rect 25498 9976 25504 9988
rect 25459 9948 25504 9976
rect 18785 9939 18843 9945
rect 17920 9936 17926 9939
rect 25498 9936 25504 9948
rect 25556 9936 25562 9988
rect 10870 9908 10876 9920
rect 10831 9880 10876 9908
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 11698 9868 11704 9920
rect 11756 9908 11762 9920
rect 11793 9911 11851 9917
rect 11793 9908 11805 9911
rect 11756 9880 11805 9908
rect 11756 9868 11762 9880
rect 11793 9877 11805 9880
rect 11839 9877 11851 9911
rect 11793 9871 11851 9877
rect 12161 9911 12219 9917
rect 12161 9877 12173 9911
rect 12207 9908 12219 9911
rect 12710 9908 12716 9920
rect 12207 9880 12716 9908
rect 12207 9877 12219 9880
rect 12161 9871 12219 9877
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 14185 9911 14243 9917
rect 14185 9877 14197 9911
rect 14231 9908 14243 9911
rect 14274 9908 14280 9920
rect 14231 9880 14280 9908
rect 14231 9877 14243 9880
rect 14185 9871 14243 9877
rect 14274 9868 14280 9880
rect 14332 9868 14338 9920
rect 14550 9868 14556 9920
rect 14608 9908 14614 9920
rect 15013 9911 15071 9917
rect 15013 9908 15025 9911
rect 14608 9880 15025 9908
rect 14608 9868 14614 9880
rect 15013 9877 15025 9880
rect 15059 9908 15071 9911
rect 15286 9908 15292 9920
rect 15059 9880 15292 9908
rect 15059 9877 15071 9880
rect 15013 9871 15071 9877
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 16209 9911 16267 9917
rect 16209 9877 16221 9911
rect 16255 9908 16267 9911
rect 16390 9908 16396 9920
rect 16255 9880 16396 9908
rect 16255 9877 16267 9880
rect 16209 9871 16267 9877
rect 16390 9868 16396 9880
rect 16448 9868 16454 9920
rect 17402 9868 17408 9920
rect 17460 9908 17466 9920
rect 18049 9911 18107 9917
rect 18049 9908 18061 9911
rect 17460 9880 18061 9908
rect 17460 9868 17466 9880
rect 18049 9877 18061 9880
rect 18095 9908 18107 9911
rect 18322 9908 18328 9920
rect 18095 9880 18328 9908
rect 18095 9877 18107 9880
rect 18049 9871 18107 9877
rect 18322 9868 18328 9880
rect 18380 9868 18386 9920
rect 18414 9868 18420 9920
rect 18472 9908 18478 9920
rect 19521 9911 19579 9917
rect 19521 9908 19533 9911
rect 18472 9880 19533 9908
rect 18472 9868 18478 9880
rect 19521 9877 19533 9880
rect 19567 9877 19579 9911
rect 19521 9871 19579 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 11790 9704 11796 9716
rect 11751 9676 11796 9704
rect 11790 9664 11796 9676
rect 11848 9664 11854 9716
rect 12710 9704 12716 9716
rect 12671 9676 12716 9704
rect 12710 9664 12716 9676
rect 12768 9664 12774 9716
rect 13081 9707 13139 9713
rect 13081 9673 13093 9707
rect 13127 9704 13139 9707
rect 13446 9704 13452 9716
rect 13127 9676 13452 9704
rect 13127 9673 13139 9676
rect 13081 9667 13139 9673
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 14074 9707 14132 9713
rect 14074 9673 14086 9707
rect 14120 9704 14132 9707
rect 14274 9704 14280 9716
rect 14120 9676 14280 9704
rect 14120 9673 14132 9676
rect 14074 9667 14132 9673
rect 14274 9664 14280 9676
rect 14332 9664 14338 9716
rect 16574 9704 16580 9716
rect 16535 9676 16580 9704
rect 16574 9664 16580 9676
rect 16632 9664 16638 9716
rect 17034 9704 17040 9716
rect 16995 9676 17040 9704
rect 17034 9664 17040 9676
rect 17092 9704 17098 9716
rect 18322 9704 18328 9716
rect 17092 9676 18328 9704
rect 17092 9664 17098 9676
rect 18322 9664 18328 9676
rect 18380 9664 18386 9716
rect 21174 9664 21180 9716
rect 21232 9704 21238 9716
rect 22189 9707 22247 9713
rect 22189 9704 22201 9707
rect 21232 9676 22201 9704
rect 21232 9664 21238 9676
rect 22189 9673 22201 9676
rect 22235 9673 22247 9707
rect 22189 9667 22247 9673
rect 23109 9707 23167 9713
rect 23109 9673 23121 9707
rect 23155 9704 23167 9707
rect 23290 9704 23296 9716
rect 23155 9676 23296 9704
rect 23155 9673 23167 9676
rect 23109 9667 23167 9673
rect 23290 9664 23296 9676
rect 23348 9664 23354 9716
rect 23385 9707 23443 9713
rect 23385 9673 23397 9707
rect 23431 9673 23443 9707
rect 24946 9704 24952 9716
rect 24907 9676 24952 9704
rect 23385 9667 23443 9673
rect 9953 9639 10011 9645
rect 9953 9605 9965 9639
rect 9999 9636 10011 9639
rect 12986 9636 12992 9648
rect 9999 9608 12992 9636
rect 9999 9605 10011 9608
rect 9953 9599 10011 9605
rect 12986 9596 12992 9608
rect 13044 9596 13050 9648
rect 14185 9639 14243 9645
rect 14185 9636 14197 9639
rect 13740 9608 14197 9636
rect 8754 9528 8760 9580
rect 8812 9568 8818 9580
rect 13740 9577 13768 9608
rect 14185 9605 14197 9608
rect 14231 9636 14243 9639
rect 15746 9636 15752 9648
rect 14231 9608 15752 9636
rect 14231 9605 14243 9608
rect 14185 9599 14243 9605
rect 15746 9596 15752 9608
rect 15804 9636 15810 9648
rect 16206 9636 16212 9648
rect 15804 9608 16212 9636
rect 15804 9596 15810 9608
rect 16206 9596 16212 9608
rect 16264 9636 16270 9648
rect 17402 9636 17408 9648
rect 16264 9608 17408 9636
rect 16264 9596 16270 9608
rect 17402 9596 17408 9608
rect 17460 9596 17466 9648
rect 22646 9596 22652 9648
rect 22704 9636 22710 9648
rect 23400 9636 23428 9667
rect 24946 9664 24952 9676
rect 25004 9664 25010 9716
rect 25774 9704 25780 9716
rect 25735 9676 25780 9704
rect 25774 9664 25780 9676
rect 25832 9664 25838 9716
rect 26050 9704 26056 9716
rect 26011 9676 26056 9704
rect 26050 9664 26056 9676
rect 26108 9664 26114 9716
rect 23842 9636 23848 9648
rect 22704 9608 23848 9636
rect 22704 9596 22710 9608
rect 23842 9596 23848 9608
rect 23900 9596 23906 9648
rect 13725 9571 13783 9577
rect 13725 9568 13737 9571
rect 8812 9540 13737 9568
rect 8812 9528 8818 9540
rect 13725 9537 13737 9540
rect 13771 9537 13783 9571
rect 14366 9568 14372 9580
rect 14327 9540 14372 9568
rect 13725 9531 13783 9537
rect 14366 9528 14372 9540
rect 14424 9528 14430 9580
rect 14642 9528 14648 9580
rect 14700 9568 14706 9580
rect 18877 9571 18935 9577
rect 18877 9568 18889 9571
rect 14700 9540 18889 9568
rect 14700 9528 14706 9540
rect 18877 9537 18889 9540
rect 18923 9568 18935 9571
rect 19150 9568 19156 9580
rect 18923 9540 19156 9568
rect 18923 9537 18935 9540
rect 18877 9531 18935 9537
rect 19150 9528 19156 9540
rect 19208 9568 19214 9580
rect 22741 9571 22799 9577
rect 19208 9540 19472 9568
rect 19208 9528 19214 9540
rect 9769 9503 9827 9509
rect 9769 9469 9781 9503
rect 9815 9469 9827 9503
rect 10870 9500 10876 9512
rect 10831 9472 10876 9500
rect 9769 9463 9827 9469
rect 9784 9432 9812 9463
rect 10870 9460 10876 9472
rect 10928 9500 10934 9512
rect 12710 9500 12716 9512
rect 10928 9472 12716 9500
rect 10928 9460 10934 9472
rect 12710 9460 12716 9472
rect 12768 9460 12774 9512
rect 12894 9500 12900 9512
rect 12855 9472 12900 9500
rect 12894 9460 12900 9472
rect 12952 9500 12958 9512
rect 13357 9503 13415 9509
rect 13357 9500 13369 9503
rect 12952 9472 13369 9500
rect 12952 9460 12958 9472
rect 13357 9469 13369 9472
rect 13403 9469 13415 9503
rect 13357 9463 13415 9469
rect 14248 9503 14306 9509
rect 14248 9469 14260 9503
rect 14294 9500 14306 9503
rect 14826 9500 14832 9512
rect 14294 9472 14832 9500
rect 14294 9469 14306 9472
rect 14248 9463 14306 9469
rect 10321 9435 10379 9441
rect 10321 9432 10333 9435
rect 9784 9404 10333 9432
rect 10321 9401 10333 9404
rect 10367 9432 10379 9435
rect 10686 9432 10692 9444
rect 10367 9404 10692 9432
rect 10367 9401 10379 9404
rect 10321 9395 10379 9401
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 11514 9432 11520 9444
rect 11475 9404 11520 9432
rect 11514 9392 11520 9404
rect 11572 9392 11578 9444
rect 11974 9392 11980 9444
rect 12032 9432 12038 9444
rect 13262 9432 13268 9444
rect 12032 9404 13268 9432
rect 12032 9392 12038 9404
rect 13262 9392 13268 9404
rect 13320 9392 13326 9444
rect 13372 9432 13400 9463
rect 14826 9460 14832 9472
rect 14884 9460 14890 9512
rect 15378 9500 15384 9512
rect 15291 9472 15384 9500
rect 15378 9460 15384 9472
rect 15436 9500 15442 9512
rect 15565 9503 15623 9509
rect 15565 9500 15577 9503
rect 15436 9472 15577 9500
rect 15436 9460 15442 9472
rect 15565 9469 15577 9472
rect 15611 9469 15623 9503
rect 15565 9463 15623 9469
rect 15838 9460 15844 9512
rect 15896 9500 15902 9512
rect 17678 9500 17684 9512
rect 15896 9472 17684 9500
rect 15896 9460 15902 9472
rect 17678 9460 17684 9472
rect 17736 9500 17742 9512
rect 17773 9503 17831 9509
rect 17773 9500 17785 9503
rect 17736 9472 17785 9500
rect 17736 9460 17742 9472
rect 17773 9469 17785 9472
rect 17819 9469 17831 9503
rect 18046 9500 18052 9512
rect 18007 9472 18052 9500
rect 17773 9463 17831 9469
rect 18046 9460 18052 9472
rect 18104 9500 18110 9512
rect 18509 9503 18567 9509
rect 18509 9500 18521 9503
rect 18104 9472 18521 9500
rect 18104 9460 18110 9472
rect 18509 9469 18521 9472
rect 18555 9500 18567 9503
rect 19245 9503 19303 9509
rect 19245 9500 19257 9503
rect 18555 9472 19257 9500
rect 18555 9469 18567 9472
rect 18509 9463 18567 9469
rect 19245 9469 19257 9472
rect 19291 9500 19303 9503
rect 19334 9500 19340 9512
rect 19291 9472 19340 9500
rect 19291 9469 19303 9472
rect 19245 9463 19303 9469
rect 19334 9460 19340 9472
rect 19392 9460 19398 9512
rect 19444 9509 19472 9540
rect 22741 9537 22753 9571
rect 22787 9568 22799 9571
rect 23382 9568 23388 9580
rect 22787 9540 23388 9568
rect 22787 9537 22799 9540
rect 22741 9531 22799 9537
rect 23382 9528 23388 9540
rect 23440 9568 23446 9580
rect 24029 9571 24087 9577
rect 24029 9568 24041 9571
rect 23440 9540 24041 9568
rect 23440 9528 23446 9540
rect 24029 9537 24041 9540
rect 24075 9537 24087 9571
rect 24029 9531 24087 9537
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9469 19487 9503
rect 19886 9500 19892 9512
rect 19847 9472 19892 9500
rect 19429 9463 19487 9469
rect 19886 9460 19892 9472
rect 19944 9460 19950 9512
rect 20165 9503 20223 9509
rect 20165 9469 20177 9503
rect 20211 9500 20223 9503
rect 20993 9503 21051 9509
rect 20993 9500 21005 9503
rect 20211 9472 21005 9500
rect 20211 9469 20223 9472
rect 20165 9463 20223 9469
rect 20993 9469 21005 9472
rect 21039 9500 21051 9503
rect 21082 9500 21088 9512
rect 21039 9472 21088 9500
rect 21039 9469 21051 9472
rect 20993 9463 21051 9469
rect 21082 9460 21088 9472
rect 21140 9460 21146 9512
rect 22554 9460 22560 9512
rect 22612 9500 22618 9512
rect 23290 9500 23296 9512
rect 22612 9472 23296 9500
rect 22612 9460 22618 9472
rect 23290 9460 23296 9472
rect 23348 9460 23354 9512
rect 25276 9503 25334 9509
rect 25276 9469 25288 9503
rect 25322 9500 25334 9503
rect 25774 9500 25780 9512
rect 25322 9472 25780 9500
rect 25322 9469 25334 9472
rect 25276 9463 25334 9469
rect 25774 9460 25780 9472
rect 25832 9460 25838 9512
rect 13906 9432 13912 9444
rect 13372 9404 13814 9432
rect 13867 9404 13912 9432
rect 10042 9324 10048 9376
rect 10100 9364 10106 9376
rect 10597 9367 10655 9373
rect 10597 9364 10609 9367
rect 10100 9336 10609 9364
rect 10100 9324 10106 9336
rect 10597 9333 10609 9336
rect 10643 9364 10655 9367
rect 11882 9364 11888 9376
rect 10643 9336 11888 9364
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 12066 9324 12072 9376
rect 12124 9364 12130 9376
rect 12161 9367 12219 9373
rect 12161 9364 12173 9367
rect 12124 9336 12173 9364
rect 12124 9324 12130 9336
rect 12161 9333 12173 9336
rect 12207 9333 12219 9367
rect 13786 9364 13814 9404
rect 13906 9392 13912 9404
rect 13964 9392 13970 9444
rect 15286 9432 15292 9444
rect 14384 9404 15292 9432
rect 14384 9364 14412 9404
rect 15286 9392 15292 9404
rect 15344 9392 15350 9444
rect 16209 9435 16267 9441
rect 16209 9401 16221 9435
rect 16255 9432 16267 9435
rect 16298 9432 16304 9444
rect 16255 9404 16304 9432
rect 16255 9401 16267 9404
rect 16209 9395 16267 9401
rect 16298 9392 16304 9404
rect 16356 9392 16362 9444
rect 21314 9435 21372 9441
rect 21314 9432 21326 9435
rect 21192 9404 21326 9432
rect 21192 9376 21220 9404
rect 21314 9401 21326 9404
rect 21360 9401 21372 9435
rect 23750 9432 23756 9444
rect 23711 9404 23756 9432
rect 21314 9395 21372 9401
rect 23750 9392 23756 9404
rect 23808 9392 23814 9444
rect 23842 9392 23848 9444
rect 23900 9432 23906 9444
rect 25363 9435 25421 9441
rect 25363 9432 25375 9435
rect 23900 9404 23945 9432
rect 24504 9404 25375 9432
rect 23900 9392 23906 9404
rect 13786 9336 14412 9364
rect 12161 9327 12219 9333
rect 14826 9324 14832 9376
rect 14884 9364 14890 9376
rect 14921 9367 14979 9373
rect 14921 9364 14933 9367
rect 14884 9336 14933 9364
rect 14884 9324 14890 9336
rect 14921 9333 14933 9336
rect 14967 9333 14979 9367
rect 14921 9327 14979 9333
rect 18233 9367 18291 9373
rect 18233 9333 18245 9367
rect 18279 9364 18291 9367
rect 19242 9364 19248 9376
rect 18279 9336 19248 9364
rect 18279 9333 18291 9336
rect 18233 9327 18291 9333
rect 19242 9324 19248 9336
rect 19300 9324 19306 9376
rect 20533 9367 20591 9373
rect 20533 9333 20545 9367
rect 20579 9364 20591 9367
rect 20809 9367 20867 9373
rect 20809 9364 20821 9367
rect 20579 9336 20821 9364
rect 20579 9333 20591 9336
rect 20533 9327 20591 9333
rect 20809 9333 20821 9336
rect 20855 9364 20867 9367
rect 21174 9364 21180 9376
rect 20855 9336 21180 9364
rect 20855 9333 20867 9336
rect 20809 9327 20867 9333
rect 21174 9324 21180 9336
rect 21232 9324 21238 9376
rect 21913 9367 21971 9373
rect 21913 9333 21925 9367
rect 21959 9364 21971 9367
rect 22922 9364 22928 9376
rect 21959 9336 22928 9364
rect 21959 9333 21971 9336
rect 21913 9327 21971 9333
rect 22922 9324 22928 9336
rect 22980 9324 22986 9376
rect 23106 9324 23112 9376
rect 23164 9364 23170 9376
rect 24504 9364 24532 9404
rect 25363 9401 25375 9404
rect 25409 9401 25421 9435
rect 25363 9395 25421 9401
rect 23164 9336 24532 9364
rect 23164 9324 23170 9336
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 10686 9120 10692 9172
rect 10744 9160 10750 9172
rect 18046 9160 18052 9172
rect 10744 9132 18052 9160
rect 10744 9120 10750 9132
rect 11514 9052 11520 9104
rect 11572 9092 11578 9104
rect 13541 9095 13599 9101
rect 13541 9092 13553 9095
rect 11572 9064 13553 9092
rect 11572 9052 11578 9064
rect 13541 9061 13553 9064
rect 13587 9092 13599 9095
rect 13722 9092 13728 9104
rect 13587 9064 13728 9092
rect 13587 9061 13599 9064
rect 13541 9055 13599 9061
rect 13722 9052 13728 9064
rect 13780 9052 13786 9104
rect 13906 9052 13912 9104
rect 13964 9092 13970 9104
rect 14461 9095 14519 9101
rect 14461 9092 14473 9095
rect 13964 9064 14473 9092
rect 13964 9052 13970 9064
rect 14461 9061 14473 9064
rect 14507 9092 14519 9095
rect 14734 9092 14740 9104
rect 14507 9064 14740 9092
rect 14507 9061 14519 9064
rect 14461 9055 14519 9061
rect 14734 9052 14740 9064
rect 14792 9052 14798 9104
rect 15304 9101 15332 9132
rect 18046 9120 18052 9132
rect 18104 9120 18110 9172
rect 21082 9160 21088 9172
rect 21043 9132 21088 9160
rect 21082 9120 21088 9132
rect 21140 9120 21146 9172
rect 22186 9160 22192 9172
rect 22147 9132 22192 9160
rect 22186 9120 22192 9132
rect 22244 9120 22250 9172
rect 22922 9120 22928 9172
rect 22980 9160 22986 9172
rect 22980 9132 24808 9160
rect 22980 9120 22986 9132
rect 15289 9095 15347 9101
rect 15289 9061 15301 9095
rect 15335 9061 15347 9095
rect 17862 9092 17868 9104
rect 15289 9055 15347 9061
rect 17144 9064 17724 9092
rect 17823 9064 17868 9092
rect 10873 9027 10931 9033
rect 10873 8993 10885 9027
rect 10919 8993 10931 9027
rect 11974 9024 11980 9036
rect 11935 8996 11980 9024
rect 10873 8987 10931 8993
rect 9674 8848 9680 8900
rect 9732 8888 9738 8900
rect 10888 8888 10916 8987
rect 11974 8984 11980 8996
rect 12032 8984 12038 9036
rect 12342 8984 12348 9036
rect 12400 9024 12406 9036
rect 15381 9027 15439 9033
rect 12400 8996 12445 9024
rect 12400 8984 12406 8996
rect 15381 8993 15393 9027
rect 15427 8993 15439 9027
rect 15381 8987 15439 8993
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8956 11023 8959
rect 12158 8956 12164 8968
rect 11011 8928 12164 8956
rect 11011 8925 11023 8928
rect 10965 8919 11023 8925
rect 12158 8916 12164 8928
rect 12216 8916 12222 8968
rect 12526 8956 12532 8968
rect 12487 8928 12532 8956
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 13446 8956 13452 8968
rect 13407 8928 13452 8956
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 15286 8916 15292 8968
rect 15344 8956 15350 8968
rect 15396 8956 15424 8987
rect 16482 8984 16488 9036
rect 16540 9024 16546 9036
rect 16942 9024 16948 9036
rect 16540 8996 16948 9024
rect 16540 8984 16546 8996
rect 16942 8984 16948 8996
rect 17000 9024 17006 9036
rect 17144 9033 17172 9064
rect 17129 9027 17187 9033
rect 17129 9024 17141 9027
rect 17000 8996 17141 9024
rect 17000 8984 17006 8996
rect 17129 8993 17141 8996
rect 17175 8993 17187 9027
rect 17310 9024 17316 9036
rect 17271 8996 17316 9024
rect 17129 8987 17187 8993
rect 17310 8984 17316 8996
rect 17368 8984 17374 9036
rect 17696 9024 17724 9064
rect 17862 9052 17868 9064
rect 17920 9052 17926 9104
rect 19978 9092 19984 9104
rect 19812 9064 19984 9092
rect 18414 9024 18420 9036
rect 17696 8996 18420 9024
rect 18414 8984 18420 8996
rect 18472 8984 18478 9036
rect 18966 8984 18972 9036
rect 19024 9024 19030 9036
rect 19812 9033 19840 9064
rect 19978 9052 19984 9064
rect 20036 9052 20042 9104
rect 21174 9052 21180 9104
rect 21232 9092 21238 9104
rect 21590 9095 21648 9101
rect 21590 9092 21602 9095
rect 21232 9064 21602 9092
rect 21232 9052 21238 9064
rect 21590 9061 21602 9064
rect 21636 9061 21648 9095
rect 21590 9055 21648 9061
rect 21726 9052 21732 9104
rect 21784 9092 21790 9104
rect 23198 9092 23204 9104
rect 21784 9064 23204 9092
rect 21784 9052 21790 9064
rect 23198 9052 23204 9064
rect 23256 9052 23262 9104
rect 24780 9101 24808 9132
rect 24765 9095 24823 9101
rect 24765 9061 24777 9095
rect 24811 9092 24823 9095
rect 24854 9092 24860 9104
rect 24811 9064 24860 9092
rect 24811 9061 24823 9064
rect 24765 9055 24823 9061
rect 24854 9052 24860 9064
rect 24912 9052 24918 9104
rect 25317 9095 25375 9101
rect 25317 9061 25329 9095
rect 25363 9092 25375 9095
rect 25498 9092 25504 9104
rect 25363 9064 25504 9092
rect 25363 9061 25375 9064
rect 25317 9055 25375 9061
rect 25498 9052 25504 9064
rect 25556 9052 25562 9104
rect 19245 9027 19303 9033
rect 19245 9024 19257 9027
rect 19024 8996 19257 9024
rect 19024 8984 19030 8996
rect 19245 8993 19257 8996
rect 19291 8993 19303 9027
rect 19245 8987 19303 8993
rect 19797 9027 19855 9033
rect 19797 8993 19809 9027
rect 19843 8993 19855 9027
rect 19797 8987 19855 8993
rect 17586 8956 17592 8968
rect 15344 8928 15424 8956
rect 17547 8928 17592 8956
rect 15344 8916 15350 8928
rect 17586 8916 17592 8928
rect 17644 8916 17650 8968
rect 19981 8959 20039 8965
rect 19981 8925 19993 8959
rect 20027 8956 20039 8959
rect 21266 8956 21272 8968
rect 20027 8928 21272 8956
rect 20027 8925 20039 8928
rect 19981 8919 20039 8925
rect 21266 8916 21272 8928
rect 21324 8916 21330 8968
rect 23106 8956 23112 8968
rect 23067 8928 23112 8956
rect 23106 8916 23112 8928
rect 23164 8916 23170 8968
rect 23382 8956 23388 8968
rect 23343 8928 23388 8956
rect 23382 8916 23388 8928
rect 23440 8916 23446 8968
rect 24673 8959 24731 8965
rect 24673 8925 24685 8959
rect 24719 8956 24731 8959
rect 24762 8956 24768 8968
rect 24719 8928 24768 8956
rect 24719 8925 24731 8928
rect 24673 8919 24731 8925
rect 24762 8916 24768 8928
rect 24820 8916 24826 8968
rect 13170 8888 13176 8900
rect 9732 8860 13176 8888
rect 9732 8848 9738 8860
rect 13170 8848 13176 8860
rect 13228 8848 13234 8900
rect 13998 8888 14004 8900
rect 13959 8860 14004 8888
rect 13998 8848 14004 8860
rect 14056 8848 14062 8900
rect 8938 8780 8944 8832
rect 8996 8820 9002 8832
rect 11517 8823 11575 8829
rect 11517 8820 11529 8823
rect 8996 8792 11529 8820
rect 8996 8780 9002 8792
rect 11517 8789 11529 8792
rect 11563 8820 11575 8823
rect 11698 8820 11704 8832
rect 11563 8792 11704 8820
rect 11563 8789 11575 8792
rect 11517 8783 11575 8789
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 13081 8823 13139 8829
rect 13081 8820 13093 8823
rect 11848 8792 13093 8820
rect 11848 8780 11854 8792
rect 13081 8789 13093 8792
rect 13127 8820 13139 8823
rect 13354 8820 13360 8832
rect 13127 8792 13360 8820
rect 13127 8789 13139 8792
rect 13081 8783 13139 8789
rect 13354 8780 13360 8792
rect 13412 8780 13418 8832
rect 15470 8780 15476 8832
rect 15528 8820 15534 8832
rect 16301 8823 16359 8829
rect 16301 8820 16313 8823
rect 15528 8792 16313 8820
rect 15528 8780 15534 8792
rect 16301 8789 16313 8792
rect 16347 8789 16359 8823
rect 18874 8820 18880 8832
rect 18835 8792 18880 8820
rect 16301 8783 16359 8789
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 22554 8820 22560 8832
rect 22515 8792 22560 8820
rect 22554 8780 22560 8792
rect 22612 8780 22618 8832
rect 23750 8780 23756 8832
rect 23808 8820 23814 8832
rect 24026 8820 24032 8832
rect 23808 8792 24032 8820
rect 23808 8780 23814 8792
rect 24026 8780 24032 8792
rect 24084 8780 24090 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 9306 8616 9312 8628
rect 9267 8588 9312 8616
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 9674 8616 9680 8628
rect 9635 8588 9680 8616
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 9950 8616 9956 8628
rect 9911 8588 9956 8616
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 11974 8616 11980 8628
rect 11931 8588 11980 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 11974 8576 11980 8588
rect 12032 8576 12038 8628
rect 12250 8616 12256 8628
rect 12211 8588 12256 8616
rect 12250 8576 12256 8588
rect 12308 8576 12314 8628
rect 13446 8576 13452 8628
rect 13504 8616 13510 8628
rect 14093 8619 14151 8625
rect 14093 8616 14105 8619
rect 13504 8588 14105 8616
rect 13504 8576 13510 8588
rect 14093 8585 14105 8588
rect 14139 8616 14151 8619
rect 14139 8588 14320 8616
rect 14139 8585 14151 8588
rect 14093 8579 14151 8585
rect 8895 8551 8953 8557
rect 8895 8517 8907 8551
rect 8941 8548 8953 8551
rect 13538 8548 13544 8560
rect 8941 8520 13544 8548
rect 8941 8517 8953 8520
rect 8895 8511 8953 8517
rect 13538 8508 13544 8520
rect 13596 8508 13602 8560
rect 13722 8548 13728 8560
rect 13683 8520 13728 8548
rect 13722 8508 13728 8520
rect 13780 8508 13786 8560
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8480 10747 8483
rect 11790 8480 11796 8492
rect 10735 8452 11796 8480
rect 10735 8449 10747 8452
rect 10689 8443 10747 8449
rect 8824 8415 8882 8421
rect 8824 8381 8836 8415
rect 8870 8412 8882 8415
rect 9306 8412 9312 8424
rect 8870 8384 9312 8412
rect 8870 8381 8882 8384
rect 8824 8375 8882 8381
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 11072 8421 11100 8452
rect 11790 8440 11796 8452
rect 11848 8440 11854 8492
rect 12526 8480 12532 8492
rect 12487 8452 12532 8480
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 14292 8489 14320 8588
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 15933 8619 15991 8625
rect 15933 8616 15945 8619
rect 14516 8588 15945 8616
rect 14516 8576 14522 8588
rect 15933 8585 15945 8588
rect 15979 8585 15991 8619
rect 16942 8616 16948 8628
rect 16903 8588 16948 8616
rect 15933 8579 15991 8585
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 17310 8616 17316 8628
rect 17271 8588 17316 8616
rect 17310 8576 17316 8588
rect 17368 8576 17374 8628
rect 19889 8619 19947 8625
rect 19889 8585 19901 8619
rect 19935 8616 19947 8619
rect 19978 8616 19984 8628
rect 19935 8588 19984 8616
rect 19935 8585 19947 8588
rect 19889 8579 19947 8585
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 23109 8619 23167 8625
rect 23109 8585 23121 8619
rect 23155 8616 23167 8619
rect 23198 8616 23204 8628
rect 23155 8588 23204 8616
rect 23155 8585 23167 8588
rect 23109 8579 23167 8585
rect 23198 8576 23204 8588
rect 23256 8576 23262 8628
rect 23290 8576 23296 8628
rect 23348 8616 23354 8628
rect 23385 8619 23443 8625
rect 23385 8616 23397 8619
rect 23348 8588 23397 8616
rect 23348 8576 23354 8588
rect 23385 8585 23397 8588
rect 23431 8616 23443 8619
rect 23842 8616 23848 8628
rect 23431 8588 23848 8616
rect 23431 8585 23443 8588
rect 23385 8579 23443 8585
rect 23842 8576 23848 8588
rect 23900 8576 23906 8628
rect 24765 8619 24823 8625
rect 24765 8585 24777 8619
rect 24811 8616 24823 8619
rect 24854 8616 24860 8628
rect 24811 8588 24860 8616
rect 24811 8585 24823 8588
rect 24765 8579 24823 8585
rect 24854 8576 24860 8588
rect 24912 8576 24918 8628
rect 25774 8616 25780 8628
rect 25735 8588 25780 8616
rect 25774 8576 25780 8588
rect 25832 8576 25838 8628
rect 15746 8548 15752 8560
rect 15707 8520 15752 8548
rect 15746 8508 15752 8520
rect 15804 8548 15810 8560
rect 16485 8551 16543 8557
rect 16485 8548 16497 8551
rect 15804 8520 16497 8548
rect 15804 8508 15810 8520
rect 16485 8517 16497 8520
rect 16531 8517 16543 8551
rect 19426 8548 19432 8560
rect 19387 8520 19432 8548
rect 16485 8511 16543 8517
rect 19426 8508 19432 8520
rect 19484 8508 19490 8560
rect 21085 8551 21143 8557
rect 21085 8517 21097 8551
rect 21131 8548 21143 8551
rect 22649 8551 22707 8557
rect 22649 8548 22661 8551
rect 21131 8520 22661 8548
rect 21131 8517 21143 8520
rect 21085 8511 21143 8517
rect 22649 8517 22661 8520
rect 22695 8548 22707 8551
rect 23014 8548 23020 8560
rect 22695 8520 23020 8548
rect 22695 8517 22707 8520
rect 22649 8511 22707 8517
rect 23014 8508 23020 8520
rect 23072 8508 23078 8560
rect 14277 8483 14335 8489
rect 14277 8449 14289 8483
rect 14323 8449 14335 8483
rect 14277 8443 14335 8449
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 15620 8483 15678 8489
rect 15620 8480 15632 8483
rect 15528 8452 15632 8480
rect 15528 8440 15534 8452
rect 15620 8449 15632 8452
rect 15666 8449 15678 8483
rect 15838 8480 15844 8492
rect 15799 8452 15844 8480
rect 15620 8443 15678 8449
rect 15838 8440 15844 8452
rect 15896 8440 15902 8492
rect 18874 8480 18880 8492
rect 18787 8452 18880 8480
rect 18874 8440 18880 8452
rect 18932 8480 18938 8492
rect 20806 8480 20812 8492
rect 18932 8452 20812 8480
rect 18932 8440 18938 8452
rect 20806 8440 20812 8452
rect 20864 8440 20870 8492
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8480 22155 8483
rect 22554 8480 22560 8492
rect 22143 8452 22560 8480
rect 22143 8449 22155 8452
rect 22097 8443 22155 8449
rect 22554 8440 22560 8452
rect 22612 8480 22618 8492
rect 25130 8480 25136 8492
rect 22612 8452 25136 8480
rect 22612 8440 22618 8452
rect 25130 8440 25136 8452
rect 25188 8440 25194 8492
rect 9769 8415 9827 8421
rect 9769 8381 9781 8415
rect 9815 8381 9827 8415
rect 9769 8375 9827 8381
rect 11057 8415 11115 8421
rect 11057 8381 11069 8415
rect 11103 8381 11115 8415
rect 11330 8412 11336 8424
rect 11291 8384 11336 8412
rect 11057 8375 11115 8381
rect 9030 8304 9036 8356
rect 9088 8344 9094 8356
rect 9784 8344 9812 8375
rect 11330 8372 11336 8384
rect 11388 8372 11394 8424
rect 12158 8372 12164 8424
rect 12216 8412 12222 8424
rect 18601 8415 18659 8421
rect 18601 8412 18613 8415
rect 12216 8384 18613 8412
rect 12216 8372 12222 8384
rect 18601 8381 18613 8384
rect 18647 8381 18659 8415
rect 18601 8375 18659 8381
rect 25292 8415 25350 8421
rect 25292 8381 25304 8415
rect 25338 8412 25350 8415
rect 25774 8412 25780 8424
rect 25338 8384 25780 8412
rect 25338 8381 25350 8384
rect 25292 8375 25350 8381
rect 10321 8347 10379 8353
rect 10321 8344 10333 8347
rect 9088 8316 10333 8344
rect 9088 8304 9094 8316
rect 10321 8313 10333 8316
rect 10367 8344 10379 8347
rect 10686 8344 10692 8356
rect 10367 8316 10692 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 10686 8304 10692 8316
rect 10744 8304 10750 8356
rect 11514 8344 11520 8356
rect 11475 8316 11520 8344
rect 11514 8304 11520 8316
rect 11572 8304 11578 8356
rect 12250 8304 12256 8356
rect 12308 8344 12314 8356
rect 12850 8347 12908 8353
rect 12850 8344 12862 8347
rect 12308 8316 12862 8344
rect 12308 8304 12314 8316
rect 12850 8313 12862 8316
rect 12896 8313 12908 8347
rect 12850 8307 12908 8313
rect 15013 8347 15071 8353
rect 15013 8313 15025 8347
rect 15059 8344 15071 8347
rect 15473 8347 15531 8353
rect 15059 8316 15424 8344
rect 15059 8313 15071 8316
rect 15013 8307 15071 8313
rect 12710 8236 12716 8288
rect 12768 8276 12774 8288
rect 13446 8276 13452 8288
rect 12768 8248 13452 8276
rect 12768 8236 12774 8248
rect 13446 8236 13452 8248
rect 13504 8236 13510 8288
rect 15286 8276 15292 8288
rect 15247 8248 15292 8276
rect 15286 8236 15292 8248
rect 15344 8236 15350 8288
rect 15396 8276 15424 8316
rect 15473 8313 15485 8347
rect 15519 8344 15531 8347
rect 15562 8344 15568 8356
rect 15519 8316 15568 8344
rect 15519 8313 15531 8316
rect 15473 8307 15531 8313
rect 15562 8304 15568 8316
rect 15620 8304 15626 8356
rect 15838 8276 15844 8288
rect 15396 8248 15844 8276
rect 15838 8236 15844 8248
rect 15896 8236 15902 8288
rect 18616 8276 18644 8375
rect 25774 8372 25780 8384
rect 25832 8372 25838 8424
rect 18969 8347 19027 8353
rect 18969 8313 18981 8347
rect 19015 8313 19027 8347
rect 20530 8344 20536 8356
rect 20491 8316 20536 8344
rect 18969 8307 19027 8313
rect 18984 8276 19012 8307
rect 20530 8304 20536 8316
rect 20588 8304 20594 8356
rect 20622 8304 20628 8356
rect 20680 8344 20686 8356
rect 22189 8347 22247 8353
rect 20680 8316 20725 8344
rect 20680 8304 20686 8316
rect 22189 8313 22201 8347
rect 22235 8313 22247 8347
rect 22189 8307 22247 8313
rect 18616 8248 19012 8276
rect 20349 8279 20407 8285
rect 20349 8245 20361 8279
rect 20395 8276 20407 8279
rect 20640 8276 20668 8304
rect 20395 8248 20668 8276
rect 20395 8245 20407 8248
rect 20349 8239 20407 8245
rect 21174 8236 21180 8288
rect 21232 8276 21238 8288
rect 21453 8279 21511 8285
rect 21453 8276 21465 8279
rect 21232 8248 21465 8276
rect 21232 8236 21238 8248
rect 21453 8245 21465 8248
rect 21499 8245 21511 8279
rect 21818 8276 21824 8288
rect 21779 8248 21824 8276
rect 21453 8239 21511 8245
rect 21818 8236 21824 8248
rect 21876 8276 21882 8288
rect 22204 8276 22232 8307
rect 22278 8304 22284 8356
rect 22336 8344 22342 8356
rect 23750 8344 23756 8356
rect 22336 8316 23756 8344
rect 22336 8304 22342 8316
rect 23750 8304 23756 8316
rect 23808 8304 23814 8356
rect 23842 8304 23848 8356
rect 23900 8344 23906 8356
rect 24394 8344 24400 8356
rect 23900 8316 23945 8344
rect 24355 8316 24400 8344
rect 23900 8304 23906 8316
rect 24394 8304 24400 8316
rect 24452 8344 24458 8356
rect 24762 8344 24768 8356
rect 24452 8316 24768 8344
rect 24452 8304 24458 8316
rect 24762 8304 24768 8316
rect 24820 8344 24826 8356
rect 25041 8347 25099 8353
rect 25041 8344 25053 8347
rect 24820 8316 25053 8344
rect 24820 8304 24826 8316
rect 25041 8313 25053 8316
rect 25087 8313 25099 8347
rect 25041 8307 25099 8313
rect 21876 8248 22232 8276
rect 21876 8236 21882 8248
rect 23934 8236 23940 8288
rect 23992 8276 23998 8288
rect 25363 8279 25421 8285
rect 25363 8276 25375 8279
rect 23992 8248 25375 8276
rect 23992 8236 23998 8248
rect 25363 8245 25375 8248
rect 25409 8245 25421 8279
rect 25363 8239 25421 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 7699 8075 7757 8081
rect 7699 8041 7711 8075
rect 7745 8072 7757 8075
rect 7834 8072 7840 8084
rect 7745 8044 7840 8072
rect 7745 8041 7757 8044
rect 7699 8035 7757 8041
rect 7834 8032 7840 8044
rect 7892 8032 7898 8084
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 12066 8072 12072 8084
rect 8803 8044 12072 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 12250 8072 12256 8084
rect 12211 8044 12256 8072
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 13081 8075 13139 8081
rect 13081 8072 13093 8075
rect 12584 8044 13093 8072
rect 12584 8032 12590 8044
rect 13081 8041 13093 8044
rect 13127 8041 13139 8075
rect 13081 8035 13139 8041
rect 13170 8032 13176 8084
rect 13228 8072 13234 8084
rect 18601 8075 18659 8081
rect 18601 8072 18613 8075
rect 13228 8044 18613 8072
rect 13228 8032 13234 8044
rect 18601 8041 18613 8044
rect 18647 8072 18659 8075
rect 18690 8072 18696 8084
rect 18647 8044 18696 8072
rect 18647 8041 18659 8044
rect 18601 8035 18659 8041
rect 18690 8032 18696 8044
rect 18748 8032 18754 8084
rect 18782 8032 18788 8084
rect 18840 8072 18846 8084
rect 19705 8075 19763 8081
rect 19705 8072 19717 8075
rect 18840 8044 19717 8072
rect 18840 8032 18846 8044
rect 19705 8041 19717 8044
rect 19751 8041 19763 8075
rect 20530 8072 20536 8084
rect 20491 8044 20536 8072
rect 19705 8035 19763 8041
rect 20530 8032 20536 8044
rect 20588 8032 20594 8084
rect 21266 8072 21272 8084
rect 21227 8044 21272 8072
rect 21266 8032 21272 8044
rect 21324 8032 21330 8084
rect 23106 8072 23112 8084
rect 23067 8044 23112 8072
rect 23106 8032 23112 8044
rect 23164 8032 23170 8084
rect 23750 8072 23756 8084
rect 23711 8044 23756 8072
rect 23750 8032 23756 8044
rect 23808 8032 23814 8084
rect 25547 8075 25605 8081
rect 25547 8041 25559 8075
rect 25593 8041 25605 8075
rect 25547 8035 25605 8041
rect 13446 8004 13452 8016
rect 13407 7976 13452 8004
rect 13446 7964 13452 7976
rect 13504 8004 13510 8016
rect 13817 8007 13875 8013
rect 13817 8004 13829 8007
rect 13504 7976 13829 8004
rect 13504 7964 13510 7976
rect 13817 7973 13829 7976
rect 13863 7973 13875 8007
rect 13817 7967 13875 7973
rect 17862 7964 17868 8016
rect 17920 8004 17926 8016
rect 18002 8007 18060 8013
rect 18002 8004 18014 8007
rect 17920 7976 18014 8004
rect 17920 7964 17926 7976
rect 18002 7973 18014 7976
rect 18048 7973 18060 8007
rect 18002 7967 18060 7973
rect 18966 7964 18972 8016
rect 19024 8004 19030 8016
rect 19245 8007 19303 8013
rect 19245 8004 19257 8007
rect 19024 7976 19257 8004
rect 19024 7964 19030 7976
rect 19245 7973 19257 7976
rect 19291 7973 19303 8007
rect 19245 7967 19303 7973
rect 21174 7964 21180 8016
rect 21232 8004 21238 8016
rect 22142 8007 22200 8013
rect 22142 8004 22154 8007
rect 21232 7976 22154 8004
rect 21232 7964 21238 7976
rect 22142 7973 22154 7976
rect 22188 7973 22200 8007
rect 24026 8004 24032 8016
rect 23987 7976 24032 8004
rect 22142 7967 22200 7973
rect 24026 7964 24032 7976
rect 24084 7964 24090 8016
rect 25130 7964 25136 8016
rect 25188 8004 25194 8016
rect 25562 8004 25590 8035
rect 25188 7976 25590 8004
rect 25188 7964 25194 7976
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7936 7527 7939
rect 7650 7936 7656 7948
rect 7515 7908 7656 7936
rect 7515 7905 7527 7908
rect 7469 7899 7527 7905
rect 7650 7896 7656 7908
rect 7708 7896 7714 7948
rect 8573 7939 8631 7945
rect 8573 7905 8585 7939
rect 8619 7936 8631 7939
rect 8846 7936 8852 7948
rect 8619 7908 8852 7936
rect 8619 7905 8631 7908
rect 8573 7899 8631 7905
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 10410 7936 10416 7948
rect 10371 7908 10416 7936
rect 10410 7896 10416 7908
rect 10468 7896 10474 7948
rect 11514 7896 11520 7948
rect 11572 7936 11578 7948
rect 11885 7939 11943 7945
rect 11885 7936 11897 7939
rect 11572 7908 11897 7936
rect 11572 7896 11578 7908
rect 11885 7905 11897 7908
rect 11931 7905 11943 7939
rect 11885 7899 11943 7905
rect 15289 7939 15347 7945
rect 15289 7905 15301 7939
rect 15335 7936 15347 7939
rect 15562 7936 15568 7948
rect 15335 7908 15568 7936
rect 15335 7905 15347 7908
rect 15289 7899 15347 7905
rect 15562 7896 15568 7908
rect 15620 7936 15626 7948
rect 16206 7936 16212 7948
rect 15620 7908 16212 7936
rect 15620 7896 15626 7908
rect 16206 7896 16212 7908
rect 16264 7896 16270 7948
rect 17586 7896 17592 7948
rect 17644 7936 17650 7948
rect 17681 7939 17739 7945
rect 17681 7936 17693 7939
rect 17644 7908 17693 7936
rect 17644 7896 17650 7908
rect 17681 7905 17693 7908
rect 17727 7905 17739 7939
rect 17681 7899 17739 7905
rect 19150 7896 19156 7948
rect 19208 7936 19214 7948
rect 19429 7939 19487 7945
rect 19429 7936 19441 7939
rect 19208 7908 19441 7936
rect 19208 7896 19214 7908
rect 19429 7905 19441 7908
rect 19475 7905 19487 7939
rect 19429 7899 19487 7905
rect 19518 7896 19524 7948
rect 19576 7936 19582 7948
rect 19613 7939 19671 7945
rect 19613 7936 19625 7939
rect 19576 7908 19625 7936
rect 19576 7896 19582 7908
rect 19613 7905 19625 7908
rect 19659 7905 19671 7939
rect 19613 7899 19671 7905
rect 22741 7939 22799 7945
rect 22741 7905 22753 7939
rect 22787 7936 22799 7939
rect 23658 7936 23664 7948
rect 22787 7908 23664 7936
rect 22787 7905 22799 7908
rect 22741 7899 22799 7905
rect 23658 7896 23664 7908
rect 23716 7896 23722 7948
rect 25476 7939 25534 7945
rect 25476 7905 25488 7939
rect 25522 7936 25534 7939
rect 25682 7936 25688 7948
rect 25522 7908 25688 7936
rect 25522 7905 25534 7908
rect 25476 7899 25534 7905
rect 25682 7896 25688 7908
rect 25740 7896 25746 7948
rect 13722 7868 13728 7880
rect 13683 7840 13728 7868
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 13998 7868 14004 7880
rect 13959 7840 14004 7868
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 14826 7828 14832 7880
rect 14884 7868 14890 7880
rect 15657 7871 15715 7877
rect 15657 7868 15669 7871
rect 14884 7840 15669 7868
rect 14884 7828 14890 7840
rect 15657 7837 15669 7840
rect 15703 7868 15715 7871
rect 16574 7868 16580 7880
rect 15703 7840 16580 7868
rect 15703 7837 15715 7840
rect 15657 7831 15715 7837
rect 16574 7828 16580 7840
rect 16632 7868 16638 7880
rect 16850 7868 16856 7880
rect 16632 7840 16856 7868
rect 16632 7828 16638 7840
rect 16850 7828 16856 7840
rect 16908 7828 16914 7880
rect 21821 7871 21879 7877
rect 21821 7837 21833 7871
rect 21867 7868 21879 7871
rect 21910 7868 21916 7880
rect 21867 7840 21916 7868
rect 21867 7837 21879 7840
rect 21821 7831 21879 7837
rect 21910 7828 21916 7840
rect 21968 7828 21974 7880
rect 23934 7868 23940 7880
rect 23895 7840 23940 7868
rect 23934 7828 23940 7840
rect 23992 7828 23998 7880
rect 24394 7868 24400 7880
rect 24355 7840 24400 7868
rect 24394 7828 24400 7840
rect 24452 7828 24458 7880
rect 10410 7760 10416 7812
rect 10468 7800 10474 7812
rect 12802 7800 12808 7812
rect 10468 7772 12808 7800
rect 10468 7760 10474 7772
rect 12802 7760 12808 7772
rect 12860 7760 12866 7812
rect 15749 7803 15807 7809
rect 15749 7800 15761 7803
rect 13924 7772 15761 7800
rect 10134 7732 10140 7744
rect 10095 7704 10140 7732
rect 10134 7692 10140 7704
rect 10192 7692 10198 7744
rect 10594 7732 10600 7744
rect 10555 7704 10600 7732
rect 10594 7692 10600 7704
rect 10652 7692 10658 7744
rect 11330 7692 11336 7744
rect 11388 7732 11394 7744
rect 11425 7735 11483 7741
rect 11425 7732 11437 7735
rect 11388 7704 11437 7732
rect 11388 7692 11394 7704
rect 11425 7701 11437 7704
rect 11471 7732 11483 7735
rect 11793 7735 11851 7741
rect 11793 7732 11805 7735
rect 11471 7704 11805 7732
rect 11471 7701 11483 7704
rect 11425 7695 11483 7701
rect 11793 7701 11805 7704
rect 11839 7732 11851 7735
rect 12342 7732 12348 7744
rect 11839 7704 12348 7732
rect 11839 7701 11851 7704
rect 11793 7695 11851 7701
rect 12342 7692 12348 7704
rect 12400 7732 12406 7744
rect 13924 7732 13952 7772
rect 15749 7769 15761 7772
rect 15795 7769 15807 7803
rect 15749 7763 15807 7769
rect 12400 7704 13952 7732
rect 12400 7692 12406 7704
rect 14550 7692 14556 7744
rect 14608 7732 14614 7744
rect 15470 7741 15476 7744
rect 14645 7735 14703 7741
rect 14645 7732 14657 7735
rect 14608 7704 14657 7732
rect 14608 7692 14614 7704
rect 14645 7701 14657 7704
rect 14691 7732 14703 7735
rect 15013 7735 15071 7741
rect 15013 7732 15025 7735
rect 14691 7704 15025 7732
rect 14691 7701 14703 7704
rect 14645 7695 14703 7701
rect 15013 7701 15025 7704
rect 15059 7732 15071 7735
rect 15427 7735 15476 7741
rect 15427 7732 15439 7735
rect 15059 7704 15439 7732
rect 15059 7701 15071 7704
rect 15013 7695 15071 7701
rect 15427 7701 15439 7704
rect 15473 7701 15476 7735
rect 15427 7695 15476 7701
rect 15470 7692 15476 7695
rect 15528 7692 15534 7744
rect 15565 7735 15623 7741
rect 15565 7701 15577 7735
rect 15611 7732 15623 7735
rect 15654 7732 15660 7744
rect 15611 7704 15660 7732
rect 15611 7701 15623 7704
rect 15565 7695 15623 7701
rect 15654 7692 15660 7704
rect 15712 7732 15718 7744
rect 15930 7732 15936 7744
rect 15712 7704 15936 7732
rect 15712 7692 15718 7704
rect 15930 7692 15936 7704
rect 15988 7692 15994 7744
rect 16206 7692 16212 7744
rect 16264 7732 16270 7744
rect 16301 7735 16359 7741
rect 16301 7732 16313 7735
rect 16264 7704 16313 7732
rect 16264 7692 16270 7704
rect 16301 7701 16313 7704
rect 16347 7701 16359 7735
rect 16301 7695 16359 7701
rect 16574 7692 16580 7744
rect 16632 7732 16638 7744
rect 16669 7735 16727 7741
rect 16669 7732 16681 7735
rect 16632 7704 16681 7732
rect 16632 7692 16638 7704
rect 16669 7701 16681 7704
rect 16715 7701 16727 7735
rect 16669 7695 16727 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 7650 7528 7656 7540
rect 7611 7500 7656 7528
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 8294 7528 8300 7540
rect 8255 7500 8300 7528
rect 8294 7488 8300 7500
rect 8352 7488 8358 7540
rect 8938 7528 8944 7540
rect 8899 7500 8944 7528
rect 8938 7488 8944 7500
rect 8996 7488 9002 7540
rect 9677 7531 9735 7537
rect 9677 7497 9689 7531
rect 9723 7528 9735 7531
rect 10410 7528 10416 7540
rect 9723 7500 10416 7528
rect 9723 7497 9735 7500
rect 9677 7491 9735 7497
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 10594 7528 10600 7540
rect 10555 7500 10600 7528
rect 10594 7488 10600 7500
rect 10652 7528 10658 7540
rect 10962 7528 10968 7540
rect 10652 7500 10968 7528
rect 10652 7488 10658 7500
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11698 7488 11704 7540
rect 11756 7528 11762 7540
rect 13909 7531 13967 7537
rect 13909 7528 13921 7531
rect 11756 7500 13921 7528
rect 11756 7488 11762 7500
rect 13909 7497 13921 7500
rect 13955 7497 13967 7531
rect 13909 7491 13967 7497
rect 14277 7531 14335 7537
rect 14277 7497 14289 7531
rect 14323 7528 14335 7531
rect 14826 7528 14832 7540
rect 14323 7500 14832 7528
rect 14323 7497 14335 7500
rect 14277 7491 14335 7497
rect 9953 7463 10011 7469
rect 9953 7429 9965 7463
rect 9999 7460 10011 7463
rect 10042 7460 10048 7472
rect 9999 7432 10048 7460
rect 9999 7429 10011 7432
rect 9953 7423 10011 7429
rect 10042 7420 10048 7432
rect 10100 7420 10106 7472
rect 11425 7463 11483 7469
rect 11425 7429 11437 7463
rect 11471 7460 11483 7463
rect 13722 7460 13728 7472
rect 11471 7432 13728 7460
rect 11471 7429 11483 7432
rect 11425 7423 11483 7429
rect 1670 7352 1676 7404
rect 1728 7392 1734 7404
rect 10134 7392 10140 7404
rect 1728 7364 10140 7392
rect 1728 7352 1734 7364
rect 10134 7352 10140 7364
rect 10192 7392 10198 7404
rect 10873 7395 10931 7401
rect 10873 7392 10885 7395
rect 10192 7364 10885 7392
rect 10192 7352 10198 7364
rect 10873 7361 10885 7364
rect 10919 7361 10931 7395
rect 10873 7355 10931 7361
rect 11330 7352 11336 7404
rect 11388 7392 11394 7404
rect 13004 7401 13032 7432
rect 13722 7420 13728 7432
rect 13780 7420 13786 7472
rect 13924 7460 13952 7491
rect 14826 7488 14832 7500
rect 14884 7528 14890 7540
rect 15381 7531 15439 7537
rect 15381 7528 15393 7531
rect 14884 7500 15393 7528
rect 14884 7488 14890 7500
rect 15381 7497 15393 7500
rect 15427 7497 15439 7531
rect 15381 7491 15439 7497
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 16071 7531 16129 7537
rect 16071 7528 16083 7531
rect 15528 7500 16083 7528
rect 15528 7488 15534 7500
rect 16071 7497 16083 7500
rect 16117 7528 16129 7531
rect 17313 7531 17371 7537
rect 17313 7528 17325 7531
rect 16117 7500 17325 7528
rect 16117 7497 16129 7500
rect 16071 7491 16129 7497
rect 17313 7497 17325 7500
rect 17359 7497 17371 7531
rect 18690 7528 18696 7540
rect 18651 7500 18696 7528
rect 17313 7491 17371 7497
rect 18690 7488 18696 7500
rect 18748 7528 18754 7540
rect 18969 7531 19027 7537
rect 18969 7528 18981 7531
rect 18748 7500 18981 7528
rect 18748 7488 18754 7500
rect 18969 7497 18981 7500
rect 19015 7497 19027 7531
rect 19150 7528 19156 7540
rect 19111 7500 19156 7528
rect 18969 7491 19027 7497
rect 19150 7488 19156 7500
rect 19208 7488 19214 7540
rect 21174 7488 21180 7540
rect 21232 7528 21238 7540
rect 21821 7531 21879 7537
rect 21821 7528 21833 7531
rect 21232 7500 21833 7528
rect 21232 7488 21238 7500
rect 21821 7497 21833 7500
rect 21867 7497 21879 7531
rect 21821 7491 21879 7497
rect 22186 7488 22192 7540
rect 22244 7528 22250 7540
rect 23385 7531 23443 7537
rect 23385 7528 23397 7531
rect 22244 7500 23397 7528
rect 22244 7488 22250 7500
rect 23385 7497 23397 7500
rect 23431 7528 23443 7531
rect 24026 7528 24032 7540
rect 23431 7500 24032 7528
rect 23431 7497 23443 7500
rect 23385 7491 23443 7497
rect 24026 7488 24032 7500
rect 24084 7488 24090 7540
rect 25501 7531 25559 7537
rect 25501 7497 25513 7531
rect 25547 7528 25559 7531
rect 25682 7528 25688 7540
rect 25547 7500 25688 7528
rect 25547 7497 25559 7500
rect 25501 7491 25559 7497
rect 25682 7488 25688 7500
rect 25740 7488 25746 7540
rect 14645 7463 14703 7469
rect 14645 7460 14657 7463
rect 13924 7432 14657 7460
rect 14645 7429 14657 7432
rect 14691 7460 14703 7463
rect 15102 7460 15108 7472
rect 14691 7432 15108 7460
rect 14691 7429 14703 7432
rect 14645 7423 14703 7429
rect 15102 7420 15108 7432
rect 15160 7460 15166 7472
rect 15654 7460 15660 7472
rect 15160 7432 15660 7460
rect 15160 7420 15166 7432
rect 15654 7420 15660 7432
rect 15712 7420 15718 7472
rect 15746 7420 15752 7472
rect 15804 7460 15810 7472
rect 16209 7463 16267 7469
rect 16209 7460 16221 7463
rect 15804 7432 16221 7460
rect 15804 7420 15810 7432
rect 16209 7429 16221 7432
rect 16255 7429 16267 7463
rect 20717 7463 20775 7469
rect 20717 7460 20729 7463
rect 16209 7423 16267 7429
rect 19352 7432 20729 7460
rect 12713 7395 12771 7401
rect 12713 7392 12725 7395
rect 11388 7364 12725 7392
rect 11388 7352 11394 7364
rect 12713 7361 12725 7364
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 14182 7352 14188 7404
rect 14240 7392 14246 7404
rect 14550 7401 14556 7404
rect 14516 7395 14556 7401
rect 14516 7392 14528 7395
rect 14240 7364 14528 7392
rect 14240 7352 14246 7364
rect 14516 7361 14528 7364
rect 14516 7355 14556 7361
rect 14550 7352 14556 7355
rect 14608 7352 14614 7404
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7392 14795 7395
rect 14826 7392 14832 7404
rect 14783 7364 14832 7392
rect 14783 7361 14795 7364
rect 14737 7355 14795 7361
rect 14826 7352 14832 7364
rect 14884 7352 14890 7404
rect 15838 7392 15844 7404
rect 15751 7364 15844 7392
rect 15838 7352 15844 7364
rect 15896 7392 15902 7404
rect 16301 7395 16359 7401
rect 16301 7392 16313 7395
rect 15896 7364 16313 7392
rect 15896 7352 15902 7364
rect 16301 7361 16313 7364
rect 16347 7361 16359 7395
rect 16301 7355 16359 7361
rect 16669 7395 16727 7401
rect 16669 7361 16681 7395
rect 16715 7392 16727 7395
rect 17310 7392 17316 7404
rect 16715 7364 17316 7392
rect 16715 7361 16727 7364
rect 16669 7355 16727 7361
rect 17310 7352 17316 7364
rect 17368 7352 17374 7404
rect 19352 7401 19380 7432
rect 20717 7429 20729 7432
rect 20763 7460 20775 7463
rect 20763 7432 24716 7460
rect 20763 7429 20775 7432
rect 20717 7423 20775 7429
rect 19337 7395 19395 7401
rect 19337 7361 19349 7395
rect 19383 7361 19395 7395
rect 19337 7355 19395 7361
rect 19426 7352 19432 7404
rect 19484 7392 19490 7404
rect 19613 7395 19671 7401
rect 19613 7392 19625 7395
rect 19484 7364 19625 7392
rect 19484 7352 19490 7364
rect 19613 7361 19625 7364
rect 19659 7361 19671 7395
rect 20806 7392 20812 7404
rect 20767 7364 20812 7392
rect 19613 7355 19671 7361
rect 20806 7352 20812 7364
rect 20864 7352 20870 7404
rect 22097 7395 22155 7401
rect 22097 7361 22109 7395
rect 22143 7392 22155 7395
rect 22278 7392 22284 7404
rect 22143 7364 22284 7392
rect 22143 7361 22155 7364
rect 22097 7355 22155 7361
rect 22278 7352 22284 7364
rect 22336 7352 22342 7404
rect 22370 7352 22376 7404
rect 22428 7392 22434 7404
rect 24394 7392 24400 7404
rect 22428 7364 24400 7392
rect 22428 7352 22434 7364
rect 24394 7352 24400 7364
rect 24452 7352 24458 7404
rect 24688 7401 24716 7432
rect 24673 7395 24731 7401
rect 24673 7361 24685 7395
rect 24719 7392 24731 7395
rect 24854 7392 24860 7404
rect 24719 7364 24860 7392
rect 24719 7361 24731 7364
rect 24673 7355 24731 7361
rect 24854 7352 24860 7364
rect 24912 7352 24918 7404
rect 7812 7327 7870 7333
rect 7812 7293 7824 7327
rect 7858 7324 7870 7327
rect 8294 7324 8300 7336
rect 7858 7296 8300 7324
rect 7858 7293 7870 7296
rect 7812 7287 7870 7293
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 8757 7327 8815 7333
rect 8757 7293 8769 7327
rect 8803 7324 8815 7327
rect 8803 7296 9168 7324
rect 8803 7293 8815 7296
rect 8757 7287 8815 7293
rect 8021 7259 8079 7265
rect 8021 7225 8033 7259
rect 8067 7256 8079 7259
rect 8938 7256 8944 7268
rect 8067 7228 8944 7256
rect 8067 7225 8079 7228
rect 8021 7219 8079 7225
rect 8938 7216 8944 7228
rect 8996 7216 9002 7268
rect 9140 7200 9168 7296
rect 9398 7284 9404 7336
rect 9456 7324 9462 7336
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 9456 7296 9781 7324
rect 9456 7284 9462 7296
rect 9769 7293 9781 7296
rect 9815 7324 9827 7327
rect 11977 7327 12035 7333
rect 9815 7296 10364 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 8665 7191 8723 7197
rect 8665 7157 8677 7191
rect 8711 7188 8723 7191
rect 8846 7188 8852 7200
rect 8711 7160 8852 7188
rect 8711 7157 8723 7160
rect 8665 7151 8723 7157
rect 8846 7148 8852 7160
rect 8904 7148 8910 7200
rect 9122 7148 9128 7200
rect 9180 7188 9186 7200
rect 10336 7197 10364 7296
rect 11977 7293 11989 7327
rect 12023 7324 12035 7327
rect 12250 7324 12256 7336
rect 12023 7296 12256 7324
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 12250 7284 12256 7296
rect 12308 7284 12314 7336
rect 14366 7324 14372 7336
rect 14327 7296 14372 7324
rect 14366 7284 14372 7296
rect 14424 7324 14430 7336
rect 15933 7327 15991 7333
rect 15933 7324 15945 7327
rect 14424 7296 15945 7324
rect 14424 7284 14430 7296
rect 15933 7293 15945 7296
rect 15979 7324 15991 7327
rect 16574 7324 16580 7336
rect 15979 7296 16580 7324
rect 15979 7293 15991 7296
rect 15933 7287 15991 7293
rect 16574 7284 16580 7296
rect 16632 7284 16638 7336
rect 17773 7327 17831 7333
rect 17773 7293 17785 7327
rect 17819 7324 17831 7327
rect 17862 7324 17868 7336
rect 17819 7296 17868 7324
rect 17819 7293 17831 7296
rect 17773 7287 17831 7293
rect 17862 7284 17868 7296
rect 17920 7284 17926 7336
rect 23658 7284 23664 7336
rect 23716 7324 23722 7336
rect 24121 7327 24179 7333
rect 24121 7324 24133 7327
rect 23716 7296 24133 7324
rect 23716 7284 23722 7296
rect 24121 7293 24133 7296
rect 24167 7293 24179 7327
rect 24121 7287 24179 7293
rect 10962 7216 10968 7268
rect 11020 7256 11026 7268
rect 11020 7228 11065 7256
rect 11164 7228 12020 7256
rect 11020 7216 11026 7228
rect 9217 7191 9275 7197
rect 9217 7188 9229 7191
rect 9180 7160 9229 7188
rect 9180 7148 9186 7160
rect 9217 7157 9229 7160
rect 9263 7157 9275 7191
rect 9217 7151 9275 7157
rect 10321 7191 10379 7197
rect 10321 7157 10333 7191
rect 10367 7188 10379 7191
rect 11164 7188 11192 7228
rect 10367 7160 11192 7188
rect 11992 7188 12020 7228
rect 12802 7216 12808 7268
rect 12860 7256 12866 7268
rect 16390 7256 16396 7268
rect 12860 7228 12905 7256
rect 13786 7228 16396 7256
rect 12860 7216 12866 7228
rect 13786 7188 13814 7228
rect 16390 7216 16396 7228
rect 16448 7216 16454 7268
rect 18233 7259 18291 7265
rect 18233 7225 18245 7259
rect 18279 7256 18291 7259
rect 18874 7256 18880 7268
rect 18279 7228 18880 7256
rect 18279 7225 18291 7228
rect 18233 7219 18291 7225
rect 18874 7216 18880 7228
rect 18932 7216 18938 7268
rect 18969 7259 19027 7265
rect 18969 7225 18981 7259
rect 19015 7256 19027 7259
rect 19429 7259 19487 7265
rect 19429 7256 19441 7259
rect 19015 7228 19441 7256
rect 19015 7225 19027 7228
rect 18969 7219 19027 7225
rect 19429 7225 19441 7228
rect 19475 7225 19487 7259
rect 19429 7219 19487 7225
rect 21545 7259 21603 7265
rect 21545 7225 21557 7259
rect 21591 7256 21603 7259
rect 22094 7256 22100 7268
rect 21591 7228 22100 7256
rect 21591 7225 21603 7228
rect 21545 7219 21603 7225
rect 22094 7216 22100 7228
rect 22152 7256 22158 7268
rect 22189 7259 22247 7265
rect 22189 7256 22201 7259
rect 22152 7228 22201 7256
rect 22152 7216 22158 7228
rect 22189 7225 22201 7228
rect 22235 7225 22247 7259
rect 22738 7256 22744 7268
rect 22699 7228 22744 7256
rect 22189 7219 22247 7225
rect 22738 7216 22744 7228
rect 22796 7216 22802 7268
rect 24136 7256 24164 7287
rect 24489 7259 24547 7265
rect 24489 7256 24501 7259
rect 24136 7228 24501 7256
rect 24489 7225 24501 7228
rect 24535 7225 24547 7259
rect 24489 7219 24547 7225
rect 11992 7160 13814 7188
rect 10367 7157 10379 7160
rect 10321 7151 10379 7157
rect 14274 7148 14280 7200
rect 14332 7188 14338 7200
rect 15013 7191 15071 7197
rect 15013 7188 15025 7191
rect 14332 7160 15025 7188
rect 14332 7148 14338 7160
rect 15013 7157 15025 7160
rect 15059 7157 15071 7191
rect 15013 7151 15071 7157
rect 15838 7148 15844 7200
rect 15896 7188 15902 7200
rect 16206 7188 16212 7200
rect 15896 7160 16212 7188
rect 15896 7148 15902 7160
rect 16206 7148 16212 7160
rect 16264 7188 16270 7200
rect 16945 7191 17003 7197
rect 16945 7188 16957 7191
rect 16264 7160 16957 7188
rect 16264 7148 16270 7160
rect 16945 7157 16957 7160
rect 16991 7157 17003 7191
rect 16945 7151 17003 7157
rect 17770 7148 17776 7200
rect 17828 7188 17834 7200
rect 19518 7188 19524 7200
rect 17828 7160 19524 7188
rect 17828 7148 17834 7160
rect 19518 7148 19524 7160
rect 19576 7188 19582 7200
rect 20257 7191 20315 7197
rect 20257 7188 20269 7191
rect 19576 7160 20269 7188
rect 19576 7148 19582 7160
rect 20257 7157 20269 7160
rect 20303 7157 20315 7191
rect 20257 7151 20315 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 6822 6984 6828 6996
rect 6783 6956 6828 6984
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 8754 6984 8760 6996
rect 8715 6956 8760 6984
rect 8754 6944 8760 6956
rect 8812 6944 8818 6996
rect 11241 6987 11299 6993
rect 11241 6953 11253 6987
rect 11287 6984 11299 6987
rect 11514 6984 11520 6996
rect 11287 6956 11520 6984
rect 11287 6953 11299 6956
rect 11241 6947 11299 6953
rect 11514 6944 11520 6956
rect 11572 6944 11578 6996
rect 11701 6987 11759 6993
rect 11701 6953 11713 6987
rect 11747 6984 11759 6987
rect 11882 6984 11888 6996
rect 11747 6956 11888 6984
rect 11747 6953 11759 6956
rect 11701 6947 11759 6953
rect 11882 6944 11888 6956
rect 11940 6984 11946 6996
rect 12250 6984 12256 6996
rect 11940 6956 12256 6984
rect 11940 6944 11946 6956
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12713 6987 12771 6993
rect 12713 6953 12725 6987
rect 12759 6984 12771 6987
rect 12802 6984 12808 6996
rect 12759 6956 12808 6984
rect 12759 6953 12771 6956
rect 12713 6947 12771 6953
rect 12802 6944 12808 6956
rect 12860 6944 12866 6996
rect 13170 6984 13176 6996
rect 13131 6956 13176 6984
rect 13170 6944 13176 6956
rect 13228 6944 13234 6996
rect 14366 6984 14372 6996
rect 14327 6956 14372 6984
rect 14366 6944 14372 6956
rect 14424 6944 14430 6996
rect 15102 6984 15108 6996
rect 15063 6956 15108 6984
rect 15102 6944 15108 6956
rect 15160 6944 15166 6996
rect 15746 6944 15752 6996
rect 15804 6984 15810 6996
rect 15933 6987 15991 6993
rect 15933 6984 15945 6987
rect 15804 6956 15945 6984
rect 15804 6944 15810 6956
rect 15933 6953 15945 6956
rect 15979 6953 15991 6987
rect 17310 6984 17316 6996
rect 17271 6956 17316 6984
rect 15933 6947 15991 6953
rect 17310 6944 17316 6956
rect 17368 6944 17374 6996
rect 17586 6944 17592 6996
rect 17644 6984 17650 6996
rect 17681 6987 17739 6993
rect 17681 6984 17693 6987
rect 17644 6956 17693 6984
rect 17644 6944 17650 6956
rect 17681 6953 17693 6956
rect 17727 6953 17739 6987
rect 17681 6947 17739 6953
rect 21174 6944 21180 6996
rect 21232 6984 21238 6996
rect 21269 6987 21327 6993
rect 21269 6984 21281 6987
rect 21232 6956 21281 6984
rect 21232 6944 21238 6956
rect 21269 6953 21281 6956
rect 21315 6953 21327 6987
rect 23934 6984 23940 6996
rect 23895 6956 23940 6984
rect 21269 6947 21327 6953
rect 23934 6944 23940 6956
rect 23992 6944 23998 6996
rect 24394 6984 24400 6996
rect 24355 6956 24400 6984
rect 24394 6944 24400 6956
rect 24452 6944 24458 6996
rect 7699 6919 7757 6925
rect 7699 6885 7711 6919
rect 7745 6916 7757 6919
rect 10781 6919 10839 6925
rect 10781 6916 10793 6919
rect 7745 6888 10793 6916
rect 7745 6885 7757 6888
rect 7699 6879 7757 6885
rect 10781 6885 10793 6888
rect 10827 6916 10839 6919
rect 11330 6916 11336 6928
rect 10827 6888 11336 6916
rect 10827 6885 10839 6888
rect 10781 6879 10839 6885
rect 11330 6876 11336 6888
rect 11388 6876 11394 6928
rect 13814 6876 13820 6928
rect 13872 6916 13878 6928
rect 13872 6888 16344 6916
rect 13872 6876 13878 6888
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 6638 6848 6644 6860
rect 6595 6820 6644 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 6638 6808 6644 6820
rect 6696 6808 6702 6860
rect 7558 6848 7564 6860
rect 7522 6820 7564 6848
rect 7558 6808 7564 6820
rect 7616 6857 7622 6860
rect 7616 6851 7670 6857
rect 7616 6817 7624 6851
rect 7658 6848 7670 6851
rect 8110 6848 8116 6860
rect 7658 6820 8116 6848
rect 7658 6817 7670 6820
rect 7616 6811 7670 6817
rect 7616 6808 7622 6811
rect 8110 6808 8116 6820
rect 8168 6808 8174 6860
rect 8294 6808 8300 6860
rect 8352 6848 8358 6860
rect 8573 6851 8631 6857
rect 8573 6848 8585 6851
rect 8352 6820 8585 6848
rect 8352 6808 8358 6820
rect 8573 6817 8585 6820
rect 8619 6817 8631 6851
rect 9122 6848 9128 6860
rect 9083 6820 9128 6848
rect 8573 6811 8631 6817
rect 9122 6808 9128 6820
rect 9180 6808 9186 6860
rect 10134 6848 10140 6860
rect 10095 6820 10140 6848
rect 10134 6808 10140 6820
rect 10192 6848 10198 6860
rect 12158 6848 12164 6860
rect 10192 6820 12164 6848
rect 10192 6808 10198 6820
rect 12158 6808 12164 6820
rect 12216 6848 12222 6860
rect 12253 6851 12311 6857
rect 12253 6848 12265 6851
rect 12216 6820 12265 6848
rect 12216 6808 12222 6820
rect 12253 6817 12265 6820
rect 12299 6817 12311 6851
rect 13354 6848 13360 6860
rect 13315 6820 13360 6848
rect 12253 6811 12311 6817
rect 13354 6808 13360 6820
rect 13412 6808 13418 6860
rect 13633 6851 13691 6857
rect 13633 6817 13645 6851
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6780 10563 6783
rect 11054 6780 11060 6792
rect 10551 6752 11060 6780
rect 10551 6749 10563 6752
rect 10505 6743 10563 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11333 6783 11391 6789
rect 11333 6749 11345 6783
rect 11379 6780 11391 6783
rect 12526 6780 12532 6792
rect 11379 6752 12532 6780
rect 11379 6749 11391 6752
rect 11333 6743 11391 6749
rect 12526 6740 12532 6752
rect 12584 6740 12590 6792
rect 13648 6780 13676 6811
rect 14826 6808 14832 6860
rect 14884 6848 14890 6860
rect 15286 6848 15292 6860
rect 14884 6820 15292 6848
rect 14884 6808 14890 6820
rect 15286 6808 15292 6820
rect 15344 6808 15350 6860
rect 16316 6857 16344 6888
rect 16301 6851 16359 6857
rect 16301 6817 16313 6851
rect 16347 6848 16359 6851
rect 16758 6848 16764 6860
rect 16347 6820 16764 6848
rect 16347 6817 16359 6820
rect 16301 6811 16359 6817
rect 16758 6808 16764 6820
rect 16816 6808 16822 6860
rect 16853 6851 16911 6857
rect 16853 6817 16865 6851
rect 16899 6848 16911 6851
rect 17328 6848 17356 6944
rect 23106 6916 23112 6928
rect 23067 6888 23112 6916
rect 23106 6876 23112 6888
rect 23164 6876 23170 6928
rect 24670 6916 24676 6928
rect 24631 6888 24676 6916
rect 24670 6876 24676 6888
rect 24728 6876 24734 6928
rect 17862 6848 17868 6860
rect 16899 6820 17356 6848
rect 17823 6820 17868 6848
rect 16899 6817 16911 6820
rect 16853 6811 16911 6817
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 19058 6848 19064 6860
rect 19019 6820 19064 6848
rect 19058 6808 19064 6820
rect 19116 6808 19122 6860
rect 19242 6808 19248 6860
rect 19300 6848 19306 6860
rect 19705 6851 19763 6857
rect 19705 6848 19717 6851
rect 19300 6820 19717 6848
rect 19300 6808 19306 6820
rect 19705 6817 19717 6820
rect 19751 6817 19763 6851
rect 19886 6848 19892 6860
rect 19847 6820 19892 6848
rect 19705 6811 19763 6817
rect 19886 6808 19892 6820
rect 19944 6808 19950 6860
rect 21910 6848 21916 6860
rect 20317 6820 21916 6848
rect 14274 6780 14280 6792
rect 13648 6752 14280 6780
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 15838 6780 15844 6792
rect 14660 6752 15844 6780
rect 9490 6712 9496 6724
rect 9451 6684 9496 6712
rect 9490 6672 9496 6684
rect 9548 6672 9554 6724
rect 7098 6644 7104 6656
rect 7059 6616 7104 6644
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 8113 6647 8171 6653
rect 8113 6613 8125 6647
rect 8159 6644 8171 6647
rect 8570 6644 8576 6656
rect 8159 6616 8576 6644
rect 8159 6613 8171 6616
rect 8113 6607 8171 6613
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 8846 6604 8852 6656
rect 8904 6644 8910 6656
rect 14660 6644 14688 6752
rect 15838 6740 15844 6752
rect 15896 6740 15902 6792
rect 17037 6783 17095 6789
rect 17037 6749 17049 6783
rect 17083 6780 17095 6783
rect 20317 6780 20345 6820
rect 21910 6808 21916 6820
rect 21968 6848 21974 6860
rect 22465 6851 22523 6857
rect 22465 6848 22477 6851
rect 21968 6820 22477 6848
rect 21968 6808 21974 6820
rect 22465 6817 22477 6820
rect 22511 6817 22523 6851
rect 22465 6811 22523 6817
rect 20898 6780 20904 6792
rect 17083 6752 20345 6780
rect 20859 6752 20904 6780
rect 17083 6749 17095 6752
rect 17037 6743 17095 6749
rect 20898 6740 20904 6752
rect 20956 6740 20962 6792
rect 23014 6780 23020 6792
rect 22975 6752 23020 6780
rect 23014 6740 23020 6752
rect 23072 6740 23078 6792
rect 24210 6740 24216 6792
rect 24268 6780 24274 6792
rect 24581 6783 24639 6789
rect 24581 6780 24593 6783
rect 24268 6752 24593 6780
rect 24268 6740 24274 6752
rect 24581 6749 24593 6752
rect 24627 6749 24639 6783
rect 24854 6780 24860 6792
rect 24815 6752 24860 6780
rect 24581 6743 24639 6749
rect 24854 6740 24860 6752
rect 24912 6740 24918 6792
rect 18690 6712 18696 6724
rect 15488 6684 18696 6712
rect 15488 6656 15516 6684
rect 18690 6672 18696 6684
rect 18748 6672 18754 6724
rect 23566 6712 23572 6724
rect 23527 6684 23572 6712
rect 23566 6672 23572 6684
rect 23624 6672 23630 6724
rect 15470 6644 15476 6656
rect 8904 6616 14688 6644
rect 15431 6616 15476 6644
rect 8904 6604 8910 6616
rect 15470 6604 15476 6616
rect 15528 6604 15534 6656
rect 18049 6647 18107 6653
rect 18049 6613 18061 6647
rect 18095 6644 18107 6647
rect 18414 6644 18420 6656
rect 18095 6616 18420 6644
rect 18095 6613 18107 6616
rect 18049 6607 18107 6613
rect 18414 6604 18420 6616
rect 18472 6604 18478 6656
rect 19978 6604 19984 6656
rect 20036 6644 20042 6656
rect 20036 6616 20081 6644
rect 20036 6604 20042 6616
rect 21266 6604 21272 6656
rect 21324 6644 21330 6656
rect 21818 6644 21824 6656
rect 21324 6616 21824 6644
rect 21324 6604 21330 6616
rect 21818 6604 21824 6616
rect 21876 6604 21882 6656
rect 22189 6647 22247 6653
rect 22189 6613 22201 6647
rect 22235 6644 22247 6647
rect 22278 6644 22284 6656
rect 22235 6616 22284 6644
rect 22235 6613 22247 6616
rect 22189 6607 22247 6613
rect 22278 6604 22284 6616
rect 22336 6604 22342 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 6638 6440 6644 6452
rect 6599 6412 6644 6440
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 7558 6440 7564 6452
rect 7519 6412 7564 6440
rect 7558 6400 7564 6412
rect 7616 6400 7622 6452
rect 9198 6443 9256 6449
rect 9198 6409 9210 6443
rect 9244 6440 9256 6443
rect 9490 6440 9496 6452
rect 9244 6412 9496 6440
rect 9244 6409 9256 6412
rect 9198 6403 9256 6409
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 10134 6440 10140 6452
rect 10095 6412 10140 6440
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 10505 6443 10563 6449
rect 10505 6409 10517 6443
rect 10551 6440 10563 6443
rect 10962 6440 10968 6452
rect 10551 6412 10968 6440
rect 10551 6409 10563 6412
rect 10505 6403 10563 6409
rect 10962 6400 10968 6412
rect 11020 6440 11026 6452
rect 11882 6440 11888 6452
rect 11020 6412 11888 6440
rect 11020 6400 11026 6412
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 11974 6400 11980 6452
rect 12032 6440 12038 6452
rect 12161 6443 12219 6449
rect 12161 6440 12173 6443
rect 12032 6412 12173 6440
rect 12032 6400 12038 6412
rect 12161 6409 12173 6412
rect 12207 6409 12219 6443
rect 12161 6403 12219 6409
rect 13354 6400 13360 6452
rect 13412 6440 13418 6452
rect 13449 6443 13507 6449
rect 13449 6440 13461 6443
rect 13412 6412 13461 6440
rect 13412 6400 13418 6412
rect 13449 6409 13461 6412
rect 13495 6409 13507 6443
rect 13449 6403 13507 6409
rect 13909 6443 13967 6449
rect 13909 6409 13921 6443
rect 13955 6440 13967 6443
rect 14274 6440 14280 6452
rect 13955 6412 14280 6440
rect 13955 6409 13967 6412
rect 13909 6403 13967 6409
rect 9306 6372 9312 6384
rect 9267 6344 9312 6372
rect 9306 6332 9312 6344
rect 9364 6332 9370 6384
rect 13464 6372 13492 6403
rect 13814 6372 13820 6384
rect 13464 6344 13820 6372
rect 13814 6332 13820 6344
rect 13872 6332 13878 6384
rect 8570 6304 8576 6316
rect 8036 6276 8576 6304
rect 6917 6239 6975 6245
rect 6917 6205 6929 6239
rect 6963 6236 6975 6239
rect 7098 6236 7104 6248
rect 6963 6208 7104 6236
rect 6963 6205 6975 6208
rect 6917 6199 6975 6205
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 8036 6245 8064 6276
rect 8570 6264 8576 6276
rect 8628 6264 8634 6316
rect 9398 6304 9404 6316
rect 9359 6276 9404 6304
rect 9398 6264 9404 6276
rect 9456 6264 9462 6316
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6304 10655 6307
rect 10686 6304 10692 6316
rect 10643 6276 10692 6304
rect 10643 6273 10655 6276
rect 10597 6267 10655 6273
rect 10686 6264 10692 6276
rect 10744 6304 10750 6316
rect 13170 6304 13176 6316
rect 10744 6276 13176 6304
rect 10744 6264 10750 6276
rect 13170 6264 13176 6276
rect 13228 6264 13234 6316
rect 8036 6239 8114 6245
rect 8036 6208 8068 6239
rect 8056 6205 8068 6208
rect 8102 6205 8114 6239
rect 8056 6199 8114 6205
rect 8159 6239 8217 6245
rect 8159 6205 8171 6239
rect 8205 6236 8217 6239
rect 10502 6236 10508 6248
rect 8205 6208 10508 6236
rect 8205 6205 8217 6208
rect 8159 6199 8217 6205
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 11974 6196 11980 6248
rect 12032 6236 12038 6248
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 12032 6208 12449 6236
rect 12032 6196 12038 6208
rect 12437 6205 12449 6208
rect 12483 6205 12495 6239
rect 12437 6199 12495 6205
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 12989 6239 13047 6245
rect 12989 6236 13001 6239
rect 12768 6208 13001 6236
rect 12768 6196 12774 6208
rect 12989 6205 13001 6208
rect 13035 6236 13047 6239
rect 13924 6236 13952 6403
rect 14274 6400 14280 6412
rect 14332 6400 14338 6452
rect 14550 6400 14556 6452
rect 14608 6440 14614 6452
rect 16114 6440 16120 6452
rect 14608 6412 16120 6440
rect 14608 6400 14614 6412
rect 16114 6400 16120 6412
rect 16172 6449 16178 6452
rect 16172 6443 16221 6449
rect 16172 6409 16175 6443
rect 16209 6409 16221 6443
rect 16298 6440 16304 6452
rect 16259 6412 16304 6440
rect 16172 6403 16221 6409
rect 16172 6400 16206 6403
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 16758 6400 16764 6452
rect 16816 6440 16822 6452
rect 17405 6443 17463 6449
rect 17405 6440 17417 6443
rect 16816 6412 17417 6440
rect 16816 6400 16822 6412
rect 17405 6409 17417 6412
rect 17451 6409 17463 6443
rect 24670 6440 24676 6452
rect 24631 6412 24676 6440
rect 17405 6403 17463 6409
rect 24670 6400 24676 6412
rect 24728 6400 24734 6452
rect 16178 6372 16206 6400
rect 17773 6375 17831 6381
rect 17773 6372 17785 6375
rect 16178 6344 17785 6372
rect 17773 6341 17785 6344
rect 17819 6341 17831 6375
rect 17773 6335 17831 6341
rect 22005 6375 22063 6381
rect 22005 6341 22017 6375
rect 22051 6372 22063 6375
rect 23017 6375 23075 6381
rect 23017 6372 23029 6375
rect 22051 6344 23029 6372
rect 22051 6341 22063 6344
rect 22005 6335 22063 6341
rect 23017 6341 23029 6344
rect 23063 6372 23075 6375
rect 23106 6372 23112 6384
rect 23063 6344 23112 6372
rect 23063 6341 23075 6344
rect 23017 6335 23075 6341
rect 23106 6332 23112 6344
rect 23164 6372 23170 6384
rect 23164 6344 23520 6372
rect 23164 6332 23170 6344
rect 15470 6304 15476 6316
rect 14476 6276 15476 6304
rect 14476 6245 14504 6276
rect 15470 6264 15476 6276
rect 15528 6264 15534 6316
rect 16390 6304 16396 6316
rect 16351 6276 16396 6304
rect 16390 6264 16396 6276
rect 16448 6304 16454 6316
rect 17037 6307 17095 6313
rect 17037 6304 17049 6307
rect 16448 6276 17049 6304
rect 16448 6264 16454 6276
rect 17037 6273 17049 6276
rect 17083 6273 17095 6307
rect 19886 6304 19892 6316
rect 19847 6276 19892 6304
rect 17037 6267 17095 6273
rect 19886 6264 19892 6276
rect 19944 6264 19950 6316
rect 19978 6264 19984 6316
rect 20036 6304 20042 6316
rect 23492 6313 23520 6344
rect 24210 6332 24216 6384
rect 24268 6372 24274 6384
rect 25041 6375 25099 6381
rect 25041 6372 25053 6375
rect 24268 6344 25053 6372
rect 24268 6332 24274 6344
rect 25041 6341 25053 6344
rect 25087 6341 25099 6375
rect 25041 6335 25099 6341
rect 25409 6375 25467 6381
rect 25409 6341 25421 6375
rect 25455 6372 25467 6375
rect 26786 6372 26792 6384
rect 25455 6344 26792 6372
rect 25455 6341 25467 6344
rect 25409 6335 25467 6341
rect 26786 6332 26792 6344
rect 26844 6332 26850 6384
rect 21085 6307 21143 6313
rect 21085 6304 21097 6307
rect 20036 6276 21097 6304
rect 20036 6264 20042 6276
rect 21085 6273 21097 6276
rect 21131 6304 21143 6307
rect 22281 6307 22339 6313
rect 22281 6304 22293 6307
rect 21131 6276 22293 6304
rect 21131 6273 21143 6276
rect 21085 6267 21143 6273
rect 22281 6273 22293 6276
rect 22327 6273 22339 6307
rect 22281 6267 22339 6273
rect 23477 6307 23535 6313
rect 23477 6273 23489 6307
rect 23523 6273 23535 6307
rect 23477 6267 23535 6273
rect 14461 6239 14519 6245
rect 14461 6236 14473 6239
rect 13035 6208 13952 6236
rect 14292 6208 14473 6236
rect 13035 6205 13047 6208
rect 12989 6199 13047 6205
rect 9030 6168 9036 6180
rect 8991 6140 9036 6168
rect 9030 6128 9036 6140
rect 9088 6128 9094 6180
rect 7147 6103 7205 6109
rect 7147 6069 7159 6103
rect 7193 6100 7205 6103
rect 7374 6100 7380 6112
rect 7193 6072 7380 6100
rect 7193 6069 7205 6072
rect 7147 6063 7205 6069
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 8573 6103 8631 6109
rect 8573 6100 8585 6103
rect 8352 6072 8585 6100
rect 8352 6060 8358 6072
rect 8573 6069 8585 6072
rect 8619 6069 8631 6103
rect 9674 6100 9680 6112
rect 9635 6072 9680 6100
rect 8573 6063 8631 6069
rect 9674 6060 9680 6072
rect 9732 6060 9738 6112
rect 10962 6100 10968 6112
rect 10923 6072 10968 6100
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 11514 6100 11520 6112
rect 11475 6072 11520 6100
rect 11514 6060 11520 6072
rect 11572 6060 11578 6112
rect 12526 6100 12532 6112
rect 12487 6072 12532 6100
rect 12526 6060 12532 6072
rect 12584 6060 12590 6112
rect 13170 6060 13176 6112
rect 13228 6100 13234 6112
rect 14292 6109 14320 6208
rect 14461 6205 14473 6208
rect 14507 6205 14519 6239
rect 14461 6199 14519 6205
rect 15013 6239 15071 6245
rect 15013 6205 15025 6239
rect 15059 6236 15071 6239
rect 15102 6236 15108 6248
rect 15059 6208 15108 6236
rect 15059 6205 15071 6208
rect 15013 6199 15071 6205
rect 15102 6196 15108 6208
rect 15160 6236 15166 6248
rect 18509 6239 18567 6245
rect 15160 6208 16804 6236
rect 15160 6196 15166 6208
rect 15197 6171 15255 6177
rect 15197 6137 15209 6171
rect 15243 6168 15255 6171
rect 15930 6168 15936 6180
rect 15243 6140 15936 6168
rect 15243 6137 15255 6140
rect 15197 6131 15255 6137
rect 15930 6128 15936 6140
rect 15988 6128 15994 6180
rect 16776 6177 16804 6208
rect 18509 6205 18521 6239
rect 18555 6236 18567 6239
rect 18877 6239 18935 6245
rect 18877 6236 18889 6239
rect 18555 6208 18889 6236
rect 18555 6205 18567 6208
rect 18509 6199 18567 6205
rect 18877 6205 18889 6208
rect 18923 6236 18935 6239
rect 18969 6239 19027 6245
rect 18969 6236 18981 6239
rect 18923 6208 18981 6236
rect 18923 6205 18935 6208
rect 18877 6199 18935 6205
rect 18969 6205 18981 6208
rect 19015 6236 19027 6239
rect 19058 6236 19064 6248
rect 19015 6208 19064 6236
rect 19015 6205 19027 6208
rect 18969 6199 19027 6205
rect 19058 6196 19064 6208
rect 19116 6196 19122 6248
rect 19518 6196 19524 6248
rect 19576 6236 19582 6248
rect 19797 6239 19855 6245
rect 19797 6236 19809 6239
rect 19576 6208 19809 6236
rect 19576 6196 19582 6208
rect 19797 6205 19809 6208
rect 19843 6205 19855 6239
rect 19797 6199 19855 6205
rect 20073 6239 20131 6245
rect 20073 6205 20085 6239
rect 20119 6236 20131 6239
rect 20898 6236 20904 6248
rect 20119 6208 20904 6236
rect 20119 6205 20131 6208
rect 20073 6199 20131 6205
rect 20898 6196 20904 6208
rect 20956 6196 20962 6248
rect 23492 6236 23520 6267
rect 23753 6239 23811 6245
rect 23753 6236 23765 6239
rect 23492 6208 23765 6236
rect 23753 6205 23765 6208
rect 23799 6205 23811 6239
rect 25222 6236 25228 6248
rect 25183 6208 25228 6236
rect 23753 6199 23811 6205
rect 25222 6196 25228 6208
rect 25280 6236 25286 6248
rect 25777 6239 25835 6245
rect 25777 6236 25789 6239
rect 25280 6208 25789 6236
rect 25280 6196 25286 6208
rect 25777 6205 25789 6208
rect 25823 6205 25835 6239
rect 25777 6199 25835 6205
rect 16025 6171 16083 6177
rect 16025 6137 16037 6171
rect 16071 6137 16083 6171
rect 16025 6131 16083 6137
rect 16761 6171 16819 6177
rect 16761 6137 16773 6171
rect 16807 6168 16819 6171
rect 17126 6168 17132 6180
rect 16807 6140 17132 6168
rect 16807 6137 16819 6140
rect 16761 6131 16819 6137
rect 14277 6103 14335 6109
rect 14277 6100 14289 6103
rect 13228 6072 14289 6100
rect 13228 6060 13234 6072
rect 14277 6069 14289 6072
rect 14323 6069 14335 6103
rect 14277 6063 14335 6069
rect 14826 6060 14832 6112
rect 14884 6100 14890 6112
rect 15473 6103 15531 6109
rect 15473 6100 15485 6103
rect 14884 6072 15485 6100
rect 14884 6060 14890 6072
rect 15473 6069 15485 6072
rect 15519 6069 15531 6103
rect 15838 6100 15844 6112
rect 15799 6072 15844 6100
rect 15473 6063 15531 6069
rect 15838 6060 15844 6072
rect 15896 6100 15902 6112
rect 16040 6100 16068 6131
rect 17126 6128 17132 6140
rect 17184 6128 17190 6180
rect 17770 6128 17776 6180
rect 17828 6168 17834 6180
rect 20533 6171 20591 6177
rect 20533 6168 20545 6171
rect 17828 6140 20545 6168
rect 17828 6128 17834 6140
rect 20533 6137 20545 6140
rect 20579 6168 20591 6171
rect 20993 6171 21051 6177
rect 20993 6168 21005 6171
rect 20579 6140 21005 6168
rect 20579 6137 20591 6140
rect 20533 6131 20591 6137
rect 20993 6137 21005 6140
rect 21039 6168 21051 6171
rect 21174 6168 21180 6180
rect 21039 6140 21180 6168
rect 21039 6137 21051 6140
rect 20993 6131 21051 6137
rect 21174 6128 21180 6140
rect 21232 6168 21238 6180
rect 21406 6171 21464 6177
rect 21406 6168 21418 6171
rect 21232 6140 21418 6168
rect 21232 6128 21238 6140
rect 21406 6137 21418 6140
rect 21452 6137 21464 6171
rect 23658 6168 23664 6180
rect 23619 6140 23664 6168
rect 21406 6131 21464 6137
rect 23658 6128 23664 6140
rect 23716 6128 23722 6180
rect 15896 6072 16068 6100
rect 15896 6060 15902 6072
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 9030 5896 9036 5908
rect 8991 5868 9036 5896
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 9398 5896 9404 5908
rect 9359 5868 9404 5896
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 10686 5896 10692 5908
rect 10647 5868 10692 5896
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 12161 5899 12219 5905
rect 12161 5865 12173 5899
rect 12207 5896 12219 5899
rect 12526 5896 12532 5908
rect 12207 5868 12532 5896
rect 12207 5865 12219 5868
rect 12161 5859 12219 5865
rect 12526 5856 12532 5868
rect 12584 5856 12590 5908
rect 13722 5896 13728 5908
rect 13683 5868 13728 5896
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 15102 5896 15108 5908
rect 15063 5868 15108 5896
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 16117 5899 16175 5905
rect 16117 5865 16129 5899
rect 16163 5896 16175 5899
rect 16298 5896 16304 5908
rect 16163 5868 16304 5896
rect 16163 5865 16175 5868
rect 16117 5859 16175 5865
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 20898 5856 20904 5908
rect 20956 5896 20962 5908
rect 21085 5899 21143 5905
rect 21085 5896 21097 5899
rect 20956 5868 21097 5896
rect 20956 5856 20962 5868
rect 21085 5865 21097 5868
rect 21131 5865 21143 5899
rect 23014 5896 23020 5908
rect 22975 5868 23020 5896
rect 21085 5859 21143 5865
rect 23014 5856 23020 5868
rect 23072 5856 23078 5908
rect 7147 5831 7205 5837
rect 7147 5797 7159 5831
rect 7193 5828 7205 5831
rect 11146 5828 11152 5840
rect 7193 5800 11152 5828
rect 7193 5797 7205 5800
rect 7147 5791 7205 5797
rect 11146 5788 11152 5800
rect 11204 5788 11210 5840
rect 11241 5831 11299 5837
rect 11241 5797 11253 5831
rect 11287 5828 11299 5831
rect 11514 5828 11520 5840
rect 11287 5800 11520 5828
rect 11287 5797 11299 5800
rect 11241 5791 11299 5797
rect 11514 5788 11520 5800
rect 11572 5788 11578 5840
rect 12437 5831 12495 5837
rect 12437 5797 12449 5831
rect 12483 5828 12495 5831
rect 12710 5828 12716 5840
rect 12483 5800 12716 5828
rect 12483 5797 12495 5800
rect 12437 5791 12495 5797
rect 12710 5788 12716 5800
rect 12768 5788 12774 5840
rect 12802 5788 12808 5840
rect 12860 5828 12866 5840
rect 18414 5828 18420 5840
rect 12860 5800 12905 5828
rect 18327 5800 18420 5828
rect 12860 5788 12866 5800
rect 18414 5788 18420 5800
rect 18472 5828 18478 5840
rect 18472 5800 19932 5828
rect 18472 5788 18478 5800
rect 6064 5763 6122 5769
rect 6064 5729 6076 5763
rect 6110 5760 6122 5763
rect 6638 5760 6644 5772
rect 6110 5732 6644 5760
rect 6110 5729 6122 5732
rect 6064 5723 6122 5729
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 7060 5763 7118 5769
rect 7060 5729 7072 5763
rect 7106 5760 7118 5763
rect 7282 5760 7288 5772
rect 7106 5732 7288 5760
rect 7106 5729 7118 5732
rect 7060 5723 7118 5729
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5760 8079 5763
rect 8478 5760 8484 5772
rect 8067 5732 8484 5760
rect 8067 5729 8079 5732
rect 8021 5723 8079 5729
rect 8478 5720 8484 5732
rect 8536 5760 8542 5772
rect 10042 5760 10048 5772
rect 8536 5732 9076 5760
rect 10003 5732 10048 5760
rect 8536 5720 8542 5732
rect 9048 5704 9076 5732
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 10183 5763 10241 5769
rect 10183 5729 10195 5763
rect 10229 5760 10241 5763
rect 10778 5760 10784 5772
rect 10229 5732 10784 5760
rect 10229 5729 10241 5732
rect 10183 5723 10241 5729
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 15286 5760 15292 5772
rect 15247 5732 15292 5760
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 17037 5763 17095 5769
rect 17037 5729 17049 5763
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 6178 5692 6184 5704
rect 6150 5652 6184 5692
rect 6236 5652 6242 5704
rect 8386 5692 8392 5704
rect 8347 5664 8392 5692
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 9030 5652 9036 5704
rect 9088 5652 9094 5704
rect 11238 5652 11244 5704
rect 11296 5692 11302 5704
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 11296 5664 11805 5692
rect 11296 5652 11302 5664
rect 11793 5661 11805 5664
rect 11839 5692 11851 5695
rect 12710 5692 12716 5704
rect 11839 5664 12716 5692
rect 11839 5661 11851 5664
rect 11793 5655 11851 5661
rect 12710 5652 12716 5664
rect 12768 5652 12774 5704
rect 12989 5695 13047 5701
rect 12989 5661 13001 5695
rect 13035 5661 13047 5695
rect 14185 5695 14243 5701
rect 14185 5692 14197 5695
rect 12989 5655 13047 5661
rect 13786 5664 14197 5692
rect 6150 5565 6178 5652
rect 7466 5584 7472 5636
rect 7524 5624 7530 5636
rect 8186 5627 8244 5633
rect 8186 5624 8198 5627
rect 7524 5596 8198 5624
rect 7524 5584 7530 5596
rect 8186 5593 8198 5596
rect 8232 5624 8244 5627
rect 9214 5624 9220 5636
rect 8232 5596 9220 5624
rect 8232 5593 8244 5596
rect 8186 5587 8244 5593
rect 9214 5584 9220 5596
rect 9272 5584 9278 5636
rect 12434 5584 12440 5636
rect 12492 5624 12498 5636
rect 13004 5624 13032 5655
rect 12492 5596 13032 5624
rect 12492 5584 12498 5596
rect 6135 5559 6193 5565
rect 6135 5525 6147 5559
rect 6181 5525 6193 5559
rect 7650 5556 7656 5568
rect 7611 5528 7656 5556
rect 6135 5519 6193 5525
rect 7650 5516 7656 5528
rect 7708 5516 7714 5568
rect 8294 5556 8300 5568
rect 8255 5528 8300 5556
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 8662 5556 8668 5568
rect 8623 5528 8668 5556
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 11606 5516 11612 5568
rect 11664 5556 11670 5568
rect 13786 5556 13814 5664
rect 14185 5661 14197 5664
rect 14231 5661 14243 5695
rect 14185 5655 14243 5661
rect 15654 5652 15660 5704
rect 15712 5692 15718 5704
rect 16393 5695 16451 5701
rect 16393 5692 16405 5695
rect 15712 5664 16405 5692
rect 15712 5652 15718 5664
rect 16393 5661 16405 5664
rect 16439 5661 16451 5695
rect 17052 5692 17080 5723
rect 18322 5720 18328 5772
rect 18380 5760 18386 5772
rect 18877 5763 18935 5769
rect 18877 5760 18889 5763
rect 18380 5732 18889 5760
rect 18380 5720 18386 5732
rect 18877 5729 18889 5732
rect 18923 5729 18935 5763
rect 19518 5760 19524 5772
rect 18877 5723 18935 5729
rect 19260 5732 19524 5760
rect 17310 5692 17316 5704
rect 17052 5664 17316 5692
rect 16393 5655 16451 5661
rect 17310 5652 17316 5664
rect 17368 5692 17374 5704
rect 18506 5692 18512 5704
rect 17368 5664 18512 5692
rect 17368 5652 17374 5664
rect 18506 5652 18512 5664
rect 18564 5692 18570 5704
rect 19150 5692 19156 5704
rect 18564 5664 19156 5692
rect 18564 5652 18570 5664
rect 19150 5652 19156 5664
rect 19208 5652 19214 5704
rect 17034 5584 17040 5636
rect 17092 5624 17098 5636
rect 18693 5627 18751 5633
rect 18693 5624 18705 5627
rect 17092 5596 18705 5624
rect 17092 5584 17098 5596
rect 18693 5593 18705 5596
rect 18739 5593 18751 5627
rect 18693 5587 18751 5593
rect 11664 5528 13814 5556
rect 14093 5559 14151 5565
rect 11664 5516 11670 5528
rect 14093 5525 14105 5559
rect 14139 5556 14151 5559
rect 14274 5556 14280 5568
rect 14139 5528 14280 5556
rect 14139 5525 14151 5528
rect 14093 5519 14151 5525
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 14642 5556 14648 5568
rect 14603 5528 14648 5556
rect 14642 5516 14648 5528
rect 14700 5516 14706 5568
rect 15470 5556 15476 5568
rect 15431 5528 15476 5556
rect 15470 5516 15476 5528
rect 15528 5516 15534 5568
rect 17862 5556 17868 5568
rect 17823 5528 17868 5556
rect 17862 5516 17868 5528
rect 17920 5516 17926 5568
rect 18708 5556 18736 5587
rect 18782 5584 18788 5636
rect 18840 5624 18846 5636
rect 19260 5624 19288 5732
rect 19518 5720 19524 5732
rect 19576 5760 19582 5772
rect 19904 5769 19932 5800
rect 20622 5788 20628 5840
rect 20680 5828 20686 5840
rect 21453 5831 21511 5837
rect 21453 5828 21465 5831
rect 20680 5800 21465 5828
rect 20680 5788 20686 5800
rect 21453 5797 21465 5800
rect 21499 5797 21511 5831
rect 21453 5791 21511 5797
rect 23477 5831 23535 5837
rect 23477 5797 23489 5831
rect 23523 5828 23535 5831
rect 23658 5828 23664 5840
rect 23523 5800 23664 5828
rect 23523 5797 23535 5800
rect 23477 5791 23535 5797
rect 23658 5788 23664 5800
rect 23716 5788 23722 5840
rect 25038 5828 25044 5840
rect 24999 5800 25044 5828
rect 25038 5788 25044 5800
rect 25096 5788 25102 5840
rect 19705 5763 19763 5769
rect 19705 5760 19717 5763
rect 19576 5732 19717 5760
rect 19576 5720 19582 5732
rect 19705 5729 19717 5732
rect 19751 5729 19763 5763
rect 19705 5723 19763 5729
rect 19889 5763 19947 5769
rect 19889 5729 19901 5763
rect 19935 5760 19947 5763
rect 20070 5760 20076 5772
rect 19935 5732 20076 5760
rect 19935 5729 19947 5732
rect 19889 5723 19947 5729
rect 20070 5720 20076 5732
rect 20128 5720 20134 5772
rect 21266 5720 21272 5772
rect 21324 5760 21330 5772
rect 21545 5763 21603 5769
rect 21545 5760 21557 5763
rect 21324 5732 21557 5760
rect 21324 5720 21330 5732
rect 21545 5729 21557 5732
rect 21591 5729 21603 5763
rect 21545 5723 21603 5729
rect 23382 5692 23388 5704
rect 23343 5664 23388 5692
rect 23382 5652 23388 5664
rect 23440 5652 23446 5704
rect 23566 5652 23572 5704
rect 23624 5692 23630 5704
rect 23661 5695 23719 5701
rect 23661 5692 23673 5695
rect 23624 5664 23673 5692
rect 23624 5652 23630 5664
rect 23661 5661 23673 5664
rect 23707 5661 23719 5695
rect 24946 5692 24952 5704
rect 24907 5664 24952 5692
rect 23661 5655 23719 5661
rect 24946 5652 24952 5664
rect 25004 5652 25010 5704
rect 25225 5695 25283 5701
rect 25225 5661 25237 5695
rect 25271 5661 25283 5695
rect 25225 5655 25283 5661
rect 18840 5596 19288 5624
rect 18840 5584 18846 5596
rect 20254 5584 20260 5636
rect 20312 5624 20318 5636
rect 22738 5624 22744 5636
rect 20312 5596 22744 5624
rect 20312 5584 20318 5596
rect 22738 5584 22744 5596
rect 22796 5624 22802 5636
rect 22796 5596 23474 5624
rect 22796 5584 22802 5596
rect 19150 5556 19156 5568
rect 18708 5528 19156 5556
rect 19150 5516 19156 5528
rect 19208 5516 19214 5568
rect 19978 5516 19984 5568
rect 20036 5556 20042 5568
rect 23446 5556 23474 5596
rect 25240 5556 25268 5655
rect 20036 5528 20081 5556
rect 23446 5528 25268 5556
rect 20036 5516 20042 5528
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 5859 5355 5917 5361
rect 5859 5321 5871 5355
rect 5905 5352 5917 5355
rect 5994 5352 6000 5364
rect 5905 5324 6000 5352
rect 5905 5321 5917 5324
rect 5859 5315 5917 5321
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 6638 5352 6644 5364
rect 6551 5324 6644 5352
rect 6638 5312 6644 5324
rect 6696 5352 6702 5364
rect 7006 5352 7012 5364
rect 6696 5324 7012 5352
rect 6696 5312 6702 5324
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 7101 5355 7159 5361
rect 7101 5321 7113 5355
rect 7147 5352 7159 5355
rect 7282 5352 7288 5364
rect 7147 5324 7288 5352
rect 7147 5321 7159 5324
rect 7101 5315 7159 5321
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 7466 5352 7472 5364
rect 7427 5324 7472 5352
rect 7466 5312 7472 5324
rect 7524 5312 7530 5364
rect 8386 5352 8392 5364
rect 8347 5324 8392 5352
rect 8386 5312 8392 5324
rect 8444 5312 8450 5364
rect 10686 5312 10692 5364
rect 10744 5352 10750 5364
rect 11241 5355 11299 5361
rect 11241 5352 11253 5355
rect 10744 5324 11253 5352
rect 10744 5312 10750 5324
rect 11241 5321 11253 5324
rect 11287 5352 11299 5355
rect 11514 5352 11520 5364
rect 11287 5324 11520 5352
rect 11287 5321 11299 5324
rect 11241 5315 11299 5321
rect 11514 5312 11520 5324
rect 11572 5312 11578 5364
rect 12158 5352 12164 5364
rect 12119 5324 12164 5352
rect 12158 5312 12164 5324
rect 12216 5352 12222 5364
rect 12802 5352 12808 5364
rect 12216 5324 12808 5352
rect 12216 5312 12222 5324
rect 12802 5312 12808 5324
rect 12860 5312 12866 5364
rect 14553 5355 14611 5361
rect 14553 5321 14565 5355
rect 14599 5352 14611 5355
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 14599 5324 14933 5352
rect 14599 5321 14611 5324
rect 14553 5315 14611 5321
rect 14921 5321 14933 5324
rect 14967 5352 14979 5355
rect 15378 5352 15384 5364
rect 14967 5324 15384 5352
rect 14967 5321 14979 5324
rect 14921 5315 14979 5321
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 15654 5352 15660 5364
rect 15615 5324 15660 5352
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 16114 5312 16120 5364
rect 16172 5352 16178 5364
rect 16301 5355 16359 5361
rect 16301 5352 16313 5355
rect 16172 5324 16313 5352
rect 16172 5312 16178 5324
rect 16301 5321 16313 5324
rect 16347 5321 16359 5355
rect 17310 5352 17316 5364
rect 17271 5324 17316 5352
rect 16301 5315 16359 5321
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 18322 5312 18328 5364
rect 18380 5352 18386 5364
rect 18509 5355 18567 5361
rect 18509 5352 18521 5355
rect 18380 5324 18521 5352
rect 18380 5312 18386 5324
rect 18509 5321 18521 5324
rect 18555 5352 18567 5355
rect 18877 5355 18935 5361
rect 18877 5352 18889 5355
rect 18555 5324 18889 5352
rect 18555 5321 18567 5324
rect 18509 5315 18567 5321
rect 18877 5321 18889 5324
rect 18923 5321 18935 5355
rect 21266 5352 21272 5364
rect 21227 5324 21272 5352
rect 18877 5315 18935 5321
rect 10042 5284 10048 5296
rect 9955 5256 10048 5284
rect 10042 5244 10048 5256
rect 10100 5284 10106 5296
rect 10778 5284 10784 5296
rect 10100 5256 10784 5284
rect 10100 5244 10106 5256
rect 10778 5244 10784 5256
rect 10836 5244 10842 5296
rect 11146 5244 11152 5296
rect 11204 5284 11210 5296
rect 11609 5287 11667 5293
rect 11609 5284 11621 5287
rect 11204 5256 11621 5284
rect 11204 5244 11210 5256
rect 11609 5253 11621 5256
rect 11655 5253 11667 5287
rect 11609 5247 11667 5253
rect 14642 5244 14648 5296
rect 14700 5284 14706 5296
rect 14700 5256 15056 5284
rect 14700 5244 14706 5256
rect 8110 5176 8116 5228
rect 8168 5216 8174 5228
rect 9950 5216 9956 5228
rect 8168 5188 9956 5216
rect 8168 5176 8174 5188
rect 9950 5176 9956 5188
rect 10008 5216 10014 5228
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 10008 5188 10241 5216
rect 10008 5176 10014 5188
rect 10229 5185 10241 5188
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5216 10931 5219
rect 11238 5216 11244 5228
rect 10919 5188 11244 5216
rect 10919 5185 10931 5188
rect 10873 5179 10931 5185
rect 11238 5176 11244 5188
rect 11296 5176 11302 5228
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5216 13047 5219
rect 13035 5188 13584 5216
rect 13035 5185 13047 5188
rect 12989 5179 13047 5185
rect 7650 5157 7656 5160
rect 4776 5151 4834 5157
rect 4776 5117 4788 5151
rect 4822 5148 4834 5151
rect 5788 5151 5846 5157
rect 4822 5120 5304 5148
rect 4822 5117 4834 5120
rect 4776 5111 4834 5117
rect 4847 5015 4905 5021
rect 4847 4981 4859 5015
rect 4893 5012 4905 5015
rect 4982 5012 4988 5024
rect 4893 4984 4988 5012
rect 4893 4981 4905 4984
rect 4847 4975 4905 4981
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 5276 5021 5304 5120
rect 5788 5117 5800 5151
rect 5834 5148 5846 5151
rect 7628 5151 7656 5157
rect 7628 5148 7640 5151
rect 5834 5120 6316 5148
rect 7563 5120 7640 5148
rect 5834 5117 5846 5120
rect 5788 5111 5846 5117
rect 6288 5024 6316 5120
rect 7628 5117 7640 5120
rect 7708 5148 7714 5160
rect 8018 5148 8024 5160
rect 7708 5120 8024 5148
rect 7628 5111 7656 5117
rect 7650 5108 7656 5111
rect 7708 5108 7714 5120
rect 8018 5108 8024 5120
rect 8076 5108 8082 5160
rect 8846 5148 8852 5160
rect 8807 5120 8852 5148
rect 8846 5108 8852 5120
rect 8904 5108 8910 5160
rect 9125 5151 9183 5157
rect 9125 5117 9137 5151
rect 9171 5148 9183 5151
rect 9674 5148 9680 5160
rect 9171 5120 9680 5148
rect 9171 5117 9183 5120
rect 9125 5111 9183 5117
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 13170 5148 13176 5160
rect 13131 5120 13176 5148
rect 13170 5108 13176 5120
rect 13228 5108 13234 5160
rect 13556 5157 13584 5188
rect 14182 5176 14188 5228
rect 14240 5216 14246 5228
rect 14734 5216 14740 5228
rect 14240 5188 14740 5216
rect 14240 5176 14246 5188
rect 14734 5176 14740 5188
rect 14792 5225 14798 5228
rect 15028 5225 15056 5256
rect 14792 5219 14850 5225
rect 14792 5185 14804 5219
rect 14838 5185 14850 5219
rect 14792 5179 14850 5185
rect 15013 5219 15071 5225
rect 15013 5185 15025 5219
rect 15059 5216 15071 5219
rect 15562 5216 15568 5228
rect 15059 5188 15568 5216
rect 15059 5185 15071 5188
rect 15013 5179 15071 5185
rect 14792 5176 14798 5179
rect 15562 5176 15568 5188
rect 15620 5176 15626 5228
rect 16022 5176 16028 5228
rect 16080 5216 16086 5228
rect 16080 5188 16804 5216
rect 16080 5176 16086 5188
rect 13541 5151 13599 5157
rect 13541 5117 13553 5151
rect 13587 5148 13599 5151
rect 13587 5120 14596 5148
rect 13587 5117 13599 5120
rect 13541 5111 13599 5117
rect 9309 5083 9367 5089
rect 9309 5049 9321 5083
rect 9355 5080 9367 5083
rect 9398 5080 9404 5092
rect 9355 5052 9404 5080
rect 9355 5049 9367 5052
rect 9309 5043 9367 5049
rect 9398 5040 9404 5052
rect 9456 5040 9462 5092
rect 10321 5083 10379 5089
rect 9876 5052 10180 5080
rect 9876 5024 9904 5052
rect 5261 5015 5319 5021
rect 5261 4981 5273 5015
rect 5307 5012 5319 5015
rect 5350 5012 5356 5024
rect 5307 4984 5356 5012
rect 5307 4981 5319 4984
rect 5261 4975 5319 4981
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 6270 5012 6276 5024
rect 6231 4984 6276 5012
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 7699 5015 7757 5021
rect 7699 4981 7711 5015
rect 7745 5012 7757 5015
rect 7834 5012 7840 5024
rect 7745 4984 7840 5012
rect 7745 4981 7757 4984
rect 7699 4975 7757 4981
rect 7834 4972 7840 4984
rect 7892 4972 7898 5024
rect 8113 5015 8171 5021
rect 8113 4981 8125 5015
rect 8159 5012 8171 5015
rect 8202 5012 8208 5024
rect 8159 4984 8208 5012
rect 8159 4981 8171 4984
rect 8113 4975 8171 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 9677 5015 9735 5021
rect 9677 4981 9689 5015
rect 9723 5012 9735 5015
rect 9858 5012 9864 5024
rect 9723 4984 9864 5012
rect 9723 4981 9735 4984
rect 9677 4975 9735 4981
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 10152 5012 10180 5052
rect 10321 5049 10333 5083
rect 10367 5049 10379 5083
rect 10321 5043 10379 5049
rect 10336 5012 10364 5043
rect 10962 5040 10968 5092
rect 11020 5080 11026 5092
rect 11020 5052 12934 5080
rect 11020 5040 11026 5052
rect 10152 4984 10364 5012
rect 12906 5012 12934 5052
rect 14568 5024 14596 5120
rect 15654 5108 15660 5160
rect 15712 5148 15718 5160
rect 16776 5157 16804 5188
rect 16209 5151 16267 5157
rect 16209 5148 16221 5151
rect 15712 5120 16221 5148
rect 15712 5108 15718 5120
rect 16209 5117 16221 5120
rect 16255 5117 16267 5151
rect 16209 5111 16267 5117
rect 16761 5151 16819 5157
rect 16761 5117 16773 5151
rect 16807 5148 16819 5151
rect 17678 5148 17684 5160
rect 16807 5120 17684 5148
rect 16807 5117 16819 5120
rect 16761 5111 16819 5117
rect 17678 5108 17684 5120
rect 17736 5108 17742 5160
rect 18892 5148 18920 5315
rect 21266 5312 21272 5324
rect 21324 5312 21330 5364
rect 21450 5312 21456 5364
rect 21508 5352 21514 5364
rect 21545 5355 21603 5361
rect 21545 5352 21557 5355
rect 21508 5324 21557 5352
rect 21508 5312 21514 5324
rect 21545 5321 21557 5324
rect 21591 5321 21603 5355
rect 21545 5315 21603 5321
rect 23109 5355 23167 5361
rect 23109 5321 23121 5355
rect 23155 5352 23167 5355
rect 23658 5352 23664 5364
rect 23155 5324 23664 5352
rect 23155 5321 23167 5324
rect 23109 5315 23167 5321
rect 23658 5312 23664 5324
rect 23716 5312 23722 5364
rect 24949 5355 25007 5361
rect 24949 5321 24961 5355
rect 24995 5352 25007 5355
rect 25038 5352 25044 5364
rect 24995 5324 25044 5352
rect 24995 5321 25007 5324
rect 24949 5315 25007 5321
rect 25038 5312 25044 5324
rect 25096 5312 25102 5364
rect 19978 5176 19984 5228
rect 20036 5216 20042 5228
rect 21726 5216 21732 5228
rect 20036 5188 21732 5216
rect 20036 5176 20042 5188
rect 21726 5176 21732 5188
rect 21784 5176 21790 5228
rect 19061 5151 19119 5157
rect 19061 5148 19073 5151
rect 18892 5120 19073 5148
rect 19061 5117 19073 5120
rect 19107 5117 19119 5151
rect 19061 5111 19119 5117
rect 19150 5108 19156 5160
rect 19208 5148 19214 5160
rect 19889 5151 19947 5157
rect 19889 5148 19901 5151
rect 19208 5120 19901 5148
rect 19208 5108 19214 5120
rect 19889 5117 19901 5120
rect 19935 5117 19947 5151
rect 20070 5148 20076 5160
rect 19983 5120 20076 5148
rect 19889 5111 19947 5117
rect 14642 5040 14648 5092
rect 14700 5080 14706 5092
rect 15838 5080 15844 5092
rect 14700 5052 15844 5080
rect 14700 5040 14706 5052
rect 15838 5040 15844 5052
rect 15896 5080 15902 5092
rect 19904 5080 19932 5111
rect 20070 5108 20076 5120
rect 20128 5148 20134 5160
rect 20809 5151 20867 5157
rect 20809 5148 20821 5151
rect 20128 5120 20821 5148
rect 20128 5108 20134 5120
rect 20809 5117 20821 5120
rect 20855 5117 20867 5151
rect 20809 5111 20867 5117
rect 25130 5108 25136 5160
rect 25188 5148 25194 5160
rect 25225 5151 25283 5157
rect 25225 5148 25237 5151
rect 25188 5120 25237 5148
rect 25188 5108 25194 5120
rect 25225 5117 25237 5120
rect 25271 5148 25283 5151
rect 25777 5151 25835 5157
rect 25777 5148 25789 5151
rect 25271 5120 25789 5148
rect 25271 5117 25283 5120
rect 25225 5111 25283 5117
rect 25777 5117 25789 5120
rect 25823 5117 25835 5151
rect 25777 5111 25835 5117
rect 20441 5083 20499 5089
rect 20441 5080 20453 5083
rect 15896 5052 19012 5080
rect 19904 5052 20453 5080
rect 15896 5040 15902 5052
rect 13173 5015 13231 5021
rect 13173 5012 13185 5015
rect 12906 4984 13185 5012
rect 13173 4981 13185 4984
rect 13219 4981 13231 5015
rect 14182 5012 14188 5024
rect 14143 4984 14188 5012
rect 13173 4975 13231 4981
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 14550 4972 14556 5024
rect 14608 5012 14614 5024
rect 15289 5015 15347 5021
rect 15289 5012 15301 5015
rect 14608 4984 15301 5012
rect 14608 4972 14614 4984
rect 15289 4981 15301 4984
rect 15335 4981 15347 5015
rect 16022 5012 16028 5024
rect 15983 4984 16028 5012
rect 15289 4975 15347 4981
rect 16022 4972 16028 4984
rect 16080 4972 16086 5024
rect 18049 5015 18107 5021
rect 18049 4981 18061 5015
rect 18095 5012 18107 5015
rect 18138 5012 18144 5024
rect 18095 4984 18144 5012
rect 18095 4981 18107 4984
rect 18049 4975 18107 4981
rect 18138 4972 18144 4984
rect 18196 4972 18202 5024
rect 18984 5012 19012 5052
rect 20441 5049 20453 5052
rect 20487 5049 20499 5083
rect 20441 5043 20499 5049
rect 21450 5040 21456 5092
rect 21508 5080 21514 5092
rect 22050 5083 22108 5089
rect 22050 5080 22062 5083
rect 21508 5052 22062 5080
rect 21508 5040 21514 5052
rect 22050 5049 22062 5052
rect 22096 5049 22108 5083
rect 23750 5080 23756 5092
rect 23711 5052 23756 5080
rect 22050 5043 22108 5049
rect 23750 5040 23756 5052
rect 23808 5040 23814 5092
rect 23845 5083 23903 5089
rect 23845 5049 23857 5083
rect 23891 5049 23903 5083
rect 23845 5043 23903 5049
rect 24397 5083 24455 5089
rect 24397 5049 24409 5083
rect 24443 5080 24455 5083
rect 24946 5080 24952 5092
rect 24443 5052 24952 5080
rect 24443 5049 24455 5052
rect 24397 5043 24455 5049
rect 19058 5012 19064 5024
rect 18984 4984 19064 5012
rect 19058 4972 19064 4984
rect 19116 4972 19122 5024
rect 20162 5012 20168 5024
rect 20123 4984 20168 5012
rect 20162 4972 20168 4984
rect 20220 4972 20226 5024
rect 22646 5012 22652 5024
rect 22607 4984 22652 5012
rect 22646 4972 22652 4984
rect 22704 4972 22710 5024
rect 23477 5015 23535 5021
rect 23477 4981 23489 5015
rect 23523 5012 23535 5015
rect 23566 5012 23572 5024
rect 23523 4984 23572 5012
rect 23523 4981 23535 4984
rect 23477 4975 23535 4981
rect 23566 4972 23572 4984
rect 23624 5012 23630 5024
rect 23860 5012 23888 5043
rect 24946 5040 24952 5052
rect 25004 5040 25010 5092
rect 23624 4984 23888 5012
rect 25409 5015 25467 5021
rect 23624 4972 23630 4984
rect 25409 4981 25421 5015
rect 25455 5012 25467 5015
rect 25682 5012 25688 5024
rect 25455 4984 25688 5012
rect 25455 4981 25467 4984
rect 25409 4975 25467 4981
rect 25682 4972 25688 4984
rect 25740 4972 25746 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 4755 4811 4813 4817
rect 4755 4777 4767 4811
rect 4801 4808 4813 4811
rect 5074 4808 5080 4820
rect 4801 4780 5080 4808
rect 4801 4777 4813 4780
rect 4755 4771 4813 4777
rect 5074 4768 5080 4780
rect 5132 4768 5138 4820
rect 5767 4811 5825 4817
rect 5767 4777 5779 4811
rect 5813 4808 5825 4811
rect 6086 4808 6092 4820
rect 5813 4780 6092 4808
rect 5813 4777 5825 4780
rect 5767 4771 5825 4777
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 7929 4811 7987 4817
rect 7929 4777 7941 4811
rect 7975 4808 7987 4811
rect 8478 4808 8484 4820
rect 7975 4780 8484 4808
rect 7975 4777 7987 4780
rect 7929 4771 7987 4777
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 8846 4768 8852 4820
rect 8904 4808 8910 4820
rect 9033 4811 9091 4817
rect 9033 4808 9045 4811
rect 8904 4780 9045 4808
rect 8904 4768 8910 4780
rect 9033 4777 9045 4780
rect 9079 4808 9091 4811
rect 9309 4811 9367 4817
rect 9309 4808 9321 4811
rect 9079 4780 9321 4808
rect 9079 4777 9091 4780
rect 9033 4771 9091 4777
rect 9309 4777 9321 4780
rect 9355 4777 9367 4811
rect 9309 4771 9367 4777
rect 9493 4811 9551 4817
rect 9493 4777 9505 4811
rect 9539 4808 9551 4811
rect 9674 4808 9680 4820
rect 9539 4780 9680 4808
rect 9539 4777 9551 4780
rect 9493 4771 9551 4777
rect 4684 4675 4742 4681
rect 4684 4641 4696 4675
rect 4730 4672 4742 4675
rect 5166 4672 5172 4684
rect 4730 4644 5172 4672
rect 4730 4641 4742 4644
rect 4684 4635 4742 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5696 4675 5754 4681
rect 5696 4641 5708 4675
rect 5742 4672 5754 4675
rect 6178 4672 6184 4684
rect 5742 4644 6184 4672
rect 5742 4641 5754 4644
rect 5696 4635 5754 4641
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 7076 4675 7134 4681
rect 7076 4641 7088 4675
rect 7122 4672 7134 4675
rect 7282 4672 7288 4684
rect 7122 4644 7288 4672
rect 7122 4641 7134 4644
rect 7076 4635 7134 4641
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 8294 4672 8300 4684
rect 8255 4644 8300 4672
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 8478 4632 8484 4684
rect 8536 4672 8542 4684
rect 8573 4675 8631 4681
rect 8573 4672 8585 4675
rect 8536 4644 8585 4672
rect 8536 4632 8542 4644
rect 8573 4641 8585 4644
rect 8619 4672 8631 4675
rect 9508 4672 9536 4771
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 9950 4768 9956 4820
rect 10008 4808 10014 4820
rect 10873 4811 10931 4817
rect 10873 4808 10885 4811
rect 10008 4780 10885 4808
rect 10008 4768 10014 4780
rect 10873 4777 10885 4780
rect 10919 4777 10931 4811
rect 10873 4771 10931 4777
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 13449 4811 13507 4817
rect 13449 4808 13461 4811
rect 12768 4780 13461 4808
rect 12768 4768 12774 4780
rect 13449 4777 13461 4780
rect 13495 4777 13507 4811
rect 13725 4811 13783 4817
rect 13725 4808 13737 4811
rect 13449 4771 13507 4777
rect 13556 4780 13737 4808
rect 9858 4740 9864 4752
rect 9819 4712 9864 4740
rect 9858 4700 9864 4712
rect 9916 4700 9922 4752
rect 11054 4700 11060 4752
rect 11112 4740 11118 4752
rect 11609 4743 11667 4749
rect 11609 4740 11621 4743
rect 11112 4712 11621 4740
rect 11112 4700 11118 4712
rect 11609 4709 11621 4712
rect 11655 4740 11667 4743
rect 11790 4740 11796 4752
rect 11655 4712 11796 4740
rect 11655 4709 11667 4712
rect 11609 4703 11667 4709
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 12618 4700 12624 4752
rect 12676 4740 12682 4752
rect 13556 4740 13584 4780
rect 13725 4777 13737 4780
rect 13771 4777 13783 4811
rect 14642 4808 14648 4820
rect 14603 4780 14648 4808
rect 13725 4771 13783 4777
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 16669 4811 16727 4817
rect 16669 4808 16681 4811
rect 15344 4780 16681 4808
rect 15344 4768 15350 4780
rect 16669 4777 16681 4780
rect 16715 4777 16727 4811
rect 16669 4771 16727 4777
rect 18414 4768 18420 4820
rect 18472 4808 18478 4820
rect 18509 4811 18567 4817
rect 18509 4808 18521 4811
rect 18472 4780 18521 4808
rect 18472 4768 18478 4780
rect 18509 4777 18521 4780
rect 18555 4777 18567 4811
rect 18509 4771 18567 4777
rect 18690 4768 18696 4820
rect 18748 4808 18754 4820
rect 18877 4811 18935 4817
rect 18877 4808 18889 4811
rect 18748 4780 18889 4808
rect 18748 4768 18754 4780
rect 18877 4777 18889 4780
rect 18923 4777 18935 4811
rect 21726 4808 21732 4820
rect 21687 4780 21732 4808
rect 18877 4771 18935 4777
rect 21726 4768 21732 4780
rect 21784 4768 21790 4820
rect 23382 4808 23388 4820
rect 23343 4780 23388 4808
rect 23382 4768 23388 4780
rect 23440 4768 23446 4820
rect 23750 4808 23756 4820
rect 23711 4780 23756 4808
rect 23750 4768 23756 4780
rect 23808 4768 23814 4820
rect 24946 4808 24952 4820
rect 24688 4780 24952 4808
rect 12676 4712 13584 4740
rect 12676 4700 12682 4712
rect 14366 4700 14372 4752
rect 14424 4740 14430 4752
rect 14424 4712 15332 4740
rect 14424 4700 14430 4712
rect 15304 4684 15332 4712
rect 18966 4700 18972 4752
rect 19024 4740 19030 4752
rect 19245 4743 19303 4749
rect 19245 4740 19257 4743
rect 19024 4712 19257 4740
rect 19024 4700 19030 4712
rect 19245 4709 19257 4712
rect 19291 4709 19303 4743
rect 19245 4703 19303 4709
rect 21450 4700 21456 4752
rect 21508 4740 21514 4752
rect 22326 4743 22384 4749
rect 22326 4740 22338 4743
rect 21508 4712 22338 4740
rect 21508 4700 21514 4712
rect 22326 4709 22338 4712
rect 22372 4709 22384 4743
rect 24118 4740 24124 4752
rect 24079 4712 24124 4740
rect 22326 4703 22384 4709
rect 24118 4700 24124 4712
rect 24176 4700 24182 4752
rect 24688 4749 24716 4780
rect 24946 4768 24952 4780
rect 25004 4768 25010 4820
rect 24673 4743 24731 4749
rect 24673 4709 24685 4743
rect 24719 4709 24731 4743
rect 24673 4703 24731 4709
rect 8619 4644 9536 4672
rect 10505 4675 10563 4681
rect 8619 4641 8631 4644
rect 8573 4635 8631 4641
rect 10505 4641 10517 4675
rect 10551 4672 10563 4675
rect 10686 4672 10692 4684
rect 10551 4644 10692 4672
rect 10551 4641 10563 4644
rect 10505 4635 10563 4641
rect 10686 4632 10692 4644
rect 10744 4632 10750 4684
rect 13446 4632 13452 4684
rect 13504 4672 13510 4684
rect 13633 4675 13691 4681
rect 13633 4672 13645 4675
rect 13504 4644 13645 4672
rect 13504 4632 13510 4644
rect 13633 4641 13645 4644
rect 13679 4641 13691 4675
rect 13633 4635 13691 4641
rect 8754 4604 8760 4616
rect 8715 4576 8760 4604
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 11517 4607 11575 4613
rect 11517 4573 11529 4607
rect 11563 4604 11575 4607
rect 11606 4604 11612 4616
rect 11563 4576 11612 4604
rect 11563 4573 11575 4576
rect 11517 4567 11575 4573
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4604 11851 4607
rect 12434 4604 12440 4616
rect 11839 4576 12440 4604
rect 11839 4573 11851 4576
rect 11793 4567 11851 4573
rect 8570 4496 8576 4548
rect 8628 4536 8634 4548
rect 11808 4536 11836 4567
rect 12434 4564 12440 4576
rect 12492 4564 12498 4616
rect 12526 4564 12532 4616
rect 12584 4604 12590 4616
rect 13081 4607 13139 4613
rect 13081 4604 13093 4607
rect 12584 4576 13093 4604
rect 12584 4564 12590 4576
rect 13081 4573 13093 4576
rect 13127 4604 13139 4607
rect 13170 4604 13176 4616
rect 13127 4576 13176 4604
rect 13127 4573 13139 4576
rect 13081 4567 13139 4573
rect 13170 4564 13176 4576
rect 13228 4564 13234 4616
rect 13648 4604 13676 4635
rect 13998 4632 14004 4684
rect 14056 4672 14062 4684
rect 14185 4675 14243 4681
rect 14185 4672 14197 4675
rect 14056 4644 14197 4672
rect 14056 4632 14062 4644
rect 14185 4641 14197 4644
rect 14231 4672 14243 4675
rect 14550 4672 14556 4684
rect 14231 4644 14556 4672
rect 14231 4641 14243 4644
rect 14185 4635 14243 4641
rect 14550 4632 14556 4644
rect 14608 4632 14614 4684
rect 15286 4672 15292 4684
rect 15199 4644 15292 4672
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 15378 4632 15384 4684
rect 15436 4672 15442 4684
rect 15519 4675 15577 4681
rect 15519 4672 15531 4675
rect 15436 4644 15531 4672
rect 15436 4632 15442 4644
rect 15519 4641 15531 4644
rect 15565 4672 15577 4675
rect 16114 4672 16120 4684
rect 15565 4644 16120 4672
rect 15565 4641 15577 4644
rect 15519 4635 15577 4641
rect 16114 4632 16120 4644
rect 16172 4632 16178 4684
rect 17126 4632 17132 4684
rect 17184 4672 17190 4684
rect 17497 4675 17555 4681
rect 17497 4672 17509 4675
rect 17184 4644 17509 4672
rect 17184 4632 17190 4644
rect 17497 4641 17509 4644
rect 17543 4641 17555 4675
rect 17497 4635 17555 4641
rect 20622 4632 20628 4684
rect 20680 4672 20686 4684
rect 20901 4675 20959 4681
rect 20901 4672 20913 4675
rect 20680 4644 20913 4672
rect 20680 4632 20686 4644
rect 20901 4641 20913 4644
rect 20947 4641 20959 4675
rect 20901 4635 20959 4641
rect 14642 4604 14648 4616
rect 13648 4576 14648 4604
rect 14642 4564 14648 4576
rect 14700 4564 14706 4616
rect 15654 4604 15660 4616
rect 15615 4576 15660 4604
rect 15654 4564 15660 4576
rect 15712 4564 15718 4616
rect 17773 4607 17831 4613
rect 17773 4573 17785 4607
rect 17819 4604 17831 4607
rect 18046 4604 18052 4616
rect 17819 4576 18052 4604
rect 17819 4573 17831 4576
rect 17773 4567 17831 4573
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 19150 4604 19156 4616
rect 19111 4576 19156 4604
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 15105 4539 15163 4545
rect 15105 4536 15117 4539
rect 8628 4508 11836 4536
rect 12728 4508 15117 4536
rect 8628 4496 8634 4508
rect 12728 4480 12756 4508
rect 15105 4505 15117 4508
rect 15151 4536 15163 4539
rect 15151 4508 15976 4536
rect 15151 4505 15163 4508
rect 15105 4499 15163 4505
rect 7147 4471 7205 4477
rect 7147 4437 7159 4471
rect 7193 4468 7205 4471
rect 7650 4468 7656 4480
rect 7193 4440 7656 4468
rect 7193 4437 7205 4440
rect 7147 4431 7205 4437
rect 7650 4428 7656 4440
rect 7708 4428 7714 4480
rect 9309 4471 9367 4477
rect 9309 4437 9321 4471
rect 9355 4468 9367 4471
rect 12434 4468 12440 4480
rect 9355 4440 12440 4468
rect 9355 4437 9367 4440
rect 9309 4431 9367 4437
rect 12434 4428 12440 4440
rect 12492 4428 12498 4480
rect 12710 4468 12716 4480
rect 12671 4440 12716 4468
rect 12710 4428 12716 4440
rect 12768 4428 12774 4480
rect 14734 4428 14740 4480
rect 14792 4468 14798 4480
rect 15948 4477 15976 4508
rect 16022 4496 16028 4548
rect 16080 4536 16086 4548
rect 16301 4539 16359 4545
rect 16301 4536 16313 4539
rect 16080 4508 16313 4536
rect 16080 4496 16086 4508
rect 16301 4505 16313 4508
rect 16347 4536 16359 4539
rect 16945 4539 17003 4545
rect 16945 4536 16957 4539
rect 16347 4508 16957 4536
rect 16347 4505 16359 4508
rect 16301 4499 16359 4505
rect 16945 4505 16957 4508
rect 16991 4536 17003 4539
rect 17034 4536 17040 4548
rect 16991 4508 17040 4536
rect 16991 4505 17003 4508
rect 16945 4499 17003 4505
rect 17034 4496 17040 4508
rect 17092 4496 17098 4548
rect 18230 4496 18236 4548
rect 18288 4536 18294 4548
rect 19444 4536 19472 4567
rect 20162 4564 20168 4616
rect 20220 4604 20226 4616
rect 22005 4607 22063 4613
rect 22005 4604 22017 4607
rect 20220 4576 22017 4604
rect 20220 4564 20226 4576
rect 22005 4573 22017 4576
rect 22051 4604 22063 4607
rect 22186 4604 22192 4616
rect 22051 4576 22192 4604
rect 22051 4573 22063 4576
rect 22005 4567 22063 4573
rect 22186 4564 22192 4576
rect 22244 4564 22250 4616
rect 22462 4564 22468 4616
rect 22520 4604 22526 4616
rect 23014 4604 23020 4616
rect 22520 4576 23020 4604
rect 22520 4564 22526 4576
rect 23014 4564 23020 4576
rect 23072 4604 23078 4616
rect 24029 4607 24087 4613
rect 24029 4604 24041 4607
rect 23072 4576 24041 4604
rect 23072 4564 23078 4576
rect 24029 4573 24041 4576
rect 24075 4573 24087 4607
rect 24029 4567 24087 4573
rect 21085 4539 21143 4545
rect 18288 4508 21036 4536
rect 18288 4496 18294 4508
rect 15427 4471 15485 4477
rect 15427 4468 15439 4471
rect 14792 4440 15439 4468
rect 14792 4428 14798 4440
rect 15427 4437 15439 4440
rect 15473 4437 15485 4471
rect 15427 4431 15485 4437
rect 15933 4471 15991 4477
rect 15933 4437 15945 4471
rect 15979 4468 15991 4471
rect 16206 4468 16212 4480
rect 15979 4440 16212 4468
rect 15979 4437 15991 4440
rect 15933 4431 15991 4437
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 17494 4428 17500 4480
rect 17552 4468 17558 4480
rect 20070 4468 20076 4480
rect 17552 4440 20076 4468
rect 17552 4428 17558 4440
rect 20070 4428 20076 4440
rect 20128 4428 20134 4480
rect 21008 4468 21036 4508
rect 21085 4505 21097 4539
rect 21131 4536 21143 4539
rect 22370 4536 22376 4548
rect 21131 4508 22376 4536
rect 21131 4505 21143 4508
rect 21085 4499 21143 4505
rect 22370 4496 22376 4508
rect 22428 4496 22434 4548
rect 22925 4539 22983 4545
rect 22925 4505 22937 4539
rect 22971 4536 22983 4539
rect 25038 4536 25044 4548
rect 22971 4508 25044 4536
rect 22971 4505 22983 4508
rect 22925 4499 22983 4505
rect 25038 4496 25044 4508
rect 25096 4496 25102 4548
rect 21542 4468 21548 4480
rect 21008 4440 21548 4468
rect 21542 4428 21548 4440
rect 21600 4428 21606 4480
rect 22462 4428 22468 4480
rect 22520 4468 22526 4480
rect 23750 4468 23756 4480
rect 22520 4440 23756 4468
rect 22520 4428 22526 4440
rect 23750 4428 23756 4440
rect 23808 4428 23814 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1535 4267 1593 4273
rect 1535 4233 1547 4267
rect 1581 4264 1593 4267
rect 3973 4267 4031 4273
rect 3973 4264 3985 4267
rect 1581 4236 3985 4264
rect 1581 4233 1593 4236
rect 1535 4227 1593 4233
rect 3973 4233 3985 4236
rect 4019 4233 4031 4267
rect 3973 4227 4031 4233
rect 4154 4224 4160 4276
rect 4212 4264 4218 4276
rect 4847 4267 4905 4273
rect 4847 4264 4859 4267
rect 4212 4236 4859 4264
rect 4212 4224 4218 4236
rect 4847 4233 4859 4236
rect 4893 4233 4905 4267
rect 4847 4227 4905 4233
rect 12434 4224 12440 4276
rect 12492 4264 12498 4276
rect 13446 4264 13452 4276
rect 12492 4236 13452 4264
rect 12492 4224 12498 4236
rect 13446 4224 13452 4236
rect 13504 4264 13510 4276
rect 13633 4267 13691 4273
rect 13633 4264 13645 4267
rect 13504 4236 13645 4264
rect 13504 4224 13510 4236
rect 13633 4233 13645 4236
rect 13679 4233 13691 4267
rect 13633 4227 13691 4233
rect 15654 4224 15660 4276
rect 15712 4264 15718 4276
rect 16761 4267 16819 4273
rect 16761 4264 16773 4267
rect 15712 4236 16773 4264
rect 15712 4224 15718 4236
rect 16761 4233 16773 4236
rect 16807 4233 16819 4267
rect 16761 4227 16819 4233
rect 17034 4224 17040 4276
rect 17092 4264 17098 4276
rect 17129 4267 17187 4273
rect 17129 4264 17141 4267
rect 17092 4236 17141 4264
rect 17092 4224 17098 4236
rect 17129 4233 17141 4236
rect 17175 4233 17187 4267
rect 17770 4264 17776 4276
rect 17731 4236 17776 4264
rect 17129 4227 17187 4233
rect 17770 4224 17776 4236
rect 17828 4224 17834 4276
rect 18966 4264 18972 4276
rect 18927 4236 18972 4264
rect 18966 4224 18972 4236
rect 19024 4264 19030 4276
rect 19245 4267 19303 4273
rect 19245 4264 19257 4267
rect 19024 4236 19257 4264
rect 19024 4224 19030 4236
rect 19245 4233 19257 4236
rect 19291 4233 19303 4267
rect 19245 4227 19303 4233
rect 22186 4224 22192 4276
rect 22244 4264 22250 4276
rect 22373 4267 22431 4273
rect 22373 4264 22385 4267
rect 22244 4236 22385 4264
rect 22244 4224 22250 4236
rect 22373 4233 22385 4236
rect 22419 4233 22431 4267
rect 22373 4227 22431 4233
rect 22646 4224 22652 4276
rect 22704 4264 22710 4276
rect 23385 4267 23443 4273
rect 23385 4264 23397 4267
rect 22704 4236 23397 4264
rect 22704 4224 22710 4236
rect 23385 4233 23397 4236
rect 23431 4264 23443 4267
rect 23474 4264 23480 4276
rect 23431 4236 23480 4264
rect 23431 4233 23443 4236
rect 23385 4227 23443 4233
rect 23474 4224 23480 4236
rect 23532 4264 23538 4276
rect 24118 4264 24124 4276
rect 23532 4236 24124 4264
rect 23532 4224 23538 4236
rect 24118 4224 24124 4236
rect 24176 4224 24182 4276
rect 2958 4196 2964 4208
rect 2919 4168 2964 4196
rect 2958 4156 2964 4168
rect 3016 4156 3022 4208
rect 4065 4199 4123 4205
rect 4065 4165 4077 4199
rect 4111 4196 4123 4199
rect 8110 4196 8116 4208
rect 4111 4168 8116 4196
rect 4111 4165 4123 4168
rect 4065 4159 4123 4165
rect 8110 4156 8116 4168
rect 8168 4156 8174 4208
rect 8294 4156 8300 4208
rect 8352 4196 8358 4208
rect 8757 4199 8815 4205
rect 8757 4196 8769 4199
rect 8352 4168 8769 4196
rect 8352 4156 8358 4168
rect 8757 4165 8769 4168
rect 8803 4196 8815 4199
rect 10321 4199 10379 4205
rect 8803 4168 9628 4196
rect 8803 4165 8815 4168
rect 8757 4159 8815 4165
rect 6270 4088 6276 4140
rect 6328 4128 6334 4140
rect 7098 4128 7104 4140
rect 6328 4100 7104 4128
rect 6328 4088 6334 4100
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4128 7619 4131
rect 8478 4128 8484 4140
rect 7607 4100 8484 4128
rect 7607 4097 7619 4100
rect 7561 4091 7619 4097
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 9600 4128 9628 4168
rect 10321 4165 10333 4199
rect 10367 4196 10379 4199
rect 10686 4196 10692 4208
rect 10367 4168 10692 4196
rect 10367 4165 10379 4168
rect 10321 4159 10379 4165
rect 10686 4156 10692 4168
rect 10744 4156 10750 4208
rect 11790 4196 11796 4208
rect 11751 4168 11796 4196
rect 11790 4156 11796 4168
rect 11848 4156 11854 4208
rect 23014 4196 23020 4208
rect 22975 4168 23020 4196
rect 23014 4156 23020 4168
rect 23072 4156 23078 4208
rect 12161 4131 12219 4137
rect 12161 4128 12173 4131
rect 9600 4100 12173 4128
rect 12161 4097 12173 4100
rect 12207 4128 12219 4131
rect 12526 4128 12532 4140
rect 12207 4100 12532 4128
rect 12207 4097 12219 4100
rect 12161 4091 12219 4097
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 18046 4128 18052 4140
rect 13188 4100 17908 4128
rect 18007 4100 18052 4128
rect 1429 4060 1435 4072
rect 1390 4032 1435 4060
rect 1429 4020 1435 4032
rect 1487 4020 1493 4072
rect 2752 4063 2810 4069
rect 2752 4029 2764 4063
rect 2798 4060 2810 4063
rect 3764 4063 3822 4069
rect 2798 4032 3280 4060
rect 2798 4029 2810 4032
rect 2752 4023 2810 4029
rect 3252 3936 3280 4032
rect 3764 4029 3776 4063
rect 3810 4060 3822 4063
rect 4776 4063 4834 4069
rect 3810 4032 4292 4060
rect 3810 4029 3822 4032
rect 3764 4023 3822 4029
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 1857 3927 1915 3933
rect 1857 3924 1869 3927
rect 1452 3896 1869 3924
rect 1452 3884 1458 3896
rect 1857 3893 1869 3896
rect 1903 3893 1915 3927
rect 3234 3924 3240 3936
rect 3195 3896 3240 3924
rect 1857 3887 1915 3893
rect 3234 3884 3240 3896
rect 3292 3884 3298 3936
rect 3835 3927 3893 3933
rect 3835 3893 3847 3927
rect 3881 3924 3893 3927
rect 4154 3924 4160 3936
rect 3881 3896 4160 3924
rect 3881 3893 3893 3896
rect 3835 3887 3893 3893
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 4264 3933 4292 4032
rect 4776 4029 4788 4063
rect 4822 4060 4834 4063
rect 5788 4063 5846 4069
rect 4822 4032 5672 4060
rect 4822 4029 4834 4032
rect 4776 4023 4834 4029
rect 5644 4001 5672 4032
rect 5788 4029 5800 4063
rect 5834 4060 5846 4063
rect 6546 4060 6552 4072
rect 5834 4032 6552 4060
rect 5834 4029 5846 4032
rect 5788 4023 5846 4029
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 8110 4060 8116 4072
rect 8071 4032 8116 4060
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 9122 4060 9128 4072
rect 9035 4032 9128 4060
rect 9122 4020 9128 4032
rect 9180 4060 9186 4072
rect 9309 4063 9367 4069
rect 9309 4060 9321 4063
rect 9180 4032 9321 4060
rect 9180 4020 9186 4032
rect 9309 4029 9321 4032
rect 9355 4029 9367 4063
rect 9309 4023 9367 4029
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 10689 4063 10747 4069
rect 9456 4032 10088 4060
rect 9456 4020 9462 4032
rect 5629 3995 5687 4001
rect 5629 3961 5641 3995
rect 5675 3992 5687 3995
rect 6270 3992 6276 4004
rect 5675 3964 6276 3992
rect 5675 3961 5687 3964
rect 5629 3955 5687 3961
rect 6270 3952 6276 3964
rect 6328 3952 6334 4004
rect 9214 3952 9220 4004
rect 9272 3992 9278 4004
rect 9950 3992 9956 4004
rect 9272 3964 9956 3992
rect 9272 3952 9278 3964
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 10060 3992 10088 4032
rect 10689 4029 10701 4063
rect 10735 4060 10747 4063
rect 11330 4060 11336 4072
rect 10735 4032 11336 4060
rect 10735 4029 10747 4032
rect 10689 4023 10747 4029
rect 11330 4020 11336 4032
rect 11388 4020 11394 4072
rect 11514 4060 11520 4072
rect 11475 4032 11520 4060
rect 11514 4020 11520 4032
rect 11572 4020 11578 4072
rect 12710 4020 12716 4072
rect 12768 4060 12774 4072
rect 13081 4063 13139 4069
rect 13081 4060 13093 4063
rect 12768 4032 13093 4060
rect 12768 4020 12774 4032
rect 13081 4029 13093 4032
rect 13127 4029 13139 4063
rect 13081 4023 13139 4029
rect 13188 3992 13216 4100
rect 15749 4063 15807 4069
rect 15749 4060 15761 4063
rect 15304 4032 15761 4060
rect 13354 3992 13360 4004
rect 10060 3964 13216 3992
rect 13315 3964 13360 3992
rect 13354 3952 13360 3964
rect 13412 3952 13418 4004
rect 14274 3992 14280 4004
rect 14235 3964 14280 3992
rect 14274 3952 14280 3964
rect 14332 3952 14338 4004
rect 14369 3995 14427 4001
rect 14369 3961 14381 3995
rect 14415 3961 14427 3995
rect 14918 3992 14924 4004
rect 14879 3964 14924 3992
rect 14369 3955 14427 3961
rect 4249 3927 4307 3933
rect 4249 3893 4261 3927
rect 4295 3924 4307 3927
rect 4430 3924 4436 3936
rect 4295 3896 4436 3924
rect 4295 3893 4307 3896
rect 4249 3887 4307 3893
rect 4430 3884 4436 3896
rect 4488 3884 4494 3936
rect 5166 3924 5172 3936
rect 5127 3896 5172 3924
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 5859 3927 5917 3933
rect 5859 3893 5871 3927
rect 5905 3924 5917 3927
rect 5994 3924 6000 3936
rect 5905 3896 6000 3924
rect 5905 3893 5917 3896
rect 5859 3887 5917 3893
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 6178 3924 6184 3936
rect 6139 3896 6184 3924
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 7101 3927 7159 3933
rect 7101 3893 7113 3927
rect 7147 3924 7159 3927
rect 7282 3924 7288 3936
rect 7147 3896 7288 3924
rect 7147 3893 7159 3896
rect 7101 3887 7159 3893
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 8481 3927 8539 3933
rect 8481 3893 8493 3927
rect 8527 3924 8539 3927
rect 9582 3924 9588 3936
rect 8527 3896 9588 3924
rect 8527 3893 8539 3896
rect 8481 3887 8539 3893
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 9677 3927 9735 3933
rect 9677 3893 9689 3927
rect 9723 3924 9735 3927
rect 9858 3924 9864 3936
rect 9723 3896 9864 3924
rect 9723 3893 9735 3896
rect 9677 3887 9735 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 13906 3884 13912 3936
rect 13964 3924 13970 3936
rect 14001 3927 14059 3933
rect 14001 3924 14013 3927
rect 13964 3896 14013 3924
rect 13964 3884 13970 3896
rect 14001 3893 14013 3896
rect 14047 3924 14059 3927
rect 14384 3924 14412 3955
rect 14918 3952 14924 3964
rect 14976 3952 14982 4004
rect 14047 3896 14412 3924
rect 14047 3893 14059 3896
rect 14001 3887 14059 3893
rect 14642 3884 14648 3936
rect 14700 3924 14706 3936
rect 15304 3924 15332 4032
rect 15749 4029 15761 4032
rect 15795 4060 15807 4063
rect 16022 4060 16028 4072
rect 15795 4032 16028 4060
rect 15795 4029 15807 4032
rect 15749 4023 15807 4029
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 16206 4060 16212 4072
rect 16167 4032 16212 4060
rect 16206 4020 16212 4032
rect 16264 4020 16270 4072
rect 17880 4060 17908 4100
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 22557 4131 22615 4137
rect 22557 4097 22569 4131
rect 22603 4128 22615 4131
rect 23382 4128 23388 4140
rect 22603 4100 23388 4128
rect 22603 4097 22615 4100
rect 22557 4091 22615 4097
rect 23382 4088 23388 4100
rect 23440 4088 23446 4140
rect 24118 4088 24124 4140
rect 24176 4128 24182 4140
rect 24176 4100 25544 4128
rect 24176 4088 24182 4100
rect 20257 4063 20315 4069
rect 20257 4060 20269 4063
rect 17880 4032 20269 4060
rect 20257 4029 20269 4032
rect 20303 4060 20315 4063
rect 20809 4063 20867 4069
rect 20809 4060 20821 4063
rect 20303 4032 20821 4060
rect 20303 4029 20315 4032
rect 20257 4023 20315 4029
rect 20809 4029 20821 4032
rect 20855 4029 20867 4063
rect 20809 4023 20867 4029
rect 22186 4020 22192 4072
rect 22244 4060 22250 4072
rect 23937 4063 23995 4069
rect 23937 4060 23949 4063
rect 22244 4032 23949 4060
rect 22244 4020 22250 4032
rect 23937 4029 23949 4032
rect 23983 4029 23995 4063
rect 23937 4023 23995 4029
rect 24394 4020 24400 4072
rect 24452 4060 24458 4072
rect 24581 4063 24639 4069
rect 24581 4060 24593 4063
rect 24452 4032 24593 4060
rect 24452 4020 24458 4032
rect 24581 4029 24593 4032
rect 24627 4060 24639 4063
rect 25038 4060 25044 4072
rect 24627 4032 25044 4060
rect 24627 4029 24639 4032
rect 24581 4023 24639 4029
rect 25038 4020 25044 4032
rect 25096 4020 25102 4072
rect 25516 4069 25544 4100
rect 25501 4063 25559 4069
rect 25501 4029 25513 4063
rect 25547 4060 25559 4063
rect 26053 4063 26111 4069
rect 26053 4060 26065 4063
rect 25547 4032 26065 4060
rect 25547 4029 25559 4032
rect 25501 4023 25559 4029
rect 26053 4029 26065 4032
rect 26099 4029 26111 4063
rect 26053 4023 26111 4029
rect 15381 3995 15439 4001
rect 15381 3961 15393 3995
rect 15427 3992 15439 3995
rect 16114 3992 16120 4004
rect 15427 3964 16120 3992
rect 15427 3961 15439 3964
rect 15381 3955 15439 3961
rect 16114 3952 16120 3964
rect 16172 3952 16178 4004
rect 17770 3952 17776 4004
rect 17828 3992 17834 4004
rect 18370 3995 18428 4001
rect 18370 3992 18382 3995
rect 17828 3964 18382 3992
rect 17828 3952 17834 3964
rect 18370 3961 18382 3964
rect 18416 3992 18428 3995
rect 21130 3995 21188 4001
rect 21130 3992 21142 3995
rect 18416 3964 21142 3992
rect 18416 3961 18428 3964
rect 18370 3955 18428 3961
rect 20732 3936 20760 3964
rect 21130 3961 21142 3964
rect 21176 3992 21188 3995
rect 21450 3992 21456 4004
rect 21176 3964 21456 3992
rect 21176 3961 21188 3964
rect 21130 3955 21188 3961
rect 21450 3952 21456 3964
rect 21508 3992 21514 4004
rect 22005 3995 22063 4001
rect 22005 3992 22017 3995
rect 21508 3964 22017 3992
rect 21508 3952 21514 3964
rect 22005 3961 22017 3964
rect 22051 3961 22063 3995
rect 22005 3955 22063 3961
rect 15838 3924 15844 3936
rect 14700 3896 15332 3924
rect 15799 3896 15844 3924
rect 14700 3884 14706 3896
rect 15838 3884 15844 3896
rect 15896 3884 15902 3936
rect 16022 3884 16028 3936
rect 16080 3924 16086 3936
rect 16298 3924 16304 3936
rect 16080 3896 16304 3924
rect 16080 3884 16086 3896
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 19150 3884 19156 3936
rect 19208 3924 19214 3936
rect 19518 3924 19524 3936
rect 19208 3896 19524 3924
rect 19208 3884 19214 3896
rect 19518 3884 19524 3896
rect 19576 3924 19582 3936
rect 19613 3927 19671 3933
rect 19613 3924 19625 3927
rect 19576 3896 19625 3924
rect 19576 3884 19582 3896
rect 19613 3893 19625 3896
rect 19659 3893 19671 3927
rect 19613 3887 19671 3893
rect 19797 3927 19855 3933
rect 19797 3893 19809 3927
rect 19843 3924 19855 3927
rect 20162 3924 20168 3936
rect 19843 3896 20168 3924
rect 19843 3893 19855 3896
rect 19797 3887 19855 3893
rect 20162 3884 20168 3896
rect 20220 3884 20226 3936
rect 20714 3924 20720 3936
rect 20675 3896 20720 3924
rect 20714 3884 20720 3896
rect 20772 3884 20778 3936
rect 21726 3924 21732 3936
rect 21687 3896 21732 3924
rect 21726 3884 21732 3896
rect 21784 3884 21790 3936
rect 25406 3884 25412 3936
rect 25464 3924 25470 3936
rect 25685 3927 25743 3933
rect 25685 3924 25697 3927
rect 25464 3896 25697 3924
rect 25464 3884 25470 3896
rect 25685 3893 25697 3896
rect 25731 3893 25743 3927
rect 25685 3887 25743 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 6730 3720 6736 3732
rect 6691 3692 6736 3720
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 9815 3723 9873 3729
rect 9815 3720 9827 3723
rect 9732 3692 9827 3720
rect 9732 3680 9738 3692
rect 9815 3689 9827 3692
rect 9861 3689 9873 3723
rect 9815 3683 9873 3689
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 11333 3723 11391 3729
rect 11333 3720 11345 3723
rect 10928 3692 11345 3720
rect 10928 3680 10934 3692
rect 11333 3689 11345 3692
rect 11379 3689 11391 3723
rect 11333 3683 11391 3689
rect 5258 3652 5264 3664
rect 5219 3624 5264 3652
rect 5258 3612 5264 3624
rect 5316 3612 5322 3664
rect 8018 3612 8024 3664
rect 8076 3652 8082 3664
rect 8076 3624 11284 3652
rect 8076 3612 8082 3624
rect 2869 3587 2927 3593
rect 2869 3553 2881 3587
rect 2915 3584 2927 3587
rect 3050 3584 3056 3596
rect 2915 3556 3056 3584
rect 2915 3553 2927 3556
rect 2869 3547 2927 3553
rect 3050 3544 3056 3556
rect 3108 3544 3114 3596
rect 4500 3587 4558 3593
rect 4500 3553 4512 3587
rect 4546 3584 4558 3587
rect 5074 3584 5080 3596
rect 4546 3556 5080 3584
rect 4546 3553 4558 3556
rect 4500 3547 4558 3553
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 6638 3584 6644 3596
rect 6599 3556 6644 3584
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 8662 3584 8668 3596
rect 8623 3556 8668 3584
rect 8662 3544 8668 3556
rect 8720 3544 8726 3596
rect 9744 3587 9802 3593
rect 9744 3553 9756 3587
rect 9790 3584 9802 3587
rect 10134 3584 10140 3596
rect 9790 3556 10140 3584
rect 9790 3553 9802 3556
rect 9744 3547 9802 3553
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 5442 3516 5448 3528
rect 5403 3488 5448 3516
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3516 8815 3519
rect 10686 3516 10692 3528
rect 8803 3488 10692 3516
rect 8803 3485 8815 3488
rect 8757 3479 8815 3485
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 10962 3516 10968 3528
rect 10875 3488 10968 3516
rect 10962 3476 10968 3488
rect 11020 3516 11026 3528
rect 11146 3516 11152 3528
rect 11020 3488 11152 3516
rect 11020 3476 11026 3488
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 11256 3516 11284 3624
rect 11348 3584 11376 3683
rect 11606 3680 11612 3732
rect 11664 3720 11670 3732
rect 12161 3723 12219 3729
rect 12161 3720 12173 3723
rect 11664 3692 12173 3720
rect 11664 3680 11670 3692
rect 12161 3689 12173 3692
rect 12207 3689 12219 3723
rect 13998 3720 14004 3732
rect 13959 3692 14004 3720
rect 12161 3683 12219 3689
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 14182 3680 14188 3732
rect 14240 3720 14246 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 14240 3692 15025 3720
rect 14240 3680 14246 3692
rect 15013 3689 15025 3692
rect 15059 3689 15071 3723
rect 15013 3683 15071 3689
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 15473 3723 15531 3729
rect 15473 3720 15485 3723
rect 15344 3692 15485 3720
rect 15344 3680 15350 3692
rect 15473 3689 15485 3692
rect 15519 3689 15531 3723
rect 17126 3720 17132 3732
rect 17087 3692 17132 3720
rect 15473 3683 15531 3689
rect 17126 3680 17132 3692
rect 17184 3680 17190 3732
rect 17770 3680 17776 3732
rect 17828 3720 17834 3732
rect 17865 3723 17923 3729
rect 17865 3720 17877 3723
rect 17828 3692 17877 3720
rect 17828 3680 17834 3692
rect 17865 3689 17877 3692
rect 17911 3689 17923 3723
rect 17865 3683 17923 3689
rect 20162 3680 20168 3732
rect 20220 3720 20226 3732
rect 23566 3720 23572 3732
rect 20220 3692 23474 3720
rect 23527 3692 23572 3720
rect 20220 3680 20226 3692
rect 12529 3655 12587 3661
rect 12529 3621 12541 3655
rect 12575 3652 12587 3655
rect 12618 3652 12624 3664
rect 12575 3624 12624 3652
rect 12575 3621 12587 3624
rect 12529 3615 12587 3621
rect 12618 3612 12624 3624
rect 12676 3612 12682 3664
rect 13075 3655 13133 3661
rect 13075 3621 13087 3655
rect 13121 3621 13133 3655
rect 13075 3615 13133 3621
rect 11882 3584 11888 3596
rect 11348 3556 11888 3584
rect 11882 3544 11888 3556
rect 11940 3584 11946 3596
rect 13090 3584 13118 3615
rect 14918 3612 14924 3664
rect 14976 3652 14982 3664
rect 15749 3655 15807 3661
rect 15749 3652 15761 3655
rect 14976 3624 15761 3652
rect 14976 3612 14982 3624
rect 15749 3621 15761 3624
rect 15795 3652 15807 3655
rect 15933 3655 15991 3661
rect 15933 3652 15945 3655
rect 15795 3624 15945 3652
rect 15795 3621 15807 3624
rect 15749 3615 15807 3621
rect 15933 3621 15945 3624
rect 15979 3621 15991 3655
rect 15933 3615 15991 3621
rect 16022 3612 16028 3664
rect 16080 3652 16086 3664
rect 16080 3624 16125 3652
rect 16080 3612 16086 3624
rect 18782 3612 18788 3664
rect 18840 3652 18846 3664
rect 19334 3652 19340 3664
rect 18840 3624 19340 3652
rect 18840 3612 18846 3624
rect 19334 3612 19340 3624
rect 19392 3652 19398 3664
rect 19429 3655 19487 3661
rect 19429 3652 19441 3655
rect 19392 3624 19441 3652
rect 19392 3612 19398 3624
rect 19429 3621 19441 3624
rect 19475 3621 19487 3655
rect 19429 3615 19487 3621
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 21222 3655 21280 3661
rect 21222 3652 21234 3655
rect 20772 3624 21234 3652
rect 20772 3612 20778 3624
rect 21222 3621 21234 3624
rect 21268 3621 21280 3655
rect 23446 3652 23474 3692
rect 23566 3680 23572 3692
rect 23624 3680 23630 3732
rect 24394 3720 24400 3732
rect 24355 3692 24400 3720
rect 24394 3680 24400 3692
rect 24452 3680 24458 3732
rect 24854 3680 24860 3732
rect 24912 3720 24918 3732
rect 24912 3692 25084 3720
rect 24912 3680 24918 3692
rect 24946 3652 24952 3664
rect 23446 3624 24952 3652
rect 21222 3615 21280 3621
rect 24946 3612 24952 3624
rect 25004 3612 25010 3664
rect 25056 3661 25084 3692
rect 25041 3655 25099 3661
rect 25041 3621 25053 3655
rect 25087 3621 25099 3655
rect 25041 3615 25099 3621
rect 11940 3556 13118 3584
rect 11940 3544 11946 3556
rect 16758 3544 16764 3596
rect 16816 3584 16822 3596
rect 19061 3587 19119 3593
rect 19061 3584 19073 3587
rect 16816 3556 19073 3584
rect 16816 3544 16822 3556
rect 19061 3553 19073 3556
rect 19107 3553 19119 3587
rect 19061 3547 19119 3553
rect 11256 3488 15884 3516
rect 4571 3451 4629 3457
rect 4571 3417 4583 3451
rect 4617 3448 4629 3451
rect 10781 3451 10839 3457
rect 10781 3448 10793 3451
rect 4617 3420 10793 3448
rect 4617 3417 4629 3420
rect 4571 3411 4629 3417
rect 10781 3417 10793 3420
rect 10827 3448 10839 3451
rect 10870 3448 10876 3460
rect 10827 3420 10876 3448
rect 10827 3417 10839 3420
rect 10781 3411 10839 3417
rect 10870 3408 10876 3420
rect 10928 3408 10934 3460
rect 12526 3408 12532 3460
rect 12584 3448 12590 3460
rect 14277 3451 14335 3457
rect 14277 3448 14289 3451
rect 12584 3420 14289 3448
rect 12584 3408 12590 3420
rect 14277 3417 14289 3420
rect 14323 3417 14335 3451
rect 15856 3448 15884 3488
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 16942 3516 16948 3528
rect 16080 3488 16948 3516
rect 16080 3476 16086 3488
rect 16942 3476 16948 3488
rect 17000 3516 17006 3528
rect 17497 3519 17555 3525
rect 17497 3516 17509 3519
rect 17000 3488 17509 3516
rect 17000 3476 17006 3488
rect 17497 3485 17509 3488
rect 17543 3485 17555 3519
rect 17497 3479 17555 3485
rect 17586 3476 17592 3528
rect 17644 3516 17650 3528
rect 18693 3519 18751 3525
rect 18693 3516 18705 3519
rect 17644 3488 18705 3516
rect 17644 3476 17650 3488
rect 18693 3485 18705 3488
rect 18739 3485 18751 3519
rect 19076 3516 19104 3547
rect 23474 3544 23480 3596
rect 23532 3584 23538 3596
rect 23532 3556 23577 3584
rect 23532 3544 23538 3556
rect 19337 3519 19395 3525
rect 19337 3516 19349 3519
rect 19076 3488 19349 3516
rect 18693 3479 18751 3485
rect 19337 3485 19349 3488
rect 19383 3485 19395 3519
rect 19337 3479 19395 3485
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 19613 3519 19671 3525
rect 19613 3516 19625 3519
rect 19576 3488 19625 3516
rect 19576 3476 19582 3488
rect 19613 3485 19625 3488
rect 19659 3485 19671 3519
rect 20898 3516 20904 3528
rect 20859 3488 20904 3516
rect 19613 3479 19671 3485
rect 20898 3476 20904 3488
rect 20956 3476 20962 3528
rect 25222 3516 25228 3528
rect 25183 3488 25228 3516
rect 25222 3476 25228 3488
rect 25280 3476 25286 3528
rect 16485 3451 16543 3457
rect 16485 3448 16497 3451
rect 15856 3420 16497 3448
rect 14277 3411 14335 3417
rect 16485 3417 16497 3420
rect 16531 3448 16543 3451
rect 18322 3448 18328 3460
rect 16531 3420 18328 3448
rect 16531 3417 16543 3420
rect 16485 3411 16543 3417
rect 18322 3408 18328 3420
rect 18380 3408 18386 3460
rect 20070 3408 20076 3460
rect 20128 3448 20134 3460
rect 23750 3448 23756 3460
rect 20128 3420 23756 3448
rect 20128 3408 20134 3420
rect 23750 3408 23756 3420
rect 23808 3408 23814 3460
rect 3099 3383 3157 3389
rect 3099 3349 3111 3383
rect 3145 3380 3157 3383
rect 7466 3380 7472 3392
rect 3145 3352 7472 3380
rect 3145 3349 3157 3352
rect 3099 3343 3157 3349
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 7745 3383 7803 3389
rect 7745 3349 7757 3383
rect 7791 3380 7803 3383
rect 8018 3380 8024 3392
rect 7791 3352 8024 3380
rect 7791 3349 7803 3352
rect 7745 3343 7803 3349
rect 8018 3340 8024 3352
rect 8076 3340 8082 3392
rect 10962 3340 10968 3392
rect 11020 3380 11026 3392
rect 11885 3383 11943 3389
rect 11885 3380 11897 3383
rect 11020 3352 11897 3380
rect 11020 3340 11026 3352
rect 11885 3349 11897 3352
rect 11931 3349 11943 3383
rect 11885 3343 11943 3349
rect 12618 3340 12624 3392
rect 12676 3380 12682 3392
rect 13633 3383 13691 3389
rect 13633 3380 13645 3383
rect 12676 3352 13645 3380
rect 12676 3340 12682 3352
rect 13633 3349 13645 3352
rect 13679 3349 13691 3383
rect 14642 3380 14648 3392
rect 14603 3352 14648 3380
rect 13633 3343 13691 3349
rect 14642 3340 14648 3352
rect 14700 3380 14706 3392
rect 15562 3380 15568 3392
rect 14700 3352 15568 3380
rect 14700 3340 14706 3352
rect 15562 3340 15568 3352
rect 15620 3340 15626 3392
rect 15749 3383 15807 3389
rect 15749 3349 15761 3383
rect 15795 3380 15807 3383
rect 16206 3380 16212 3392
rect 15795 3352 16212 3380
rect 15795 3349 15807 3352
rect 15749 3343 15807 3349
rect 16206 3340 16212 3352
rect 16264 3380 16270 3392
rect 17586 3380 17592 3392
rect 16264 3352 17592 3380
rect 16264 3340 16270 3352
rect 17586 3340 17592 3352
rect 17644 3340 17650 3392
rect 18414 3380 18420 3392
rect 18375 3352 18420 3380
rect 18414 3340 18420 3352
rect 18472 3340 18478 3392
rect 20254 3380 20260 3392
rect 20215 3352 20260 3380
rect 20254 3340 20260 3352
rect 20312 3340 20318 3392
rect 20622 3380 20628 3392
rect 20583 3352 20628 3380
rect 20622 3340 20628 3352
rect 20680 3340 20686 3392
rect 21358 3340 21364 3392
rect 21416 3380 21422 3392
rect 21821 3383 21879 3389
rect 21821 3380 21833 3383
rect 21416 3352 21833 3380
rect 21416 3340 21422 3352
rect 21821 3349 21833 3352
rect 21867 3349 21879 3383
rect 21821 3343 21879 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 2409 3179 2467 3185
rect 2409 3145 2421 3179
rect 2455 3176 2467 3179
rect 2498 3176 2504 3188
rect 2455 3148 2504 3176
rect 2455 3145 2467 3148
rect 2409 3139 2467 3145
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 3050 3176 3056 3188
rect 3011 3148 3056 3176
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 3283 3179 3341 3185
rect 3283 3145 3295 3179
rect 3329 3176 3341 3179
rect 8938 3176 8944 3188
rect 3329 3148 8944 3176
rect 3329 3145 3341 3148
rect 3283 3139 3341 3145
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9306 3176 9312 3188
rect 9267 3148 9312 3176
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 11422 3176 11428 3188
rect 9548 3148 11428 3176
rect 9548 3136 9554 3148
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 11514 3136 11520 3188
rect 11572 3176 11578 3188
rect 19334 3176 19340 3188
rect 11572 3148 19012 3176
rect 19295 3148 19340 3176
rect 11572 3136 11578 3148
rect 3694 3108 3700 3120
rect 3655 3080 3700 3108
rect 3694 3068 3700 3080
rect 3752 3068 3758 3120
rect 5258 3108 5264 3120
rect 3804 3080 5264 3108
rect 2200 2975 2258 2981
rect 2200 2941 2212 2975
rect 2246 2941 2258 2975
rect 2200 2935 2258 2941
rect 3212 2975 3270 2981
rect 3212 2941 3224 2975
rect 3258 2972 3270 2975
rect 3712 2972 3740 3068
rect 3258 2944 3740 2972
rect 3258 2941 3270 2944
rect 3212 2935 3270 2941
rect 2215 2904 2243 2935
rect 2685 2907 2743 2913
rect 2685 2904 2697 2907
rect 2215 2876 2697 2904
rect 2685 2873 2697 2876
rect 2731 2904 2743 2907
rect 3804 2904 3832 3080
rect 5258 3068 5264 3080
rect 5316 3068 5322 3120
rect 8662 3108 8668 3120
rect 8623 3080 8668 3108
rect 8662 3068 8668 3080
rect 8720 3068 8726 3120
rect 9122 3068 9128 3120
rect 9180 3108 9186 3120
rect 10597 3111 10655 3117
rect 10597 3108 10609 3111
rect 9180 3080 10609 3108
rect 9180 3068 9186 3080
rect 10597 3077 10609 3080
rect 10643 3077 10655 3111
rect 11882 3108 11888 3120
rect 11843 3080 11888 3108
rect 10597 3071 10655 3077
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9079 3012 9812 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 9784 2984 9812 3012
rect 4192 2975 4250 2981
rect 4192 2941 4204 2975
rect 4238 2941 4250 2975
rect 5350 2972 5356 2984
rect 5311 2944 5356 2972
rect 4192 2935 4250 2941
rect 4207 2904 4235 2935
rect 5350 2932 5356 2944
rect 5408 2932 5414 2984
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2972 7619 2975
rect 8294 2972 8300 2984
rect 7607 2944 8300 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 8294 2932 8300 2944
rect 8352 2932 8358 2984
rect 9490 2972 9496 2984
rect 9451 2944 9496 2972
rect 9490 2932 9496 2944
rect 9548 2932 9554 2984
rect 9766 2972 9772 2984
rect 9727 2944 9772 2972
rect 9766 2932 9772 2944
rect 9824 2932 9830 2984
rect 4617 2907 4675 2913
rect 4617 2904 4629 2907
rect 2731 2876 3832 2904
rect 4126 2876 4629 2904
rect 2731 2873 2743 2876
rect 2685 2867 2743 2873
rect 1854 2796 1860 2848
rect 1912 2836 1918 2848
rect 4126 2836 4154 2876
rect 4617 2873 4629 2876
rect 4663 2873 4675 2907
rect 4617 2867 4675 2873
rect 5905 2907 5963 2913
rect 5905 2873 5917 2907
rect 5951 2904 5963 2907
rect 8202 2904 8208 2916
rect 5951 2876 8208 2904
rect 5951 2873 5963 2876
rect 5905 2867 5963 2873
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 8386 2904 8392 2916
rect 8347 2876 8392 2904
rect 8386 2864 8392 2876
rect 8444 2864 8450 2916
rect 8662 2864 8668 2916
rect 8720 2904 8726 2916
rect 10612 2904 10640 3071
rect 11882 3068 11888 3080
rect 11940 3108 11946 3120
rect 13449 3111 13507 3117
rect 13449 3108 13461 3111
rect 11940 3080 13461 3108
rect 11940 3068 11946 3080
rect 13449 3077 13461 3080
rect 13495 3108 13507 3111
rect 13909 3111 13967 3117
rect 13909 3108 13921 3111
rect 13495 3080 13921 3108
rect 13495 3077 13507 3080
rect 13449 3071 13507 3077
rect 13909 3077 13921 3080
rect 13955 3077 13967 3111
rect 13909 3071 13967 3077
rect 10870 3040 10876 3052
rect 10831 3012 10876 3040
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11112 3012 11529 3040
rect 11112 3000 11118 3012
rect 11517 3009 11529 3012
rect 11563 3040 11575 3043
rect 12526 3040 12532 3052
rect 11563 3012 12532 3040
rect 11563 3009 11575 3012
rect 11517 3003 11575 3009
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 12802 3040 12808 3052
rect 12763 3012 12808 3040
rect 12802 3000 12808 3012
rect 12860 3000 12866 3052
rect 13354 3000 13360 3052
rect 13412 3040 13418 3052
rect 13924 3040 13952 3071
rect 15565 3043 15623 3049
rect 15565 3040 15577 3043
rect 13412 3012 13814 3040
rect 13924 3012 15577 3040
rect 13412 3000 13418 3012
rect 13786 2972 13814 3012
rect 14090 2972 14096 2984
rect 13786 2944 14096 2972
rect 14090 2932 14096 2944
rect 14148 2932 14154 2984
rect 10962 2904 10968 2916
rect 8720 2876 10364 2904
rect 10612 2876 10968 2904
rect 8720 2864 8726 2876
rect 1912 2808 4154 2836
rect 4295 2839 4353 2845
rect 1912 2796 1918 2808
rect 4295 2805 4307 2839
rect 4341 2836 4353 2839
rect 4890 2836 4896 2848
rect 4341 2808 4896 2836
rect 4341 2805 4353 2808
rect 4295 2799 4353 2805
rect 4890 2796 4896 2808
rect 4948 2796 4954 2848
rect 5074 2836 5080 2848
rect 5035 2808 5080 2836
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 6546 2836 6552 2848
rect 6507 2808 6552 2836
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 10229 2839 10287 2845
rect 10229 2836 10241 2839
rect 10192 2808 10241 2836
rect 10192 2796 10198 2808
rect 10229 2805 10241 2808
rect 10275 2805 10287 2839
rect 10336 2836 10364 2876
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 12161 2907 12219 2913
rect 12161 2904 12173 2907
rect 11624 2876 12173 2904
rect 11624 2836 11652 2876
rect 12161 2873 12173 2876
rect 12207 2873 12219 2907
rect 12161 2867 12219 2873
rect 10336 2808 11652 2836
rect 12176 2836 12204 2867
rect 12618 2864 12624 2916
rect 12676 2904 12682 2916
rect 14470 2913 14498 3012
rect 15565 3009 15577 3012
rect 15611 3040 15623 3043
rect 15657 3043 15715 3049
rect 15657 3040 15669 3043
rect 15611 3012 15669 3040
rect 15611 3009 15623 3012
rect 15565 3003 15623 3009
rect 15657 3009 15669 3012
rect 15703 3009 15715 3043
rect 15838 3040 15844 3052
rect 15799 3012 15844 3040
rect 15657 3003 15715 3009
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 17221 3043 17279 3049
rect 17221 3009 17233 3043
rect 17267 3040 17279 3043
rect 18138 3040 18144 3052
rect 17267 3012 18144 3040
rect 17267 3009 17279 3012
rect 17221 3003 17279 3009
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 18322 3000 18328 3052
rect 18380 3040 18386 3052
rect 18417 3043 18475 3049
rect 18417 3040 18429 3043
rect 18380 3012 18429 3040
rect 18380 3000 18386 3012
rect 18417 3009 18429 3012
rect 18463 3009 18475 3043
rect 18417 3003 18475 3009
rect 16298 2972 16304 2984
rect 15304 2944 16304 2972
rect 14455 2907 14513 2913
rect 12676 2876 12769 2904
rect 12676 2864 12682 2876
rect 14455 2873 14467 2907
rect 14501 2873 14513 2907
rect 14455 2867 14513 2873
rect 12636 2836 12664 2864
rect 15304 2848 15332 2944
rect 16298 2932 16304 2944
rect 16356 2972 16362 2984
rect 16761 2975 16819 2981
rect 16761 2972 16773 2975
rect 16356 2944 16773 2972
rect 16356 2932 16362 2944
rect 16761 2941 16773 2944
rect 16807 2941 16819 2975
rect 18984 2972 19012 3148
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 19889 3179 19947 3185
rect 19889 3176 19901 3179
rect 19628 3148 19901 3176
rect 19058 3068 19064 3120
rect 19116 3108 19122 3120
rect 19628 3108 19656 3148
rect 19889 3145 19901 3148
rect 19935 3145 19947 3179
rect 19889 3139 19947 3145
rect 20898 3136 20904 3188
rect 20956 3176 20962 3188
rect 22465 3179 22523 3185
rect 22465 3176 22477 3179
rect 20956 3148 22477 3176
rect 20956 3136 20962 3148
rect 22465 3145 22477 3148
rect 22511 3145 22523 3179
rect 22465 3139 22523 3145
rect 23109 3179 23167 3185
rect 23109 3145 23121 3179
rect 23155 3176 23167 3179
rect 23474 3176 23480 3188
rect 23155 3148 23480 3176
rect 23155 3145 23167 3148
rect 23109 3139 23167 3145
rect 23474 3136 23480 3148
rect 23532 3136 23538 3188
rect 19116 3080 19656 3108
rect 19116 3068 19122 3080
rect 23382 3068 23388 3120
rect 23440 3108 23446 3120
rect 25409 3111 25467 3117
rect 25409 3108 25421 3111
rect 23440 3080 25421 3108
rect 23440 3068 23446 3080
rect 25409 3077 25421 3080
rect 25455 3077 25467 3111
rect 25409 3071 25467 3077
rect 20254 3000 20260 3052
rect 20312 3040 20318 3052
rect 21177 3043 21235 3049
rect 21177 3040 21189 3043
rect 20312 3012 21189 3040
rect 20312 3000 20318 3012
rect 21177 3009 21189 3012
rect 21223 3009 21235 3043
rect 23750 3040 23756 3052
rect 23711 3012 23756 3040
rect 21177 3003 21235 3009
rect 23750 3000 23756 3012
rect 23808 3000 23814 3052
rect 23934 3000 23940 3052
rect 23992 3040 23998 3052
rect 24029 3043 24087 3049
rect 24029 3040 24041 3043
rect 23992 3012 24041 3040
rect 23992 3000 23998 3012
rect 24029 3009 24041 3012
rect 24075 3009 24087 3043
rect 24029 3003 24087 3009
rect 19426 2972 19432 2984
rect 18984 2944 19432 2972
rect 16761 2935 16819 2941
rect 19426 2932 19432 2944
rect 19484 2972 19490 2984
rect 19613 2975 19671 2981
rect 19613 2972 19625 2975
rect 19484 2944 19625 2972
rect 19484 2932 19490 2944
rect 19613 2941 19625 2944
rect 19659 2941 19671 2975
rect 19613 2935 19671 2941
rect 19797 2975 19855 2981
rect 19797 2941 19809 2975
rect 19843 2941 19855 2975
rect 19797 2935 19855 2941
rect 21821 2975 21879 2981
rect 21821 2941 21833 2975
rect 21867 2972 21879 2975
rect 23290 2972 23296 2984
rect 21867 2944 23296 2972
rect 21867 2941 21879 2944
rect 21821 2935 21879 2941
rect 15565 2907 15623 2913
rect 15565 2873 15577 2907
rect 15611 2904 15623 2907
rect 16162 2907 16220 2913
rect 16162 2904 16174 2907
rect 15611 2876 16174 2904
rect 15611 2873 15623 2876
rect 15565 2867 15623 2873
rect 16162 2873 16174 2876
rect 16208 2904 16220 2907
rect 17497 2907 17555 2913
rect 17497 2904 17509 2907
rect 16208 2876 17509 2904
rect 16208 2873 16220 2876
rect 16162 2867 16220 2873
rect 17497 2873 17509 2876
rect 17543 2904 17555 2907
rect 17770 2904 17776 2916
rect 17543 2876 17776 2904
rect 17543 2873 17555 2876
rect 17497 2867 17555 2873
rect 17770 2864 17776 2876
rect 17828 2864 17834 2916
rect 18233 2907 18291 2913
rect 18233 2873 18245 2907
rect 18279 2873 18291 2907
rect 18233 2867 18291 2873
rect 12176 2808 12664 2836
rect 10229 2799 10287 2805
rect 14734 2796 14740 2848
rect 14792 2836 14798 2848
rect 15013 2839 15071 2845
rect 15013 2836 15025 2839
rect 14792 2808 15025 2836
rect 14792 2796 14798 2808
rect 15013 2805 15025 2808
rect 15059 2805 15071 2839
rect 15286 2836 15292 2848
rect 15247 2808 15292 2836
rect 15013 2799 15071 2805
rect 15286 2796 15292 2808
rect 15344 2796 15350 2848
rect 18046 2796 18052 2848
rect 18104 2836 18110 2848
rect 18248 2836 18276 2867
rect 19334 2864 19340 2916
rect 19392 2904 19398 2916
rect 19812 2904 19840 2935
rect 23290 2932 23296 2944
rect 23348 2932 23354 2984
rect 25130 2932 25136 2984
rect 25188 2972 25194 2984
rect 25225 2975 25283 2981
rect 25225 2972 25237 2975
rect 25188 2944 25237 2972
rect 25188 2932 25194 2944
rect 25225 2941 25237 2944
rect 25271 2972 25283 2975
rect 25777 2975 25835 2981
rect 25777 2972 25789 2975
rect 25271 2944 25789 2972
rect 25271 2941 25283 2944
rect 25225 2935 25283 2941
rect 25777 2941 25789 2944
rect 25823 2941 25835 2975
rect 25777 2935 25835 2941
rect 20441 2907 20499 2913
rect 20441 2904 20453 2907
rect 19392 2876 20453 2904
rect 19392 2864 19398 2876
rect 20441 2873 20453 2876
rect 20487 2873 20499 2907
rect 20441 2867 20499 2873
rect 21269 2907 21327 2913
rect 21269 2873 21281 2907
rect 21315 2904 21327 2907
rect 22097 2907 22155 2913
rect 22097 2904 22109 2907
rect 21315 2876 22109 2904
rect 21315 2873 21327 2876
rect 21269 2867 21327 2873
rect 22097 2873 22109 2876
rect 22143 2873 22155 2907
rect 22097 2867 22155 2873
rect 18104 2808 18276 2836
rect 18104 2796 18110 2808
rect 19978 2796 19984 2848
rect 20036 2836 20042 2848
rect 20714 2836 20720 2848
rect 20036 2808 20720 2836
rect 20036 2796 20042 2808
rect 20714 2796 20720 2808
rect 20772 2836 20778 2848
rect 20901 2839 20959 2845
rect 20901 2836 20913 2839
rect 20772 2808 20913 2836
rect 20772 2796 20778 2808
rect 20901 2805 20913 2808
rect 20947 2805 20959 2839
rect 20901 2799 20959 2805
rect 20990 2796 20996 2848
rect 21048 2836 21054 2848
rect 21284 2836 21312 2867
rect 23842 2864 23848 2916
rect 23900 2904 23906 2916
rect 23900 2876 23945 2904
rect 23900 2864 23906 2876
rect 21048 2808 21312 2836
rect 21048 2796 21054 2808
rect 21358 2796 21364 2848
rect 21416 2836 21422 2848
rect 23385 2839 23443 2845
rect 23385 2836 23397 2839
rect 21416 2808 23397 2836
rect 21416 2796 21422 2808
rect 23385 2805 23397 2808
rect 23431 2836 23443 2839
rect 23658 2836 23664 2848
rect 23431 2808 23664 2836
rect 23431 2805 23443 2808
rect 23385 2799 23443 2805
rect 23658 2796 23664 2808
rect 23716 2796 23722 2848
rect 24854 2836 24860 2848
rect 24815 2808 24860 2836
rect 24854 2796 24860 2808
rect 24912 2796 24918 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1535 2635 1593 2641
rect 1535 2601 1547 2635
rect 1581 2632 1593 2635
rect 1670 2632 1676 2644
rect 1581 2604 1676 2632
rect 1581 2601 1593 2604
rect 1535 2595 1593 2601
rect 1670 2592 1676 2604
rect 1728 2592 1734 2644
rect 2547 2635 2605 2641
rect 2547 2601 2559 2635
rect 2593 2632 2605 2635
rect 4246 2632 4252 2644
rect 2593 2604 4252 2632
rect 2593 2601 2605 2604
rect 2547 2595 2605 2601
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 4387 2635 4445 2641
rect 4387 2601 4399 2635
rect 4433 2632 4445 2635
rect 4522 2632 4528 2644
rect 4433 2604 4528 2632
rect 4433 2601 4445 2604
rect 4387 2595 4445 2601
rect 4522 2592 4528 2604
rect 4580 2592 4586 2644
rect 7239 2635 7297 2641
rect 7239 2601 7251 2635
rect 7285 2632 7297 2635
rect 7926 2632 7932 2644
rect 7285 2604 7932 2632
rect 7285 2601 7297 2604
rect 7239 2595 7297 2601
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 9309 2635 9367 2641
rect 9309 2601 9321 2635
rect 9355 2632 9367 2635
rect 9490 2632 9496 2644
rect 9355 2604 9496 2632
rect 9355 2601 9367 2604
rect 9309 2595 9367 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 9858 2592 9864 2644
rect 9916 2632 9922 2644
rect 9953 2635 10011 2641
rect 9953 2632 9965 2635
rect 9916 2604 9965 2632
rect 9916 2592 9922 2604
rect 9953 2601 9965 2604
rect 9999 2632 10011 2635
rect 11146 2632 11152 2644
rect 9999 2604 10364 2632
rect 11107 2604 11152 2632
rect 9999 2601 10011 2604
rect 9953 2595 10011 2601
rect 4890 2524 4896 2576
rect 4948 2564 4954 2576
rect 10226 2564 10232 2576
rect 4948 2536 10232 2564
rect 4948 2524 4954 2536
rect 10226 2524 10232 2536
rect 10284 2524 10290 2576
rect 10336 2573 10364 2604
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11974 2632 11980 2644
rect 11935 2604 11980 2632
rect 11974 2592 11980 2604
rect 12032 2632 12038 2644
rect 12710 2632 12716 2644
rect 12032 2604 12716 2632
rect 12032 2592 12038 2604
rect 12710 2592 12716 2604
rect 12768 2592 12774 2644
rect 14090 2632 14096 2644
rect 14051 2604 14096 2632
rect 14090 2592 14096 2604
rect 14148 2592 14154 2644
rect 15838 2592 15844 2644
rect 15896 2632 15902 2644
rect 16485 2635 16543 2641
rect 16485 2632 16497 2635
rect 15896 2604 16497 2632
rect 15896 2592 15902 2604
rect 16485 2601 16497 2604
rect 16531 2601 16543 2635
rect 16942 2632 16948 2644
rect 16903 2604 16948 2632
rect 16485 2595 16543 2601
rect 16942 2592 16948 2604
rect 17000 2592 17006 2644
rect 17313 2635 17371 2641
rect 17313 2601 17325 2635
rect 17359 2632 17371 2635
rect 20070 2632 20076 2644
rect 17359 2604 20076 2632
rect 17359 2601 17371 2604
rect 17313 2595 17371 2601
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 21726 2592 21732 2644
rect 21784 2632 21790 2644
rect 23753 2635 23811 2641
rect 23753 2632 23765 2635
rect 21784 2604 23765 2632
rect 21784 2592 21790 2604
rect 23753 2601 23765 2604
rect 23799 2632 23811 2635
rect 23799 2604 24256 2632
rect 23799 2601 23811 2604
rect 23753 2595 23811 2601
rect 10321 2567 10379 2573
rect 10321 2533 10333 2567
rect 10367 2533 10379 2567
rect 10321 2527 10379 2533
rect 10873 2567 10931 2573
rect 10873 2533 10885 2567
rect 10919 2564 10931 2567
rect 11054 2564 11060 2576
rect 10919 2536 11060 2564
rect 10919 2533 10931 2536
rect 10873 2527 10931 2533
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 12805 2567 12863 2573
rect 12805 2564 12817 2567
rect 12360 2536 12817 2564
rect 658 2456 664 2508
rect 716 2496 722 2508
rect 1432 2499 1490 2505
rect 1432 2496 1444 2499
rect 716 2468 1444 2496
rect 716 2456 722 2468
rect 1432 2465 1444 2468
rect 1478 2496 1490 2499
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 1478 2468 1869 2496
rect 1478 2465 1490 2468
rect 1432 2459 1490 2465
rect 1857 2465 1869 2468
rect 1903 2465 1915 2499
rect 1857 2459 1915 2465
rect 2476 2499 2534 2505
rect 2476 2465 2488 2499
rect 2522 2496 2534 2499
rect 2866 2496 2872 2508
rect 2522 2468 2872 2496
rect 2522 2465 2534 2468
rect 2476 2459 2534 2465
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 4316 2499 4374 2505
rect 4316 2465 4328 2499
rect 4362 2496 4374 2499
rect 5169 2499 5227 2505
rect 4362 2468 4844 2496
rect 4362 2465 4374 2468
rect 4316 2459 4374 2465
rect 2866 2292 2872 2304
rect 2827 2264 2872 2292
rect 2866 2252 2872 2264
rect 2924 2252 2930 2304
rect 4816 2301 4844 2468
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5905 2499 5963 2505
rect 5905 2496 5917 2499
rect 5215 2468 5917 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5905 2465 5917 2468
rect 5951 2496 5963 2499
rect 6086 2496 6092 2508
rect 5951 2468 6092 2496
rect 5951 2465 5963 2468
rect 5905 2459 5963 2465
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 7168 2499 7226 2505
rect 7168 2465 7180 2499
rect 7214 2496 7226 2499
rect 8021 2499 8079 2505
rect 7214 2468 7696 2496
rect 7214 2465 7226 2468
rect 7168 2459 7226 2465
rect 5994 2428 6000 2440
rect 5955 2400 6000 2428
rect 5994 2388 6000 2400
rect 6052 2388 6058 2440
rect 7668 2369 7696 2468
rect 8021 2465 8033 2499
rect 8067 2496 8079 2499
rect 8754 2496 8760 2508
rect 8067 2468 8760 2496
rect 8067 2465 8079 2468
rect 8021 2459 8079 2465
rect 8754 2456 8760 2468
rect 8812 2456 8818 2508
rect 8849 2499 8907 2505
rect 8849 2465 8861 2499
rect 8895 2496 8907 2499
rect 10042 2496 10048 2508
rect 8895 2468 10048 2496
rect 8895 2465 8907 2468
rect 8849 2459 8907 2465
rect 10042 2456 10048 2468
rect 10100 2456 10106 2508
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 10284 2400 11529 2428
rect 10284 2388 10290 2400
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 7653 2363 7711 2369
rect 7653 2329 7665 2363
rect 7699 2360 7711 2363
rect 8846 2360 8852 2372
rect 7699 2332 8852 2360
rect 7699 2329 7711 2332
rect 7653 2323 7711 2329
rect 8846 2320 8852 2332
rect 8904 2320 8910 2372
rect 8956 2332 10364 2360
rect 4801 2295 4859 2301
rect 4801 2261 4813 2295
rect 4847 2292 4859 2295
rect 8956 2292 8984 2332
rect 4847 2264 8984 2292
rect 10336 2292 10364 2332
rect 10686 2320 10692 2372
rect 10744 2360 10750 2372
rect 12360 2369 12388 2536
rect 12805 2533 12817 2536
rect 12851 2533 12863 2567
rect 15657 2567 15715 2573
rect 15657 2564 15669 2567
rect 12805 2527 12863 2533
rect 15212 2536 15669 2564
rect 13630 2456 13636 2508
rect 13688 2496 13694 2508
rect 13725 2499 13783 2505
rect 13725 2496 13737 2499
rect 13688 2468 13737 2496
rect 13688 2456 13694 2468
rect 13725 2465 13737 2468
rect 13771 2496 13783 2499
rect 14277 2499 14335 2505
rect 14277 2496 14289 2499
rect 13771 2468 14289 2496
rect 13771 2465 13783 2468
rect 13725 2459 13783 2465
rect 14277 2465 14289 2468
rect 14323 2465 14335 2499
rect 14277 2459 14335 2465
rect 12710 2428 12716 2440
rect 12671 2400 12716 2428
rect 12710 2388 12716 2400
rect 12768 2388 12774 2440
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 12989 2431 13047 2437
rect 12989 2428 13001 2431
rect 12860 2400 13001 2428
rect 12860 2388 12866 2400
rect 12989 2397 13001 2400
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 13596 2400 13814 2428
rect 13596 2388 13602 2400
rect 12345 2363 12403 2369
rect 12345 2360 12357 2363
rect 10744 2332 12357 2360
rect 10744 2320 10750 2332
rect 12345 2329 12357 2332
rect 12391 2329 12403 2363
rect 13786 2360 13814 2400
rect 14734 2388 14740 2440
rect 14792 2428 14798 2440
rect 15212 2437 15240 2536
rect 15657 2533 15669 2536
rect 15703 2533 15715 2567
rect 16206 2564 16212 2576
rect 16167 2536 16212 2564
rect 15657 2527 15715 2533
rect 16206 2524 16212 2536
rect 16264 2524 16270 2576
rect 17586 2524 17592 2576
rect 17644 2564 17650 2576
rect 18414 2564 18420 2576
rect 17644 2536 18420 2564
rect 17644 2524 17650 2536
rect 18414 2524 18420 2536
rect 18472 2564 18478 2576
rect 18785 2567 18843 2573
rect 18785 2564 18797 2567
rect 18472 2536 18797 2564
rect 18472 2524 18478 2536
rect 18785 2533 18797 2536
rect 18831 2533 18843 2567
rect 18785 2527 18843 2533
rect 19337 2567 19395 2573
rect 19337 2533 19349 2567
rect 19383 2564 19395 2567
rect 19518 2564 19524 2576
rect 19383 2536 19524 2564
rect 19383 2533 19395 2536
rect 19337 2527 19395 2533
rect 19518 2524 19524 2536
rect 19576 2524 19582 2576
rect 20898 2524 20904 2576
rect 20956 2564 20962 2576
rect 21361 2567 21419 2573
rect 21361 2564 21373 2567
rect 20956 2536 21373 2564
rect 20956 2524 20962 2536
rect 21361 2533 21373 2536
rect 21407 2533 21419 2567
rect 21361 2527 21419 2533
rect 23290 2524 23296 2576
rect 23348 2564 23354 2576
rect 23934 2564 23940 2576
rect 23348 2536 23940 2564
rect 23348 2524 23354 2536
rect 23934 2524 23940 2536
rect 23992 2564 23998 2576
rect 24228 2573 24256 2604
rect 24121 2567 24179 2573
rect 24121 2564 24133 2567
rect 23992 2536 24133 2564
rect 23992 2524 23998 2536
rect 24121 2533 24133 2536
rect 24167 2533 24179 2567
rect 24121 2527 24179 2533
rect 24213 2567 24271 2573
rect 24213 2533 24225 2567
rect 24259 2533 24271 2567
rect 24213 2527 24271 2533
rect 24765 2567 24823 2573
rect 24765 2533 24777 2567
rect 24811 2564 24823 2567
rect 25222 2564 25228 2576
rect 24811 2536 25228 2564
rect 24811 2533 24823 2536
rect 24765 2527 24823 2533
rect 25222 2524 25228 2536
rect 25280 2524 25286 2576
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 16224 2468 17141 2496
rect 15197 2431 15255 2437
rect 15197 2428 15209 2431
rect 14792 2400 15209 2428
rect 14792 2388 14798 2400
rect 15197 2397 15209 2400
rect 15243 2397 15255 2431
rect 15562 2428 15568 2440
rect 15523 2400 15568 2428
rect 15197 2391 15255 2397
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 16224 2428 16252 2468
rect 17129 2465 17141 2468
rect 17175 2465 17187 2499
rect 17129 2459 17187 2465
rect 19426 2456 19432 2508
rect 19484 2496 19490 2508
rect 19613 2499 19671 2505
rect 19613 2496 19625 2499
rect 19484 2468 19625 2496
rect 19484 2456 19490 2468
rect 19613 2465 19625 2468
rect 19659 2465 19671 2499
rect 19613 2459 19671 2465
rect 22462 2456 22468 2508
rect 22520 2496 22526 2508
rect 22741 2499 22799 2505
rect 22741 2496 22753 2499
rect 22520 2468 22753 2496
rect 22520 2456 22526 2468
rect 22741 2465 22753 2468
rect 22787 2465 22799 2499
rect 22741 2459 22799 2465
rect 23477 2499 23535 2505
rect 23477 2465 23489 2499
rect 23523 2496 23535 2499
rect 23750 2496 23756 2508
rect 23523 2468 23756 2496
rect 23523 2465 23535 2468
rect 23477 2459 23535 2465
rect 23750 2456 23756 2468
rect 23808 2456 23814 2508
rect 24946 2456 24952 2508
rect 25004 2496 25010 2508
rect 25041 2499 25099 2505
rect 25041 2496 25053 2499
rect 25004 2468 25053 2496
rect 25004 2456 25010 2468
rect 25041 2465 25053 2468
rect 25087 2465 25099 2499
rect 25041 2459 25099 2465
rect 15672 2400 16252 2428
rect 14921 2363 14979 2369
rect 14921 2360 14933 2363
rect 13786 2332 14933 2360
rect 12345 2323 12403 2329
rect 14921 2329 14933 2332
rect 14967 2360 14979 2363
rect 15672 2360 15700 2400
rect 18414 2388 18420 2440
rect 18472 2428 18478 2440
rect 18693 2431 18751 2437
rect 18693 2428 18705 2431
rect 18472 2400 18705 2428
rect 18472 2388 18478 2400
rect 18693 2397 18705 2400
rect 18739 2428 18751 2431
rect 19981 2431 20039 2437
rect 19981 2428 19993 2431
rect 18739 2400 19993 2428
rect 18739 2397 18751 2400
rect 18693 2391 18751 2397
rect 19981 2397 19993 2400
rect 20027 2397 20039 2431
rect 19981 2391 20039 2397
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2397 21327 2431
rect 21542 2428 21548 2440
rect 21503 2400 21548 2428
rect 21269 2391 21327 2397
rect 14967 2332 15700 2360
rect 14967 2329 14979 2332
rect 14921 2323 14979 2329
rect 18874 2320 18880 2372
rect 18932 2360 18938 2372
rect 20533 2363 20591 2369
rect 20533 2360 20545 2363
rect 18932 2332 20545 2360
rect 18932 2320 18938 2332
rect 20533 2329 20545 2332
rect 20579 2360 20591 2363
rect 21284 2360 21312 2391
rect 21542 2388 21548 2400
rect 21600 2388 21606 2440
rect 22278 2388 22284 2440
rect 22336 2428 22342 2440
rect 25593 2431 25651 2437
rect 25593 2428 25605 2431
rect 22336 2400 23474 2428
rect 22336 2388 22342 2400
rect 20579 2332 21312 2360
rect 23446 2360 23474 2400
rect 24228 2400 25605 2428
rect 24228 2360 24256 2400
rect 25593 2397 25605 2400
rect 25639 2397 25651 2431
rect 25593 2391 25651 2397
rect 23446 2332 24256 2360
rect 20579 2329 20591 2332
rect 20533 2323 20591 2329
rect 11238 2292 11244 2304
rect 10336 2264 11244 2292
rect 4847 2261 4859 2264
rect 4801 2255 4859 2261
rect 11238 2252 11244 2264
rect 11296 2252 11302 2304
rect 11422 2252 11428 2304
rect 11480 2292 11486 2304
rect 13722 2292 13728 2304
rect 11480 2264 13728 2292
rect 11480 2252 11486 2264
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 14458 2292 14464 2304
rect 14419 2264 14464 2292
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 17586 2252 17592 2304
rect 17644 2292 17650 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17644 2264 17693 2292
rect 17644 2252 17650 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 18046 2292 18052 2304
rect 18007 2264 18052 2292
rect 17681 2255 17739 2261
rect 18046 2252 18052 2264
rect 18104 2252 18110 2304
rect 20898 2292 20904 2304
rect 20859 2264 20904 2292
rect 20898 2252 20904 2264
rect 20956 2252 20962 2304
rect 22462 2252 22468 2304
rect 22520 2292 22526 2304
rect 22557 2295 22615 2301
rect 22557 2292 22569 2295
rect 22520 2264 22569 2292
rect 22520 2252 22526 2264
rect 22557 2261 22569 2264
rect 22603 2261 22615 2295
rect 22557 2255 22615 2261
rect 22646 2252 22652 2304
rect 22704 2292 22710 2304
rect 22925 2295 22983 2301
rect 22925 2292 22937 2295
rect 22704 2264 22937 2292
rect 22704 2252 22710 2264
rect 22925 2261 22937 2264
rect 22971 2261 22983 2295
rect 22925 2255 22983 2261
rect 23934 2252 23940 2304
rect 23992 2292 23998 2304
rect 25409 2295 25467 2301
rect 25409 2292 25421 2295
rect 23992 2264 25421 2292
rect 23992 2252 23998 2264
rect 25409 2261 25421 2264
rect 25455 2261 25467 2295
rect 25409 2255 25467 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 10042 2048 10048 2100
rect 10100 2088 10106 2100
rect 18046 2088 18052 2100
rect 10100 2060 18052 2088
rect 10100 2048 10106 2060
rect 18046 2048 18052 2060
rect 18104 2048 18110 2100
rect 6270 1980 6276 2032
rect 6328 2020 6334 2032
rect 11974 2020 11980 2032
rect 6328 1992 11980 2020
rect 6328 1980 6334 1992
rect 11974 1980 11980 1992
rect 12032 1980 12038 2032
rect 15470 144 15476 196
rect 15528 184 15534 196
rect 15528 156 21956 184
rect 15528 144 15534 156
rect 21928 128 21956 156
rect 6914 76 6920 128
rect 6972 116 6978 128
rect 8294 116 8300 128
rect 6972 88 8300 116
rect 6972 76 6978 88
rect 8294 76 8300 88
rect 8352 76 8358 128
rect 9766 76 9772 128
rect 9824 116 9830 128
rect 9824 88 13814 116
rect 9824 76 9830 88
rect 13786 48 13814 88
rect 14458 76 14464 128
rect 14516 116 14522 128
rect 21082 116 21088 128
rect 14516 88 21088 116
rect 14516 76 14522 88
rect 21082 76 21088 88
rect 21140 76 21146 128
rect 21910 76 21916 128
rect 21968 76 21974 128
rect 22370 76 22376 128
rect 22428 116 22434 128
rect 24302 116 24308 128
rect 22428 88 24308 116
rect 22428 76 22434 88
rect 24302 76 24308 88
rect 24360 76 24366 128
rect 26234 76 26240 128
rect 26292 116 26298 128
rect 27522 116 27528 128
rect 26292 88 27528 116
rect 26292 76 26298 88
rect 27522 76 27528 88
rect 27580 76 27586 128
rect 15562 48 15568 60
rect 13786 20 15568 48
rect 15562 8 15568 20
rect 15620 48 15626 60
rect 19334 48 19340 60
rect 15620 20 19340 48
rect 15620 8 15626 20
rect 19334 8 19340 20
rect 19392 8 19398 60
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 24768 24395 24820 24404
rect 24768 24361 24777 24395
rect 24777 24361 24811 24395
rect 24811 24361 24820 24395
rect 24768 24352 24820 24361
rect 25136 24216 25188 24268
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 24952 23808 25004 23860
rect 25136 23851 25188 23860
rect 25136 23817 25145 23851
rect 25145 23817 25179 23851
rect 25179 23817 25188 23851
rect 25136 23808 25188 23817
rect 23664 23468 23716 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 27620 23264 27672 23316
rect 15568 23128 15620 23180
rect 18972 23171 19024 23180
rect 18972 23137 18981 23171
rect 18981 23137 19015 23171
rect 19015 23137 19024 23171
rect 18972 23128 19024 23137
rect 24676 23128 24728 23180
rect 20904 23060 20956 23112
rect 23296 22924 23348 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 15568 22380 15620 22432
rect 18328 22380 18380 22432
rect 18972 22380 19024 22432
rect 24584 22423 24636 22432
rect 24584 22389 24593 22423
rect 24593 22389 24627 22423
rect 24627 22389 24636 22423
rect 24584 22380 24636 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 24860 21632 24912 21684
rect 25320 21292 25372 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 24768 21131 24820 21140
rect 24768 21097 24777 21131
rect 24777 21097 24811 21131
rect 24811 21097 24820 21131
rect 24768 21088 24820 21097
rect 24676 20952 24728 21004
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 24676 20476 24728 20528
rect 24952 20204 25004 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 24768 20043 24820 20052
rect 24768 20009 24777 20043
rect 24777 20009 24811 20043
rect 24811 20009 24820 20043
rect 24768 20000 24820 20009
rect 24676 19864 24728 19916
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 24676 19388 24728 19440
rect 24860 19159 24912 19168
rect 24860 19125 24869 19159
rect 24869 19125 24903 19159
rect 24903 19125 24912 19159
rect 24860 19116 24912 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 24768 18955 24820 18964
rect 24768 18921 24777 18955
rect 24777 18921 24811 18955
rect 24811 18921 24820 18955
rect 24768 18912 24820 18921
rect 23572 18819 23624 18828
rect 23572 18785 23581 18819
rect 23581 18785 23615 18819
rect 23615 18785 23624 18819
rect 23572 18776 23624 18785
rect 24676 18776 24728 18828
rect 23756 18708 23808 18760
rect 25228 18572 25280 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 24676 18368 24728 18420
rect 24124 18300 24176 18352
rect 23940 18164 23992 18216
rect 24216 18164 24268 18216
rect 22100 18028 22152 18080
rect 23572 18028 23624 18080
rect 25504 18028 25556 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 16396 17867 16448 17876
rect 16396 17833 16405 17867
rect 16405 17833 16439 17867
rect 16439 17833 16448 17867
rect 16396 17824 16448 17833
rect 16120 17731 16172 17740
rect 16120 17697 16129 17731
rect 16129 17697 16163 17731
rect 16163 17697 16172 17731
rect 16120 17688 16172 17697
rect 17776 17731 17828 17740
rect 17776 17697 17785 17731
rect 17785 17697 17819 17731
rect 17819 17697 17828 17731
rect 17776 17688 17828 17697
rect 21548 17731 21600 17740
rect 21548 17697 21557 17731
rect 21557 17697 21591 17731
rect 21591 17697 21600 17731
rect 21548 17688 21600 17697
rect 22836 17731 22888 17740
rect 22836 17697 22845 17731
rect 22845 17697 22879 17731
rect 22879 17697 22888 17731
rect 22836 17688 22888 17697
rect 25044 17688 25096 17740
rect 21824 17663 21876 17672
rect 21824 17629 21833 17663
rect 21833 17629 21867 17663
rect 21867 17629 21876 17663
rect 21824 17620 21876 17629
rect 23848 17620 23900 17672
rect 18144 17527 18196 17536
rect 18144 17493 18153 17527
rect 18153 17493 18187 17527
rect 18187 17493 18196 17527
rect 18144 17484 18196 17493
rect 23296 17484 23348 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 16120 17280 16172 17332
rect 17776 17323 17828 17332
rect 17776 17289 17785 17323
rect 17785 17289 17819 17323
rect 17819 17289 17828 17323
rect 17776 17280 17828 17289
rect 21548 17323 21600 17332
rect 21548 17289 21557 17323
rect 21557 17289 21591 17323
rect 21591 17289 21600 17323
rect 21548 17280 21600 17289
rect 21916 17280 21968 17332
rect 25044 17280 25096 17332
rect 25412 17323 25464 17332
rect 25412 17289 25421 17323
rect 25421 17289 25455 17323
rect 25455 17289 25464 17323
rect 25412 17280 25464 17289
rect 15476 17076 15528 17128
rect 17040 17076 17092 17128
rect 18972 17076 19024 17128
rect 20812 17076 20864 17128
rect 22008 17076 22060 17128
rect 23204 17076 23256 17128
rect 25228 17119 25280 17128
rect 25228 17085 25237 17119
rect 25237 17085 25271 17119
rect 25271 17085 25280 17119
rect 25228 17076 25280 17085
rect 16396 17051 16448 17060
rect 16396 17017 16405 17051
rect 16405 17017 16439 17051
rect 16439 17017 16448 17051
rect 16396 17008 16448 17017
rect 22744 17051 22796 17060
rect 22744 17017 22753 17051
rect 22753 17017 22787 17051
rect 22787 17017 22796 17051
rect 22744 17008 22796 17017
rect 23480 17008 23532 17060
rect 15292 16983 15344 16992
rect 15292 16949 15301 16983
rect 15301 16949 15335 16983
rect 15335 16949 15344 16983
rect 15292 16940 15344 16949
rect 19064 16983 19116 16992
rect 19064 16949 19073 16983
rect 19073 16949 19107 16983
rect 19107 16949 19116 16983
rect 19064 16940 19116 16949
rect 20720 16983 20772 16992
rect 20720 16949 20729 16983
rect 20729 16949 20763 16983
rect 20763 16949 20772 16983
rect 20720 16940 20772 16949
rect 22192 16940 22244 16992
rect 22836 16940 22888 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 24216 16736 24268 16788
rect 16212 16668 16264 16720
rect 18144 16668 18196 16720
rect 19524 16600 19576 16652
rect 21640 16643 21692 16652
rect 21640 16609 21649 16643
rect 21649 16609 21683 16643
rect 21683 16609 21692 16643
rect 21640 16600 21692 16609
rect 22560 16600 22612 16652
rect 23388 16643 23440 16652
rect 23388 16609 23397 16643
rect 23397 16609 23431 16643
rect 23431 16609 23440 16643
rect 23388 16600 23440 16609
rect 25044 16643 25096 16652
rect 25044 16609 25053 16643
rect 25053 16609 25087 16643
rect 25087 16609 25096 16643
rect 25044 16600 25096 16609
rect 15660 16575 15712 16584
rect 15660 16541 15669 16575
rect 15669 16541 15703 16575
rect 15703 16541 15712 16575
rect 15660 16532 15712 16541
rect 18144 16575 18196 16584
rect 18144 16541 18153 16575
rect 18153 16541 18187 16575
rect 18187 16541 18196 16575
rect 18144 16532 18196 16541
rect 18328 16532 18380 16584
rect 22652 16532 22704 16584
rect 24124 16532 24176 16584
rect 16672 16464 16724 16516
rect 19248 16439 19300 16448
rect 19248 16405 19257 16439
rect 19257 16405 19291 16439
rect 19291 16405 19300 16439
rect 19248 16396 19300 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 15292 16192 15344 16244
rect 18236 16192 18288 16244
rect 19064 16235 19116 16244
rect 19064 16201 19073 16235
rect 19073 16201 19107 16235
rect 19107 16201 19116 16235
rect 19064 16192 19116 16201
rect 21548 16235 21600 16244
rect 21548 16201 21557 16235
rect 21557 16201 21591 16235
rect 21591 16201 21600 16235
rect 21548 16192 21600 16201
rect 21824 16235 21876 16244
rect 21824 16201 21833 16235
rect 21833 16201 21867 16235
rect 21867 16201 21876 16235
rect 21824 16192 21876 16201
rect 25320 16192 25372 16244
rect 16120 16056 16172 16108
rect 18144 16056 18196 16108
rect 19248 16099 19300 16108
rect 19248 16065 19257 16099
rect 19257 16065 19291 16099
rect 19291 16065 19300 16099
rect 19248 16056 19300 16065
rect 19524 16099 19576 16108
rect 19524 16065 19533 16099
rect 19533 16065 19567 16099
rect 19567 16065 19576 16099
rect 19524 16056 19576 16065
rect 22100 16099 22152 16108
rect 22100 16065 22109 16099
rect 22109 16065 22143 16099
rect 22143 16065 22152 16099
rect 22100 16056 22152 16065
rect 22468 16099 22520 16108
rect 22468 16065 22477 16099
rect 22477 16065 22511 16099
rect 22511 16065 22520 16099
rect 22468 16056 22520 16065
rect 21548 15988 21600 16040
rect 15384 15963 15436 15972
rect 15384 15929 15393 15963
rect 15393 15929 15427 15963
rect 15427 15929 15436 15963
rect 15384 15920 15436 15929
rect 16212 15895 16264 15904
rect 16212 15861 16221 15895
rect 16221 15861 16255 15895
rect 16255 15861 16264 15895
rect 16212 15852 16264 15861
rect 16672 15895 16724 15904
rect 16672 15861 16681 15895
rect 16681 15861 16715 15895
rect 16715 15861 16724 15895
rect 16672 15852 16724 15861
rect 19064 15852 19116 15904
rect 19432 15852 19484 15904
rect 21824 15852 21876 15904
rect 22928 15920 22980 15972
rect 24952 15920 25004 15972
rect 22284 15852 22336 15904
rect 23388 15895 23440 15904
rect 23388 15861 23397 15895
rect 23397 15861 23431 15895
rect 23431 15861 23440 15895
rect 23388 15852 23440 15861
rect 25044 15895 25096 15904
rect 25044 15861 25053 15895
rect 25053 15861 25087 15895
rect 25087 15861 25096 15895
rect 25044 15852 25096 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 18144 15648 18196 15700
rect 19432 15648 19484 15700
rect 21640 15691 21692 15700
rect 21640 15657 21649 15691
rect 21649 15657 21683 15691
rect 21683 15657 21692 15691
rect 21640 15648 21692 15657
rect 13820 15623 13872 15632
rect 13820 15589 13829 15623
rect 13829 15589 13863 15623
rect 13863 15589 13872 15623
rect 15476 15623 15528 15632
rect 13820 15580 13872 15589
rect 15476 15589 15485 15623
rect 15485 15589 15519 15623
rect 15519 15589 15528 15623
rect 15476 15580 15528 15589
rect 16120 15580 16172 15632
rect 17776 15580 17828 15632
rect 18328 15580 18380 15632
rect 18972 15580 19024 15632
rect 21916 15623 21968 15632
rect 21916 15589 21925 15623
rect 21925 15589 21959 15623
rect 21959 15589 21968 15623
rect 21916 15580 21968 15589
rect 22468 15623 22520 15632
rect 22468 15589 22477 15623
rect 22477 15589 22511 15623
rect 22511 15589 22520 15623
rect 22468 15580 22520 15589
rect 24216 15555 24268 15564
rect 24216 15521 24225 15555
rect 24225 15521 24259 15555
rect 24259 15521 24268 15555
rect 24216 15512 24268 15521
rect 13728 15487 13780 15496
rect 13728 15453 13737 15487
rect 13737 15453 13771 15487
rect 13771 15453 13780 15487
rect 13728 15444 13780 15453
rect 15660 15444 15712 15496
rect 17408 15487 17460 15496
rect 17408 15453 17417 15487
rect 17417 15453 17451 15487
rect 17451 15453 17460 15487
rect 17408 15444 17460 15453
rect 19432 15444 19484 15496
rect 21824 15487 21876 15496
rect 21824 15453 21833 15487
rect 21833 15453 21867 15487
rect 21867 15453 21876 15487
rect 21824 15444 21876 15453
rect 24768 15487 24820 15496
rect 24768 15453 24777 15487
rect 24777 15453 24811 15487
rect 24811 15453 24820 15487
rect 24768 15444 24820 15453
rect 19524 15419 19576 15428
rect 19524 15385 19533 15419
rect 19533 15385 19567 15419
rect 19567 15385 19576 15419
rect 19524 15376 19576 15385
rect 16488 15351 16540 15360
rect 16488 15317 16497 15351
rect 16497 15317 16531 15351
rect 16531 15317 16540 15351
rect 16488 15308 16540 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 13820 15147 13872 15156
rect 13820 15113 13829 15147
rect 13829 15113 13863 15147
rect 13863 15113 13872 15147
rect 13820 15104 13872 15113
rect 15476 15104 15528 15156
rect 16396 15104 16448 15156
rect 17776 15104 17828 15156
rect 18972 15104 19024 15156
rect 20720 15104 20772 15156
rect 21916 15104 21968 15156
rect 23112 15147 23164 15156
rect 23112 15113 23121 15147
rect 23121 15113 23155 15147
rect 23155 15113 23164 15147
rect 23112 15104 23164 15113
rect 23664 15104 23716 15156
rect 24216 15104 24268 15156
rect 25780 15147 25832 15156
rect 25780 15113 25789 15147
rect 25789 15113 25823 15147
rect 25823 15113 25832 15147
rect 25780 15104 25832 15113
rect 24308 15036 24360 15088
rect 17408 14968 17460 15020
rect 19248 14968 19300 15020
rect 23756 15011 23808 15020
rect 23756 14977 23765 15011
rect 23765 14977 23799 15011
rect 23799 14977 23808 15011
rect 23756 14968 23808 14977
rect 13452 14943 13504 14952
rect 13452 14909 13461 14943
rect 13461 14909 13495 14943
rect 13495 14909 13504 14943
rect 13452 14900 13504 14909
rect 14372 14943 14424 14952
rect 14372 14909 14381 14943
rect 14381 14909 14415 14943
rect 14415 14909 14424 14943
rect 14372 14900 14424 14909
rect 23112 14900 23164 14952
rect 25780 14900 25832 14952
rect 16488 14875 16540 14884
rect 16488 14841 16497 14875
rect 16497 14841 16531 14875
rect 16531 14841 16540 14875
rect 16488 14832 16540 14841
rect 18144 14875 18196 14884
rect 14280 14807 14332 14816
rect 14280 14773 14289 14807
rect 14289 14773 14323 14807
rect 14323 14773 14332 14807
rect 14280 14764 14332 14773
rect 16396 14764 16448 14816
rect 18144 14841 18153 14875
rect 18153 14841 18187 14875
rect 18187 14841 18196 14875
rect 18144 14832 18196 14841
rect 17040 14764 17092 14816
rect 19432 14807 19484 14816
rect 19432 14773 19441 14807
rect 19441 14773 19475 14807
rect 19475 14773 19484 14807
rect 19432 14764 19484 14773
rect 20168 14807 20220 14816
rect 20168 14773 20177 14807
rect 20177 14773 20211 14807
rect 20211 14773 20220 14807
rect 20168 14764 20220 14773
rect 20720 14764 20772 14816
rect 21824 14832 21876 14884
rect 23388 14832 23440 14884
rect 23848 14875 23900 14884
rect 23848 14841 23857 14875
rect 23857 14841 23891 14875
rect 23891 14841 23900 14875
rect 23848 14832 23900 14841
rect 24584 14832 24636 14884
rect 24860 14832 24912 14884
rect 20996 14764 21048 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 13728 14560 13780 14612
rect 15660 14560 15712 14612
rect 17040 14603 17092 14612
rect 17040 14569 17049 14603
rect 17049 14569 17083 14603
rect 17083 14569 17092 14603
rect 17040 14560 17092 14569
rect 17408 14603 17460 14612
rect 17408 14569 17417 14603
rect 17417 14569 17451 14603
rect 17451 14569 17460 14603
rect 17408 14560 17460 14569
rect 18972 14560 19024 14612
rect 14280 14492 14332 14544
rect 16856 14492 16908 14544
rect 21916 14560 21968 14612
rect 23756 14603 23808 14612
rect 23756 14569 23765 14603
rect 23765 14569 23799 14603
rect 23799 14569 23808 14603
rect 23756 14560 23808 14569
rect 22836 14535 22888 14544
rect 6368 14467 6420 14476
rect 6368 14433 6377 14467
rect 6377 14433 6411 14467
rect 6411 14433 6420 14467
rect 6368 14424 6420 14433
rect 13084 14424 13136 14476
rect 13360 14424 13412 14476
rect 14096 14467 14148 14476
rect 14096 14433 14105 14467
rect 14105 14433 14139 14467
rect 14139 14433 14148 14467
rect 14096 14424 14148 14433
rect 20812 14424 20864 14476
rect 22836 14501 22845 14535
rect 22845 14501 22879 14535
rect 22879 14501 22888 14535
rect 22836 14492 22888 14501
rect 23388 14535 23440 14544
rect 23388 14501 23397 14535
rect 23397 14501 23431 14535
rect 23431 14501 23440 14535
rect 23388 14492 23440 14501
rect 25136 14492 25188 14544
rect 15936 14356 15988 14408
rect 16120 14399 16172 14408
rect 16120 14365 16129 14399
rect 16129 14365 16163 14399
rect 16163 14365 16172 14399
rect 16120 14356 16172 14365
rect 17868 14399 17920 14408
rect 17868 14365 17877 14399
rect 17877 14365 17911 14399
rect 17911 14365 17920 14399
rect 17868 14356 17920 14365
rect 20720 14356 20772 14408
rect 20904 14399 20956 14408
rect 20904 14365 20913 14399
rect 20913 14365 20947 14399
rect 20947 14365 20956 14399
rect 20904 14356 20956 14365
rect 23572 14356 23624 14408
rect 24032 14356 24084 14408
rect 24584 14399 24636 14408
rect 24584 14365 24593 14399
rect 24593 14365 24627 14399
rect 24627 14365 24636 14399
rect 24584 14356 24636 14365
rect 12624 14288 12676 14340
rect 14372 14220 14424 14272
rect 18880 14220 18932 14272
rect 21916 14220 21968 14272
rect 23756 14220 23808 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 13084 13948 13136 14000
rect 14096 14016 14148 14068
rect 15936 14016 15988 14068
rect 17868 14016 17920 14068
rect 19800 14016 19852 14068
rect 20812 14016 20864 14068
rect 25136 14016 25188 14068
rect 25780 14059 25832 14068
rect 25780 14025 25789 14059
rect 25789 14025 25823 14059
rect 25823 14025 25832 14059
rect 25780 14016 25832 14025
rect 13452 13948 13504 14000
rect 16212 13948 16264 14000
rect 16856 13991 16908 14000
rect 16856 13957 16865 13991
rect 16865 13957 16899 13991
rect 16899 13957 16908 13991
rect 16856 13948 16908 13957
rect 18788 13948 18840 14000
rect 19432 13948 19484 14000
rect 20536 13948 20588 14000
rect 21916 13948 21968 14000
rect 22836 13948 22888 14000
rect 12348 13812 12400 13864
rect 13728 13812 13780 13864
rect 13268 13744 13320 13796
rect 6368 13676 6420 13728
rect 13360 13676 13412 13728
rect 13820 13719 13872 13728
rect 13820 13685 13829 13719
rect 13829 13685 13863 13719
rect 13863 13685 13872 13719
rect 14280 13812 14332 13864
rect 18880 13880 18932 13932
rect 19156 13880 19208 13932
rect 21824 13880 21876 13932
rect 22008 13880 22060 13932
rect 15936 13812 15988 13864
rect 21916 13812 21968 13864
rect 23204 13880 23256 13932
rect 24032 13923 24084 13932
rect 24032 13889 24041 13923
rect 24041 13889 24075 13923
rect 24075 13889 24084 13923
rect 24032 13880 24084 13889
rect 16120 13719 16172 13728
rect 13820 13676 13872 13685
rect 16120 13685 16129 13719
rect 16129 13685 16163 13719
rect 16163 13685 16172 13719
rect 16120 13676 16172 13685
rect 18328 13676 18380 13728
rect 19800 13744 19852 13796
rect 21272 13719 21324 13728
rect 21272 13685 21281 13719
rect 21281 13685 21315 13719
rect 21315 13685 21324 13719
rect 21272 13676 21324 13685
rect 25780 13812 25832 13864
rect 23756 13787 23808 13796
rect 23756 13753 23765 13787
rect 23765 13753 23799 13787
rect 23799 13753 23808 13787
rect 23756 13744 23808 13753
rect 24308 13676 24360 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 16120 13472 16172 13524
rect 17776 13472 17828 13524
rect 14372 13447 14424 13456
rect 14372 13413 14381 13447
rect 14381 13413 14415 13447
rect 14415 13413 14424 13447
rect 14372 13404 14424 13413
rect 16856 13404 16908 13456
rect 12624 13379 12676 13388
rect 12624 13345 12633 13379
rect 12633 13345 12667 13379
rect 12667 13345 12676 13379
rect 12624 13336 12676 13345
rect 13912 13379 13964 13388
rect 13912 13345 13921 13379
rect 13921 13345 13955 13379
rect 13955 13345 13964 13379
rect 13912 13336 13964 13345
rect 14464 13336 14516 13388
rect 19248 13404 19300 13456
rect 22744 13404 22796 13456
rect 23204 13447 23256 13456
rect 23204 13413 23213 13447
rect 23213 13413 23247 13447
rect 23247 13413 23256 13447
rect 23204 13404 23256 13413
rect 24216 13447 24268 13456
rect 24216 13413 24225 13447
rect 24225 13413 24259 13447
rect 24259 13413 24268 13447
rect 24216 13404 24268 13413
rect 24860 13404 24912 13456
rect 20812 13336 20864 13388
rect 15384 13268 15436 13320
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 14556 13200 14608 13252
rect 18788 13268 18840 13320
rect 21640 13311 21692 13320
rect 21640 13277 21649 13311
rect 21649 13277 21683 13311
rect 21683 13277 21692 13311
rect 21640 13268 21692 13277
rect 22836 13268 22888 13320
rect 24124 13311 24176 13320
rect 20720 13200 20772 13252
rect 24124 13277 24133 13311
rect 24133 13277 24167 13311
rect 24167 13277 24176 13311
rect 24124 13268 24176 13277
rect 24676 13243 24728 13252
rect 24676 13209 24685 13243
rect 24685 13209 24719 13243
rect 24719 13209 24728 13243
rect 24676 13200 24728 13209
rect 13728 13132 13780 13184
rect 15844 13175 15896 13184
rect 15844 13141 15853 13175
rect 15853 13141 15887 13175
rect 15887 13141 15896 13175
rect 15844 13132 15896 13141
rect 18328 13175 18380 13184
rect 18328 13141 18337 13175
rect 18337 13141 18371 13175
rect 18371 13141 18380 13175
rect 18328 13132 18380 13141
rect 18420 13132 18472 13184
rect 20260 13132 20312 13184
rect 20904 13132 20956 13184
rect 23020 13132 23072 13184
rect 23572 13175 23624 13184
rect 23572 13141 23581 13175
rect 23581 13141 23615 13175
rect 23615 13141 23624 13175
rect 23572 13132 23624 13141
rect 23940 13175 23992 13184
rect 23940 13141 23949 13175
rect 23949 13141 23983 13175
rect 23983 13141 23992 13175
rect 23940 13132 23992 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 12624 12928 12676 12980
rect 18328 12928 18380 12980
rect 19248 12971 19300 12980
rect 19248 12937 19257 12971
rect 19257 12937 19291 12971
rect 19291 12937 19300 12971
rect 19248 12928 19300 12937
rect 22008 12928 22060 12980
rect 22744 12928 22796 12980
rect 24860 12971 24912 12980
rect 24860 12937 24869 12971
rect 24869 12937 24903 12971
rect 24903 12937 24912 12971
rect 24860 12928 24912 12937
rect 12532 12860 12584 12912
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 14832 12792 14884 12844
rect 15568 12792 15620 12844
rect 16764 12835 16816 12844
rect 16764 12801 16773 12835
rect 16773 12801 16807 12835
rect 16807 12801 16816 12835
rect 16764 12792 16816 12801
rect 23756 12860 23808 12912
rect 18696 12792 18748 12844
rect 20536 12835 20588 12844
rect 12716 12724 12768 12776
rect 13268 12767 13320 12776
rect 13268 12733 13277 12767
rect 13277 12733 13311 12767
rect 13311 12733 13320 12767
rect 13268 12724 13320 12733
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 14464 12724 14516 12776
rect 16028 12724 16080 12776
rect 16672 12767 16724 12776
rect 16672 12733 16681 12767
rect 16681 12733 16715 12767
rect 16715 12733 16724 12767
rect 16672 12724 16724 12733
rect 14740 12699 14792 12708
rect 14740 12665 14749 12699
rect 14749 12665 14783 12699
rect 14783 12665 14792 12699
rect 14740 12656 14792 12665
rect 15844 12656 15896 12708
rect 13268 12588 13320 12640
rect 13912 12588 13964 12640
rect 14464 12631 14516 12640
rect 14464 12597 14473 12631
rect 14473 12597 14507 12631
rect 14507 12597 14516 12631
rect 14464 12588 14516 12597
rect 16028 12631 16080 12640
rect 16028 12597 16037 12631
rect 16037 12597 16071 12631
rect 16071 12597 16080 12631
rect 16028 12588 16080 12597
rect 19524 12588 19576 12640
rect 20260 12767 20312 12776
rect 20260 12733 20269 12767
rect 20269 12733 20303 12767
rect 20303 12733 20312 12767
rect 20260 12724 20312 12733
rect 20536 12801 20545 12835
rect 20545 12801 20579 12835
rect 20579 12801 20588 12835
rect 20536 12792 20588 12801
rect 21640 12792 21692 12844
rect 23940 12835 23992 12844
rect 23940 12801 23949 12835
rect 23949 12801 23983 12835
rect 23983 12801 23992 12835
rect 23940 12792 23992 12801
rect 24676 12792 24728 12844
rect 27620 12724 27672 12776
rect 22100 12656 22152 12708
rect 25044 12656 25096 12708
rect 20812 12631 20864 12640
rect 20812 12597 20821 12631
rect 20821 12597 20855 12631
rect 20855 12597 20864 12631
rect 20812 12588 20864 12597
rect 21272 12631 21324 12640
rect 21272 12597 21281 12631
rect 21281 12597 21315 12631
rect 21315 12597 21324 12631
rect 21272 12588 21324 12597
rect 22836 12588 22888 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 8300 12384 8352 12436
rect 13544 12384 13596 12436
rect 15292 12384 15344 12436
rect 16764 12427 16816 12436
rect 12532 12359 12584 12368
rect 12532 12325 12541 12359
rect 12541 12325 12575 12359
rect 12575 12325 12584 12359
rect 12532 12316 12584 12325
rect 16764 12393 16773 12427
rect 16773 12393 16807 12427
rect 16807 12393 16816 12427
rect 16764 12384 16816 12393
rect 18696 12427 18748 12436
rect 18696 12393 18705 12427
rect 18705 12393 18739 12427
rect 18739 12393 18748 12427
rect 18696 12384 18748 12393
rect 20260 12384 20312 12436
rect 22100 12427 22152 12436
rect 22100 12393 22109 12427
rect 22109 12393 22143 12427
rect 22143 12393 22152 12427
rect 22100 12384 22152 12393
rect 23020 12427 23072 12436
rect 23020 12393 23029 12427
rect 23029 12393 23063 12427
rect 23063 12393 23072 12427
rect 23020 12384 23072 12393
rect 24124 12427 24176 12436
rect 24124 12393 24133 12427
rect 24133 12393 24167 12427
rect 24167 12393 24176 12427
rect 24124 12384 24176 12393
rect 18420 12359 18472 12368
rect 18420 12325 18429 12359
rect 18429 12325 18463 12359
rect 18463 12325 18472 12359
rect 18420 12316 18472 12325
rect 7932 12291 7984 12300
rect 7932 12257 7941 12291
rect 7941 12257 7975 12291
rect 7975 12257 7984 12291
rect 7932 12248 7984 12257
rect 12348 12291 12400 12300
rect 11888 12180 11940 12232
rect 12348 12257 12357 12291
rect 12357 12257 12391 12291
rect 12391 12257 12400 12291
rect 12348 12248 12400 12257
rect 13268 12248 13320 12300
rect 13820 12291 13872 12300
rect 13820 12257 13829 12291
rect 13829 12257 13863 12291
rect 13863 12257 13872 12291
rect 13820 12248 13872 12257
rect 17224 12248 17276 12300
rect 20812 12316 20864 12368
rect 21272 12316 21324 12368
rect 21824 12316 21876 12368
rect 12624 12180 12676 12232
rect 14096 12223 14148 12232
rect 14096 12189 14105 12223
rect 14105 12189 14139 12223
rect 14139 12189 14148 12223
rect 14096 12180 14148 12189
rect 15384 12223 15436 12232
rect 15384 12189 15393 12223
rect 15393 12189 15427 12223
rect 15427 12189 15436 12223
rect 15384 12180 15436 12189
rect 15568 12180 15620 12232
rect 17868 12223 17920 12232
rect 17868 12189 17874 12223
rect 17874 12189 17920 12223
rect 17868 12180 17920 12189
rect 18052 12223 18104 12232
rect 18052 12189 18061 12223
rect 18061 12189 18095 12223
rect 18095 12189 18104 12223
rect 18052 12180 18104 12189
rect 23020 12291 23072 12300
rect 23020 12257 23029 12291
rect 23029 12257 23063 12291
rect 23063 12257 23072 12291
rect 23020 12248 23072 12257
rect 23204 12248 23256 12300
rect 24676 12291 24728 12300
rect 24676 12257 24685 12291
rect 24685 12257 24719 12291
rect 24719 12257 24728 12291
rect 24676 12248 24728 12257
rect 19984 12223 20036 12232
rect 18972 12112 19024 12164
rect 19984 12189 19993 12223
rect 19993 12189 20027 12223
rect 20027 12189 20036 12223
rect 19984 12180 20036 12189
rect 20260 12180 20312 12232
rect 20812 12112 20864 12164
rect 24676 12112 24728 12164
rect 14556 12087 14608 12096
rect 14556 12053 14565 12087
rect 14565 12053 14599 12087
rect 14599 12053 14608 12087
rect 14556 12044 14608 12053
rect 14832 12044 14884 12096
rect 15752 12044 15804 12096
rect 17960 12087 18012 12096
rect 17960 12053 17969 12087
rect 17969 12053 18003 12087
rect 18003 12053 18012 12087
rect 17960 12044 18012 12053
rect 19064 12087 19116 12096
rect 19064 12053 19073 12087
rect 19073 12053 19107 12087
rect 19107 12053 19116 12087
rect 19064 12044 19116 12053
rect 23204 12044 23256 12096
rect 25044 12044 25096 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 13820 11840 13872 11892
rect 15384 11840 15436 11892
rect 11980 11772 12032 11824
rect 14556 11772 14608 11824
rect 20996 11840 21048 11892
rect 22008 11883 22060 11892
rect 22008 11849 22017 11883
rect 22017 11849 22051 11883
rect 22051 11849 22060 11883
rect 22008 11840 22060 11849
rect 23388 11883 23440 11892
rect 23388 11849 23397 11883
rect 23397 11849 23431 11883
rect 23431 11849 23440 11883
rect 23388 11840 23440 11849
rect 24676 11883 24728 11892
rect 24676 11849 24685 11883
rect 24685 11849 24719 11883
rect 24719 11849 24728 11883
rect 24676 11840 24728 11849
rect 25044 11883 25096 11892
rect 25044 11849 25053 11883
rect 25053 11849 25087 11883
rect 25087 11849 25096 11883
rect 25044 11840 25096 11849
rect 25780 11883 25832 11892
rect 25780 11849 25789 11883
rect 25789 11849 25823 11883
rect 25823 11849 25832 11883
rect 25780 11840 25832 11849
rect 16856 11772 16908 11824
rect 23204 11772 23256 11824
rect 23572 11772 23624 11824
rect 13636 11704 13688 11756
rect 14832 11704 14884 11756
rect 18972 11747 19024 11756
rect 18972 11713 18981 11747
rect 18981 11713 19015 11747
rect 19015 11713 19024 11747
rect 18972 11704 19024 11713
rect 20260 11747 20312 11756
rect 20260 11713 20269 11747
rect 20269 11713 20303 11747
rect 20303 11713 20312 11747
rect 20260 11704 20312 11713
rect 23940 11704 23992 11756
rect 13452 11636 13504 11688
rect 14096 11636 14148 11688
rect 14556 11636 14608 11688
rect 12348 11568 12400 11620
rect 13544 11568 13596 11620
rect 15108 11568 15160 11620
rect 15752 11611 15804 11620
rect 15752 11577 15761 11611
rect 15761 11577 15795 11611
rect 15795 11577 15804 11611
rect 15752 11568 15804 11577
rect 17868 11568 17920 11620
rect 6920 11500 6972 11552
rect 7932 11500 7984 11552
rect 13268 11543 13320 11552
rect 13268 11509 13277 11543
rect 13277 11509 13311 11543
rect 13311 11509 13320 11543
rect 13268 11500 13320 11509
rect 13728 11543 13780 11552
rect 13728 11509 13737 11543
rect 13737 11509 13771 11543
rect 13771 11509 13780 11543
rect 13728 11500 13780 11509
rect 15292 11543 15344 11552
rect 15292 11509 15301 11543
rect 15301 11509 15335 11543
rect 15335 11509 15344 11543
rect 15292 11500 15344 11509
rect 17224 11500 17276 11552
rect 18052 11500 18104 11552
rect 19156 11636 19208 11688
rect 19524 11679 19576 11688
rect 19524 11645 19533 11679
rect 19533 11645 19567 11679
rect 19567 11645 19576 11679
rect 19524 11636 19576 11645
rect 21088 11679 21140 11688
rect 19064 11568 19116 11620
rect 21088 11645 21097 11679
rect 21097 11645 21131 11679
rect 21131 11645 21140 11679
rect 21088 11636 21140 11645
rect 25780 11636 25832 11688
rect 18788 11500 18840 11552
rect 19156 11500 19208 11552
rect 20628 11543 20680 11552
rect 20628 11509 20637 11543
rect 20637 11509 20671 11543
rect 20671 11509 20680 11543
rect 20628 11500 20680 11509
rect 21272 11568 21324 11620
rect 23756 11611 23808 11620
rect 23756 11577 23765 11611
rect 23765 11577 23799 11611
rect 23799 11577 23808 11611
rect 23756 11568 23808 11577
rect 23020 11500 23072 11552
rect 23388 11500 23440 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 12072 11296 12124 11348
rect 14556 11339 14608 11348
rect 12808 11228 12860 11280
rect 13728 11228 13780 11280
rect 14556 11305 14565 11339
rect 14565 11305 14599 11339
rect 14599 11305 14608 11339
rect 14556 11296 14608 11305
rect 15108 11339 15160 11348
rect 15108 11305 15117 11339
rect 15117 11305 15151 11339
rect 15151 11305 15160 11339
rect 15108 11296 15160 11305
rect 17040 11296 17092 11348
rect 16856 11271 16908 11280
rect 11888 11203 11940 11212
rect 11888 11169 11897 11203
rect 11897 11169 11931 11203
rect 11931 11169 11940 11203
rect 11888 11160 11940 11169
rect 15292 11160 15344 11212
rect 16856 11237 16865 11271
rect 16865 11237 16899 11271
rect 16899 11237 16908 11271
rect 16856 11228 16908 11237
rect 19984 11296 20036 11348
rect 21088 11296 21140 11348
rect 21180 11339 21232 11348
rect 21180 11305 21189 11339
rect 21189 11305 21223 11339
rect 21223 11305 21232 11339
rect 21180 11296 21232 11305
rect 19064 11228 19116 11280
rect 19156 11160 19208 11212
rect 19340 11160 19392 11212
rect 22008 11228 22060 11280
rect 20812 11160 20864 11212
rect 21456 11203 21508 11212
rect 21456 11169 21465 11203
rect 21465 11169 21499 11203
rect 21499 11169 21508 11203
rect 21456 11160 21508 11169
rect 25320 11228 25372 11280
rect 13176 10999 13228 11008
rect 13176 10965 13185 10999
rect 13185 10965 13219 10999
rect 13219 10965 13228 10999
rect 16212 11092 16264 11144
rect 13452 11024 13504 11076
rect 15752 11024 15804 11076
rect 16580 11092 16632 11144
rect 18052 11135 18104 11144
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 21088 11092 21140 11144
rect 23020 11092 23072 11144
rect 23572 11135 23624 11144
rect 23572 11101 23581 11135
rect 23581 11101 23615 11135
rect 23615 11101 23624 11135
rect 23572 11092 23624 11101
rect 23940 11135 23992 11144
rect 23940 11101 23949 11135
rect 23949 11101 23983 11135
rect 23983 11101 23992 11135
rect 23940 11092 23992 11101
rect 17960 11067 18012 11076
rect 17960 11033 17969 11067
rect 17969 11033 18003 11067
rect 18003 11033 18012 11067
rect 17960 11024 18012 11033
rect 15568 10999 15620 11008
rect 13176 10956 13228 10965
rect 15568 10965 15577 10999
rect 15577 10965 15611 10999
rect 15611 10965 15620 10999
rect 15568 10956 15620 10965
rect 16304 10999 16356 11008
rect 16304 10965 16328 10999
rect 16328 10965 16356 10999
rect 16304 10956 16356 10965
rect 17224 10999 17276 11008
rect 17224 10965 17233 10999
rect 17233 10965 17267 10999
rect 17267 10965 17276 10999
rect 17224 10956 17276 10965
rect 17868 10999 17920 11008
rect 17868 10965 17892 10999
rect 17892 10965 17920 10999
rect 17868 10956 17920 10965
rect 18328 10956 18380 11008
rect 23756 10956 23808 11008
rect 24676 10956 24728 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 11888 10795 11940 10804
rect 11888 10761 11897 10795
rect 11897 10761 11931 10795
rect 11931 10761 11940 10795
rect 11888 10752 11940 10761
rect 12532 10752 12584 10804
rect 12624 10727 12676 10736
rect 12624 10693 12633 10727
rect 12633 10693 12667 10727
rect 12667 10693 12676 10727
rect 12624 10684 12676 10693
rect 14832 10616 14884 10668
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 15292 10591 15344 10600
rect 15292 10557 15301 10591
rect 15301 10557 15335 10591
rect 15335 10557 15344 10591
rect 15292 10548 15344 10557
rect 16672 10752 16724 10804
rect 20812 10752 20864 10804
rect 21456 10752 21508 10804
rect 23020 10795 23072 10804
rect 23020 10761 23029 10795
rect 23029 10761 23063 10795
rect 23063 10761 23072 10795
rect 23020 10752 23072 10761
rect 25320 10752 25372 10804
rect 17960 10684 18012 10736
rect 18328 10727 18380 10736
rect 18328 10693 18337 10727
rect 18337 10693 18371 10727
rect 18371 10693 18380 10727
rect 18328 10684 18380 10693
rect 16672 10659 16724 10668
rect 16672 10625 16681 10659
rect 16681 10625 16715 10659
rect 16715 10625 16724 10659
rect 16672 10616 16724 10625
rect 17684 10616 17736 10668
rect 18052 10616 18104 10668
rect 22008 10684 22060 10736
rect 19340 10616 19392 10668
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 23480 10727 23532 10736
rect 23480 10693 23489 10727
rect 23489 10693 23523 10727
rect 23523 10693 23532 10727
rect 23480 10684 23532 10693
rect 23572 10684 23624 10736
rect 24676 10727 24728 10736
rect 24676 10693 24685 10727
rect 24685 10693 24719 10727
rect 24719 10693 24728 10727
rect 24676 10684 24728 10693
rect 24032 10659 24084 10668
rect 24032 10625 24041 10659
rect 24041 10625 24075 10659
rect 24075 10625 24084 10659
rect 24032 10616 24084 10625
rect 12992 10480 13044 10532
rect 13636 10523 13688 10532
rect 13636 10489 13645 10523
rect 13645 10489 13679 10523
rect 13679 10489 13688 10523
rect 13636 10480 13688 10489
rect 7564 10412 7616 10464
rect 7748 10455 7800 10464
rect 7748 10421 7757 10455
rect 7757 10421 7791 10455
rect 7791 10421 7800 10455
rect 7748 10412 7800 10421
rect 12256 10412 12308 10464
rect 12808 10412 12860 10464
rect 15936 10523 15988 10532
rect 15936 10489 15945 10523
rect 15945 10489 15979 10523
rect 15979 10489 15988 10523
rect 15936 10480 15988 10489
rect 17868 10548 17920 10600
rect 18696 10548 18748 10600
rect 23296 10548 23348 10600
rect 18052 10523 18104 10532
rect 15476 10455 15528 10464
rect 15476 10421 15485 10455
rect 15485 10421 15519 10455
rect 15519 10421 15528 10455
rect 15476 10412 15528 10421
rect 16212 10455 16264 10464
rect 16212 10421 16221 10455
rect 16221 10421 16255 10455
rect 16255 10421 16264 10455
rect 16212 10412 16264 10421
rect 17224 10412 17276 10464
rect 17684 10455 17736 10464
rect 17684 10421 17693 10455
rect 17693 10421 17727 10455
rect 17727 10421 17736 10455
rect 17684 10412 17736 10421
rect 18052 10489 18061 10523
rect 18061 10489 18095 10523
rect 18095 10489 18104 10523
rect 18052 10480 18104 10489
rect 19064 10480 19116 10532
rect 23480 10480 23532 10532
rect 18788 10412 18840 10464
rect 19156 10412 19208 10464
rect 20628 10412 20680 10464
rect 21272 10412 21324 10464
rect 25228 10455 25280 10464
rect 25228 10421 25237 10455
rect 25237 10421 25271 10455
rect 25271 10421 25280 10455
rect 25228 10412 25280 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 7564 10208 7616 10260
rect 12992 10208 13044 10260
rect 13176 10251 13228 10260
rect 13176 10217 13185 10251
rect 13185 10217 13219 10251
rect 13219 10217 13228 10251
rect 13176 10208 13228 10217
rect 14740 10208 14792 10260
rect 17224 10251 17276 10260
rect 17224 10217 17233 10251
rect 17233 10217 17267 10251
rect 17267 10217 17276 10251
rect 17224 10208 17276 10217
rect 18052 10208 18104 10260
rect 19340 10208 19392 10260
rect 21272 10251 21324 10260
rect 21272 10217 21281 10251
rect 21281 10217 21315 10251
rect 21315 10217 21324 10251
rect 21272 10208 21324 10217
rect 21732 10208 21784 10260
rect 23296 10208 23348 10260
rect 12072 10140 12124 10192
rect 12716 10140 12768 10192
rect 11796 10072 11848 10124
rect 12532 10072 12584 10124
rect 11888 10047 11940 10056
rect 11888 10013 11897 10047
rect 11897 10013 11931 10047
rect 11931 10013 11940 10047
rect 12808 10072 12860 10124
rect 13268 10140 13320 10192
rect 16028 10140 16080 10192
rect 16488 10140 16540 10192
rect 17040 10140 17092 10192
rect 24032 10183 24084 10192
rect 24032 10149 24041 10183
rect 24041 10149 24075 10183
rect 24075 10149 24084 10183
rect 24032 10140 24084 10149
rect 24952 10140 25004 10192
rect 13452 10072 13504 10124
rect 13820 10072 13872 10124
rect 16580 10072 16632 10124
rect 18696 10072 18748 10124
rect 19340 10115 19392 10124
rect 19340 10081 19349 10115
rect 19349 10081 19383 10115
rect 19383 10081 19392 10115
rect 19340 10072 19392 10081
rect 11888 10004 11940 10013
rect 12808 9936 12860 9988
rect 14832 10004 14884 10056
rect 15568 10047 15620 10056
rect 15568 10013 15577 10047
rect 15577 10013 15611 10047
rect 15611 10013 15620 10047
rect 15568 10004 15620 10013
rect 16672 10004 16724 10056
rect 17684 10004 17736 10056
rect 19892 10004 19944 10056
rect 21180 10004 21232 10056
rect 23388 10047 23440 10056
rect 23388 10013 23397 10047
rect 23397 10013 23431 10047
rect 23431 10013 23440 10047
rect 23388 10004 23440 10013
rect 25228 10004 25280 10056
rect 26056 10004 26108 10056
rect 16304 9936 16356 9988
rect 17868 9936 17920 9988
rect 25504 9979 25556 9988
rect 25504 9945 25513 9979
rect 25513 9945 25547 9979
rect 25547 9945 25556 9979
rect 25504 9936 25556 9945
rect 10876 9911 10928 9920
rect 10876 9877 10885 9911
rect 10885 9877 10919 9911
rect 10919 9877 10928 9911
rect 10876 9868 10928 9877
rect 11704 9868 11756 9920
rect 12716 9868 12768 9920
rect 14280 9868 14332 9920
rect 14556 9868 14608 9920
rect 15292 9868 15344 9920
rect 16396 9868 16448 9920
rect 17408 9868 17460 9920
rect 18328 9868 18380 9920
rect 18420 9868 18472 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 11796 9707 11848 9716
rect 11796 9673 11805 9707
rect 11805 9673 11839 9707
rect 11839 9673 11848 9707
rect 11796 9664 11848 9673
rect 12716 9707 12768 9716
rect 12716 9673 12725 9707
rect 12725 9673 12759 9707
rect 12759 9673 12768 9707
rect 12716 9664 12768 9673
rect 13452 9664 13504 9716
rect 14280 9664 14332 9716
rect 16580 9707 16632 9716
rect 16580 9673 16589 9707
rect 16589 9673 16623 9707
rect 16623 9673 16632 9707
rect 16580 9664 16632 9673
rect 17040 9707 17092 9716
rect 17040 9673 17049 9707
rect 17049 9673 17083 9707
rect 17083 9673 17092 9707
rect 17040 9664 17092 9673
rect 18328 9664 18380 9716
rect 21180 9664 21232 9716
rect 23296 9664 23348 9716
rect 24952 9707 25004 9716
rect 12992 9596 13044 9648
rect 8760 9528 8812 9580
rect 15752 9596 15804 9648
rect 16212 9596 16264 9648
rect 17408 9639 17460 9648
rect 17408 9605 17417 9639
rect 17417 9605 17451 9639
rect 17451 9605 17460 9639
rect 17408 9596 17460 9605
rect 22652 9596 22704 9648
rect 24952 9673 24961 9707
rect 24961 9673 24995 9707
rect 24995 9673 25004 9707
rect 24952 9664 25004 9673
rect 25780 9707 25832 9716
rect 25780 9673 25789 9707
rect 25789 9673 25823 9707
rect 25823 9673 25832 9707
rect 25780 9664 25832 9673
rect 26056 9707 26108 9716
rect 26056 9673 26065 9707
rect 26065 9673 26099 9707
rect 26099 9673 26108 9707
rect 26056 9664 26108 9673
rect 23848 9596 23900 9648
rect 14372 9571 14424 9580
rect 14372 9537 14381 9571
rect 14381 9537 14415 9571
rect 14415 9537 14424 9571
rect 14372 9528 14424 9537
rect 14648 9528 14700 9580
rect 19156 9528 19208 9580
rect 10876 9503 10928 9512
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 12716 9460 12768 9512
rect 12900 9503 12952 9512
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 10692 9392 10744 9444
rect 11520 9435 11572 9444
rect 11520 9401 11529 9435
rect 11529 9401 11563 9435
rect 11563 9401 11572 9435
rect 11520 9392 11572 9401
rect 11980 9392 12032 9444
rect 13268 9392 13320 9444
rect 14832 9460 14884 9512
rect 15384 9503 15436 9512
rect 15384 9469 15393 9503
rect 15393 9469 15427 9503
rect 15427 9469 15436 9503
rect 15384 9460 15436 9469
rect 15844 9460 15896 9512
rect 17684 9460 17736 9512
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 19340 9460 19392 9512
rect 23388 9528 23440 9580
rect 19892 9503 19944 9512
rect 19892 9469 19901 9503
rect 19901 9469 19935 9503
rect 19935 9469 19944 9503
rect 19892 9460 19944 9469
rect 21088 9460 21140 9512
rect 22560 9460 22612 9512
rect 23296 9460 23348 9512
rect 25780 9460 25832 9512
rect 13912 9435 13964 9444
rect 10048 9324 10100 9376
rect 11888 9324 11940 9376
rect 12072 9324 12124 9376
rect 13912 9401 13921 9435
rect 13921 9401 13955 9435
rect 13955 9401 13964 9435
rect 13912 9392 13964 9401
rect 15292 9392 15344 9444
rect 16304 9392 16356 9444
rect 23756 9435 23808 9444
rect 23756 9401 23765 9435
rect 23765 9401 23799 9435
rect 23799 9401 23808 9435
rect 23756 9392 23808 9401
rect 23848 9435 23900 9444
rect 23848 9401 23857 9435
rect 23857 9401 23891 9435
rect 23891 9401 23900 9435
rect 23848 9392 23900 9401
rect 14832 9324 14884 9376
rect 19248 9324 19300 9376
rect 21180 9324 21232 9376
rect 22928 9324 22980 9376
rect 23112 9324 23164 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 10692 9120 10744 9172
rect 11520 9052 11572 9104
rect 13728 9052 13780 9104
rect 13912 9052 13964 9104
rect 14740 9052 14792 9104
rect 18052 9120 18104 9172
rect 21088 9163 21140 9172
rect 21088 9129 21097 9163
rect 21097 9129 21131 9163
rect 21131 9129 21140 9163
rect 21088 9120 21140 9129
rect 22192 9163 22244 9172
rect 22192 9129 22201 9163
rect 22201 9129 22235 9163
rect 22235 9129 22244 9163
rect 22192 9120 22244 9129
rect 22928 9120 22980 9172
rect 17868 9095 17920 9104
rect 11980 9027 12032 9036
rect 9680 8848 9732 8900
rect 11980 8993 11989 9027
rect 11989 8993 12023 9027
rect 12023 8993 12032 9027
rect 11980 8984 12032 8993
rect 12348 9027 12400 9036
rect 12348 8993 12357 9027
rect 12357 8993 12391 9027
rect 12391 8993 12400 9027
rect 12348 8984 12400 8993
rect 12164 8916 12216 8968
rect 12532 8959 12584 8968
rect 12532 8925 12541 8959
rect 12541 8925 12575 8959
rect 12575 8925 12584 8959
rect 12532 8916 12584 8925
rect 13452 8959 13504 8968
rect 13452 8925 13461 8959
rect 13461 8925 13495 8959
rect 13495 8925 13504 8959
rect 13452 8916 13504 8925
rect 15292 8916 15344 8968
rect 16488 8984 16540 9036
rect 16948 8984 17000 9036
rect 17316 9027 17368 9036
rect 17316 8993 17325 9027
rect 17325 8993 17359 9027
rect 17359 8993 17368 9027
rect 17316 8984 17368 8993
rect 17868 9061 17877 9095
rect 17877 9061 17911 9095
rect 17911 9061 17920 9095
rect 17868 9052 17920 9061
rect 18420 8984 18472 9036
rect 18972 8984 19024 9036
rect 19984 9052 20036 9104
rect 21180 9052 21232 9104
rect 21732 9052 21784 9104
rect 23204 9095 23256 9104
rect 23204 9061 23213 9095
rect 23213 9061 23247 9095
rect 23247 9061 23256 9095
rect 23204 9052 23256 9061
rect 24860 9052 24912 9104
rect 25504 9052 25556 9104
rect 17592 8959 17644 8968
rect 17592 8925 17601 8959
rect 17601 8925 17635 8959
rect 17635 8925 17644 8959
rect 17592 8916 17644 8925
rect 21272 8959 21324 8968
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 23112 8959 23164 8968
rect 23112 8925 23121 8959
rect 23121 8925 23155 8959
rect 23155 8925 23164 8959
rect 23112 8916 23164 8925
rect 23388 8959 23440 8968
rect 23388 8925 23397 8959
rect 23397 8925 23431 8959
rect 23431 8925 23440 8959
rect 23388 8916 23440 8925
rect 24768 8916 24820 8968
rect 13176 8848 13228 8900
rect 14004 8891 14056 8900
rect 14004 8857 14013 8891
rect 14013 8857 14047 8891
rect 14047 8857 14056 8891
rect 14004 8848 14056 8857
rect 8944 8780 8996 8832
rect 11704 8780 11756 8832
rect 11796 8780 11848 8832
rect 13360 8780 13412 8832
rect 15476 8780 15528 8832
rect 18880 8823 18932 8832
rect 18880 8789 18889 8823
rect 18889 8789 18923 8823
rect 18923 8789 18932 8823
rect 18880 8780 18932 8789
rect 22560 8823 22612 8832
rect 22560 8789 22569 8823
rect 22569 8789 22603 8823
rect 22603 8789 22612 8823
rect 22560 8780 22612 8789
rect 23756 8780 23808 8832
rect 24032 8823 24084 8832
rect 24032 8789 24041 8823
rect 24041 8789 24075 8823
rect 24075 8789 24084 8823
rect 24032 8780 24084 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 9312 8619 9364 8628
rect 9312 8585 9321 8619
rect 9321 8585 9355 8619
rect 9355 8585 9364 8619
rect 9312 8576 9364 8585
rect 9680 8619 9732 8628
rect 9680 8585 9689 8619
rect 9689 8585 9723 8619
rect 9723 8585 9732 8619
rect 9680 8576 9732 8585
rect 9956 8619 10008 8628
rect 9956 8585 9965 8619
rect 9965 8585 9999 8619
rect 9999 8585 10008 8619
rect 9956 8576 10008 8585
rect 11980 8576 12032 8628
rect 12256 8619 12308 8628
rect 12256 8585 12265 8619
rect 12265 8585 12299 8619
rect 12299 8585 12308 8619
rect 12256 8576 12308 8585
rect 13452 8576 13504 8628
rect 13544 8508 13596 8560
rect 13728 8551 13780 8560
rect 13728 8517 13737 8551
rect 13737 8517 13771 8551
rect 13771 8517 13780 8551
rect 13728 8508 13780 8517
rect 9312 8372 9364 8424
rect 11796 8440 11848 8492
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 14464 8576 14516 8628
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 17316 8619 17368 8628
rect 17316 8585 17325 8619
rect 17325 8585 17359 8619
rect 17359 8585 17368 8619
rect 17316 8576 17368 8585
rect 19984 8576 20036 8628
rect 23204 8576 23256 8628
rect 23296 8576 23348 8628
rect 23848 8576 23900 8628
rect 24860 8576 24912 8628
rect 25780 8619 25832 8628
rect 25780 8585 25789 8619
rect 25789 8585 25823 8619
rect 25823 8585 25832 8619
rect 25780 8576 25832 8585
rect 15752 8551 15804 8560
rect 15752 8517 15761 8551
rect 15761 8517 15795 8551
rect 15795 8517 15804 8551
rect 15752 8508 15804 8517
rect 19432 8551 19484 8560
rect 19432 8517 19441 8551
rect 19441 8517 19475 8551
rect 19475 8517 19484 8551
rect 19432 8508 19484 8517
rect 23020 8508 23072 8560
rect 15476 8440 15528 8492
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 18880 8440 18932 8449
rect 20812 8440 20864 8492
rect 22560 8440 22612 8492
rect 25136 8440 25188 8492
rect 11336 8415 11388 8424
rect 9036 8304 9088 8356
rect 11336 8381 11345 8415
rect 11345 8381 11379 8415
rect 11379 8381 11388 8415
rect 11336 8372 11388 8381
rect 12164 8372 12216 8424
rect 10692 8304 10744 8356
rect 11520 8347 11572 8356
rect 11520 8313 11529 8347
rect 11529 8313 11563 8347
rect 11563 8313 11572 8347
rect 11520 8304 11572 8313
rect 12256 8304 12308 8356
rect 12716 8236 12768 8288
rect 13452 8279 13504 8288
rect 13452 8245 13461 8279
rect 13461 8245 13495 8279
rect 13495 8245 13504 8279
rect 13452 8236 13504 8245
rect 15292 8279 15344 8288
rect 15292 8245 15301 8279
rect 15301 8245 15335 8279
rect 15335 8245 15344 8279
rect 15292 8236 15344 8245
rect 15568 8304 15620 8356
rect 15844 8236 15896 8288
rect 25780 8372 25832 8424
rect 20536 8347 20588 8356
rect 20536 8313 20545 8347
rect 20545 8313 20579 8347
rect 20579 8313 20588 8347
rect 20536 8304 20588 8313
rect 20628 8347 20680 8356
rect 20628 8313 20637 8347
rect 20637 8313 20671 8347
rect 20671 8313 20680 8347
rect 20628 8304 20680 8313
rect 21180 8236 21232 8288
rect 21824 8279 21876 8288
rect 21824 8245 21833 8279
rect 21833 8245 21867 8279
rect 21867 8245 21876 8279
rect 22284 8304 22336 8356
rect 23756 8347 23808 8356
rect 23756 8313 23765 8347
rect 23765 8313 23799 8347
rect 23799 8313 23808 8347
rect 23756 8304 23808 8313
rect 23848 8347 23900 8356
rect 23848 8313 23857 8347
rect 23857 8313 23891 8347
rect 23891 8313 23900 8347
rect 24400 8347 24452 8356
rect 23848 8304 23900 8313
rect 24400 8313 24409 8347
rect 24409 8313 24443 8347
rect 24443 8313 24452 8347
rect 24400 8304 24452 8313
rect 24768 8304 24820 8356
rect 21824 8236 21876 8245
rect 23940 8236 23992 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 7840 8032 7892 8084
rect 12072 8032 12124 8084
rect 12256 8075 12308 8084
rect 12256 8041 12265 8075
rect 12265 8041 12299 8075
rect 12299 8041 12308 8075
rect 12256 8032 12308 8041
rect 12532 8032 12584 8084
rect 13176 8032 13228 8084
rect 18696 8032 18748 8084
rect 18788 8032 18840 8084
rect 20536 8075 20588 8084
rect 20536 8041 20545 8075
rect 20545 8041 20579 8075
rect 20579 8041 20588 8075
rect 20536 8032 20588 8041
rect 21272 8075 21324 8084
rect 21272 8041 21281 8075
rect 21281 8041 21315 8075
rect 21315 8041 21324 8075
rect 21272 8032 21324 8041
rect 23112 8075 23164 8084
rect 23112 8041 23121 8075
rect 23121 8041 23155 8075
rect 23155 8041 23164 8075
rect 23112 8032 23164 8041
rect 23756 8075 23808 8084
rect 23756 8041 23765 8075
rect 23765 8041 23799 8075
rect 23799 8041 23808 8075
rect 23756 8032 23808 8041
rect 13452 8007 13504 8016
rect 13452 7973 13461 8007
rect 13461 7973 13495 8007
rect 13495 7973 13504 8007
rect 13452 7964 13504 7973
rect 17868 7964 17920 8016
rect 18972 7964 19024 8016
rect 21180 7964 21232 8016
rect 24032 8007 24084 8016
rect 24032 7973 24041 8007
rect 24041 7973 24075 8007
rect 24075 7973 24084 8007
rect 24032 7964 24084 7973
rect 25136 7964 25188 8016
rect 7656 7896 7708 7948
rect 8852 7896 8904 7948
rect 10416 7939 10468 7948
rect 10416 7905 10425 7939
rect 10425 7905 10459 7939
rect 10459 7905 10468 7939
rect 10416 7896 10468 7905
rect 11520 7896 11572 7948
rect 15568 7896 15620 7948
rect 16212 7896 16264 7948
rect 17592 7896 17644 7948
rect 19156 7896 19208 7948
rect 19524 7896 19576 7948
rect 23664 7896 23716 7948
rect 25688 7896 25740 7948
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 14004 7871 14056 7880
rect 14004 7837 14013 7871
rect 14013 7837 14047 7871
rect 14047 7837 14056 7871
rect 14004 7828 14056 7837
rect 14832 7828 14884 7880
rect 16580 7828 16632 7880
rect 16856 7828 16908 7880
rect 21916 7828 21968 7880
rect 23940 7871 23992 7880
rect 23940 7837 23949 7871
rect 23949 7837 23983 7871
rect 23983 7837 23992 7871
rect 23940 7828 23992 7837
rect 24400 7871 24452 7880
rect 24400 7837 24409 7871
rect 24409 7837 24443 7871
rect 24443 7837 24452 7871
rect 24400 7828 24452 7837
rect 10416 7760 10468 7812
rect 12808 7803 12860 7812
rect 12808 7769 12817 7803
rect 12817 7769 12851 7803
rect 12851 7769 12860 7803
rect 12808 7760 12860 7769
rect 10140 7735 10192 7744
rect 10140 7701 10149 7735
rect 10149 7701 10183 7735
rect 10183 7701 10192 7735
rect 10140 7692 10192 7701
rect 10600 7735 10652 7744
rect 10600 7701 10609 7735
rect 10609 7701 10643 7735
rect 10643 7701 10652 7735
rect 10600 7692 10652 7701
rect 11336 7692 11388 7744
rect 12348 7692 12400 7744
rect 14556 7692 14608 7744
rect 15476 7692 15528 7744
rect 15660 7692 15712 7744
rect 15936 7692 15988 7744
rect 16212 7692 16264 7744
rect 16580 7692 16632 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 7656 7531 7708 7540
rect 7656 7497 7665 7531
rect 7665 7497 7699 7531
rect 7699 7497 7708 7531
rect 7656 7488 7708 7497
rect 8300 7531 8352 7540
rect 8300 7497 8309 7531
rect 8309 7497 8343 7531
rect 8343 7497 8352 7531
rect 8300 7488 8352 7497
rect 8944 7531 8996 7540
rect 8944 7497 8953 7531
rect 8953 7497 8987 7531
rect 8987 7497 8996 7531
rect 8944 7488 8996 7497
rect 10416 7488 10468 7540
rect 10600 7531 10652 7540
rect 10600 7497 10609 7531
rect 10609 7497 10643 7531
rect 10643 7497 10652 7531
rect 10600 7488 10652 7497
rect 10968 7488 11020 7540
rect 11704 7488 11756 7540
rect 10048 7420 10100 7472
rect 1676 7352 1728 7404
rect 10140 7352 10192 7404
rect 11336 7352 11388 7404
rect 13728 7420 13780 7472
rect 14832 7488 14884 7540
rect 15476 7488 15528 7540
rect 18696 7531 18748 7540
rect 18696 7497 18705 7531
rect 18705 7497 18739 7531
rect 18739 7497 18748 7531
rect 18696 7488 18748 7497
rect 19156 7531 19208 7540
rect 19156 7497 19165 7531
rect 19165 7497 19199 7531
rect 19199 7497 19208 7531
rect 19156 7488 19208 7497
rect 21180 7488 21232 7540
rect 22192 7488 22244 7540
rect 24032 7488 24084 7540
rect 25688 7488 25740 7540
rect 15108 7420 15160 7472
rect 15660 7420 15712 7472
rect 15752 7420 15804 7472
rect 14188 7352 14240 7404
rect 14556 7395 14608 7404
rect 14556 7361 14562 7395
rect 14562 7361 14608 7395
rect 14556 7352 14608 7361
rect 14832 7352 14884 7404
rect 15844 7395 15896 7404
rect 15844 7361 15853 7395
rect 15853 7361 15887 7395
rect 15887 7361 15896 7395
rect 15844 7352 15896 7361
rect 17316 7352 17368 7404
rect 19432 7352 19484 7404
rect 20812 7395 20864 7404
rect 20812 7361 20821 7395
rect 20821 7361 20855 7395
rect 20855 7361 20864 7395
rect 20812 7352 20864 7361
rect 22284 7352 22336 7404
rect 22376 7352 22428 7404
rect 24400 7395 24452 7404
rect 24400 7361 24409 7395
rect 24409 7361 24443 7395
rect 24443 7361 24452 7395
rect 24400 7352 24452 7361
rect 24860 7352 24912 7404
rect 8300 7284 8352 7336
rect 8944 7216 8996 7268
rect 9404 7284 9456 7336
rect 8852 7148 8904 7200
rect 9128 7148 9180 7200
rect 12256 7284 12308 7336
rect 14372 7327 14424 7336
rect 14372 7293 14381 7327
rect 14381 7293 14415 7327
rect 14415 7293 14424 7327
rect 14372 7284 14424 7293
rect 16580 7284 16632 7336
rect 17868 7284 17920 7336
rect 23664 7284 23716 7336
rect 10968 7259 11020 7268
rect 10968 7225 10977 7259
rect 10977 7225 11011 7259
rect 11011 7225 11020 7259
rect 10968 7216 11020 7225
rect 12808 7259 12860 7268
rect 12808 7225 12817 7259
rect 12817 7225 12851 7259
rect 12851 7225 12860 7259
rect 12808 7216 12860 7225
rect 16396 7216 16448 7268
rect 18880 7216 18932 7268
rect 22100 7216 22152 7268
rect 22744 7259 22796 7268
rect 22744 7225 22753 7259
rect 22753 7225 22787 7259
rect 22787 7225 22796 7259
rect 22744 7216 22796 7225
rect 14280 7148 14332 7200
rect 15844 7148 15896 7200
rect 16212 7148 16264 7200
rect 17776 7148 17828 7200
rect 19524 7148 19576 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 6828 6987 6880 6996
rect 6828 6953 6837 6987
rect 6837 6953 6871 6987
rect 6871 6953 6880 6987
rect 6828 6944 6880 6953
rect 8760 6987 8812 6996
rect 8760 6953 8769 6987
rect 8769 6953 8803 6987
rect 8803 6953 8812 6987
rect 8760 6944 8812 6953
rect 11520 6944 11572 6996
rect 11888 6944 11940 6996
rect 12256 6944 12308 6996
rect 12808 6944 12860 6996
rect 13176 6987 13228 6996
rect 13176 6953 13185 6987
rect 13185 6953 13219 6987
rect 13219 6953 13228 6987
rect 13176 6944 13228 6953
rect 14372 6987 14424 6996
rect 14372 6953 14381 6987
rect 14381 6953 14415 6987
rect 14415 6953 14424 6987
rect 14372 6944 14424 6953
rect 15108 6987 15160 6996
rect 15108 6953 15117 6987
rect 15117 6953 15151 6987
rect 15151 6953 15160 6987
rect 15108 6944 15160 6953
rect 15752 6944 15804 6996
rect 17316 6987 17368 6996
rect 17316 6953 17325 6987
rect 17325 6953 17359 6987
rect 17359 6953 17368 6987
rect 17316 6944 17368 6953
rect 17592 6944 17644 6996
rect 21180 6944 21232 6996
rect 23940 6987 23992 6996
rect 23940 6953 23949 6987
rect 23949 6953 23983 6987
rect 23983 6953 23992 6987
rect 23940 6944 23992 6953
rect 24400 6987 24452 6996
rect 24400 6953 24409 6987
rect 24409 6953 24443 6987
rect 24443 6953 24452 6987
rect 24400 6944 24452 6953
rect 11336 6876 11388 6928
rect 13820 6876 13872 6928
rect 6644 6808 6696 6860
rect 7564 6808 7616 6860
rect 8116 6808 8168 6860
rect 8300 6808 8352 6860
rect 9128 6851 9180 6860
rect 9128 6817 9137 6851
rect 9137 6817 9171 6851
rect 9171 6817 9180 6851
rect 9128 6808 9180 6817
rect 10140 6851 10192 6860
rect 10140 6817 10149 6851
rect 10149 6817 10183 6851
rect 10183 6817 10192 6851
rect 10140 6808 10192 6817
rect 12164 6808 12216 6860
rect 13360 6851 13412 6860
rect 13360 6817 13369 6851
rect 13369 6817 13403 6851
rect 13403 6817 13412 6851
rect 13360 6808 13412 6817
rect 11060 6740 11112 6792
rect 12532 6740 12584 6792
rect 14832 6808 14884 6860
rect 15292 6851 15344 6860
rect 15292 6817 15301 6851
rect 15301 6817 15335 6851
rect 15335 6817 15344 6851
rect 15292 6808 15344 6817
rect 16764 6808 16816 6860
rect 23112 6919 23164 6928
rect 23112 6885 23121 6919
rect 23121 6885 23155 6919
rect 23155 6885 23164 6919
rect 23112 6876 23164 6885
rect 24676 6919 24728 6928
rect 24676 6885 24685 6919
rect 24685 6885 24719 6919
rect 24719 6885 24728 6919
rect 24676 6876 24728 6885
rect 17868 6851 17920 6860
rect 17868 6817 17877 6851
rect 17877 6817 17911 6851
rect 17911 6817 17920 6851
rect 17868 6808 17920 6817
rect 19064 6851 19116 6860
rect 19064 6817 19073 6851
rect 19073 6817 19107 6851
rect 19107 6817 19116 6851
rect 19064 6808 19116 6817
rect 19248 6808 19300 6860
rect 19892 6851 19944 6860
rect 19892 6817 19901 6851
rect 19901 6817 19935 6851
rect 19935 6817 19944 6851
rect 19892 6808 19944 6817
rect 14280 6740 14332 6792
rect 9496 6715 9548 6724
rect 9496 6681 9505 6715
rect 9505 6681 9539 6715
rect 9539 6681 9548 6715
rect 9496 6672 9548 6681
rect 7104 6647 7156 6656
rect 7104 6613 7113 6647
rect 7113 6613 7147 6647
rect 7147 6613 7156 6647
rect 7104 6604 7156 6613
rect 8576 6604 8628 6656
rect 8852 6604 8904 6656
rect 15844 6740 15896 6792
rect 21916 6808 21968 6860
rect 20904 6783 20956 6792
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 23020 6783 23072 6792
rect 23020 6749 23029 6783
rect 23029 6749 23063 6783
rect 23063 6749 23072 6783
rect 23020 6740 23072 6749
rect 24216 6740 24268 6792
rect 24860 6783 24912 6792
rect 24860 6749 24869 6783
rect 24869 6749 24903 6783
rect 24903 6749 24912 6783
rect 24860 6740 24912 6749
rect 18696 6715 18748 6724
rect 18696 6681 18705 6715
rect 18705 6681 18739 6715
rect 18739 6681 18748 6715
rect 18696 6672 18748 6681
rect 23572 6715 23624 6724
rect 23572 6681 23581 6715
rect 23581 6681 23615 6715
rect 23615 6681 23624 6715
rect 23572 6672 23624 6681
rect 15476 6647 15528 6656
rect 15476 6613 15485 6647
rect 15485 6613 15519 6647
rect 15519 6613 15528 6647
rect 15476 6604 15528 6613
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 19984 6647 20036 6656
rect 19984 6613 19993 6647
rect 19993 6613 20027 6647
rect 20027 6613 20036 6647
rect 19984 6604 20036 6613
rect 21272 6604 21324 6656
rect 21824 6647 21876 6656
rect 21824 6613 21833 6647
rect 21833 6613 21867 6647
rect 21867 6613 21876 6647
rect 21824 6604 21876 6613
rect 22284 6604 22336 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 6644 6443 6696 6452
rect 6644 6409 6653 6443
rect 6653 6409 6687 6443
rect 6687 6409 6696 6443
rect 6644 6400 6696 6409
rect 7564 6443 7616 6452
rect 7564 6409 7573 6443
rect 7573 6409 7607 6443
rect 7607 6409 7616 6443
rect 7564 6400 7616 6409
rect 9496 6400 9548 6452
rect 10140 6443 10192 6452
rect 10140 6409 10149 6443
rect 10149 6409 10183 6443
rect 10183 6409 10192 6443
rect 10140 6400 10192 6409
rect 10968 6400 11020 6452
rect 11888 6443 11940 6452
rect 11888 6409 11897 6443
rect 11897 6409 11931 6443
rect 11931 6409 11940 6443
rect 11888 6400 11940 6409
rect 11980 6400 12032 6452
rect 13360 6400 13412 6452
rect 9312 6375 9364 6384
rect 9312 6341 9321 6375
rect 9321 6341 9355 6375
rect 9355 6341 9364 6375
rect 9312 6332 9364 6341
rect 13820 6332 13872 6384
rect 7104 6196 7156 6248
rect 8576 6264 8628 6316
rect 9404 6307 9456 6316
rect 9404 6273 9413 6307
rect 9413 6273 9447 6307
rect 9447 6273 9456 6307
rect 9404 6264 9456 6273
rect 10692 6264 10744 6316
rect 13176 6264 13228 6316
rect 10508 6196 10560 6248
rect 11980 6196 12032 6248
rect 12716 6196 12768 6248
rect 14280 6400 14332 6452
rect 14556 6400 14608 6452
rect 16120 6400 16172 6452
rect 16304 6443 16356 6452
rect 16304 6409 16313 6443
rect 16313 6409 16347 6443
rect 16347 6409 16356 6443
rect 16304 6400 16356 6409
rect 16764 6400 16816 6452
rect 24676 6443 24728 6452
rect 24676 6409 24685 6443
rect 24685 6409 24719 6443
rect 24719 6409 24728 6443
rect 24676 6400 24728 6409
rect 23112 6332 23164 6384
rect 15476 6264 15528 6316
rect 16396 6307 16448 6316
rect 16396 6273 16405 6307
rect 16405 6273 16439 6307
rect 16439 6273 16448 6307
rect 16396 6264 16448 6273
rect 19892 6307 19944 6316
rect 19892 6273 19901 6307
rect 19901 6273 19935 6307
rect 19935 6273 19944 6307
rect 19892 6264 19944 6273
rect 19984 6264 20036 6316
rect 24216 6332 24268 6384
rect 26792 6332 26844 6384
rect 9036 6171 9088 6180
rect 9036 6137 9045 6171
rect 9045 6137 9079 6171
rect 9079 6137 9088 6171
rect 9036 6128 9088 6137
rect 7380 6060 7432 6112
rect 8300 6060 8352 6112
rect 9680 6103 9732 6112
rect 9680 6069 9689 6103
rect 9689 6069 9723 6103
rect 9723 6069 9732 6103
rect 9680 6060 9732 6069
rect 10968 6103 11020 6112
rect 10968 6069 10977 6103
rect 10977 6069 11011 6103
rect 11011 6069 11020 6103
rect 10968 6060 11020 6069
rect 11520 6103 11572 6112
rect 11520 6069 11529 6103
rect 11529 6069 11563 6103
rect 11563 6069 11572 6103
rect 11520 6060 11572 6069
rect 12532 6103 12584 6112
rect 12532 6069 12541 6103
rect 12541 6069 12575 6103
rect 12575 6069 12584 6103
rect 12532 6060 12584 6069
rect 13176 6060 13228 6112
rect 15108 6196 15160 6248
rect 15936 6128 15988 6180
rect 19064 6196 19116 6248
rect 19524 6196 19576 6248
rect 20904 6196 20956 6248
rect 25228 6239 25280 6248
rect 25228 6205 25237 6239
rect 25237 6205 25271 6239
rect 25271 6205 25280 6239
rect 25228 6196 25280 6205
rect 14832 6060 14884 6112
rect 15844 6103 15896 6112
rect 15844 6069 15853 6103
rect 15853 6069 15887 6103
rect 15887 6069 15896 6103
rect 17132 6128 17184 6180
rect 17776 6128 17828 6180
rect 21180 6128 21232 6180
rect 23664 6171 23716 6180
rect 23664 6137 23673 6171
rect 23673 6137 23707 6171
rect 23707 6137 23716 6171
rect 23664 6128 23716 6137
rect 15844 6060 15896 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 9036 5899 9088 5908
rect 9036 5865 9045 5899
rect 9045 5865 9079 5899
rect 9079 5865 9088 5899
rect 9036 5856 9088 5865
rect 9404 5899 9456 5908
rect 9404 5865 9413 5899
rect 9413 5865 9447 5899
rect 9447 5865 9456 5899
rect 9404 5856 9456 5865
rect 10692 5899 10744 5908
rect 10692 5865 10701 5899
rect 10701 5865 10735 5899
rect 10735 5865 10744 5899
rect 10692 5856 10744 5865
rect 12532 5856 12584 5908
rect 13728 5899 13780 5908
rect 13728 5865 13737 5899
rect 13737 5865 13771 5899
rect 13771 5865 13780 5899
rect 13728 5856 13780 5865
rect 15108 5899 15160 5908
rect 15108 5865 15117 5899
rect 15117 5865 15151 5899
rect 15151 5865 15160 5899
rect 15108 5856 15160 5865
rect 16304 5856 16356 5908
rect 20904 5856 20956 5908
rect 23020 5899 23072 5908
rect 23020 5865 23029 5899
rect 23029 5865 23063 5899
rect 23063 5865 23072 5899
rect 23020 5856 23072 5865
rect 11152 5831 11204 5840
rect 11152 5797 11161 5831
rect 11161 5797 11195 5831
rect 11195 5797 11204 5831
rect 11152 5788 11204 5797
rect 11520 5788 11572 5840
rect 12716 5788 12768 5840
rect 12808 5831 12860 5840
rect 12808 5797 12817 5831
rect 12817 5797 12851 5831
rect 12851 5797 12860 5831
rect 18420 5831 18472 5840
rect 12808 5788 12860 5797
rect 18420 5797 18429 5831
rect 18429 5797 18463 5831
rect 18463 5797 18472 5831
rect 18420 5788 18472 5797
rect 6644 5720 6696 5772
rect 7288 5720 7340 5772
rect 8484 5720 8536 5772
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 10784 5720 10836 5772
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 6184 5652 6236 5704
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 9036 5652 9088 5704
rect 11244 5652 11296 5704
rect 12716 5695 12768 5704
rect 12716 5661 12725 5695
rect 12725 5661 12759 5695
rect 12759 5661 12768 5695
rect 12716 5652 12768 5661
rect 7472 5584 7524 5636
rect 9220 5584 9272 5636
rect 12440 5584 12492 5636
rect 7656 5559 7708 5568
rect 7656 5525 7665 5559
rect 7665 5525 7699 5559
rect 7699 5525 7708 5559
rect 7656 5516 7708 5525
rect 8300 5559 8352 5568
rect 8300 5525 8309 5559
rect 8309 5525 8343 5559
rect 8343 5525 8352 5559
rect 8300 5516 8352 5525
rect 8668 5559 8720 5568
rect 8668 5525 8677 5559
rect 8677 5525 8711 5559
rect 8711 5525 8720 5559
rect 8668 5516 8720 5525
rect 11612 5516 11664 5568
rect 15660 5652 15712 5704
rect 18328 5720 18380 5772
rect 17316 5652 17368 5704
rect 18512 5652 18564 5704
rect 19156 5652 19208 5704
rect 17040 5584 17092 5636
rect 14280 5516 14332 5568
rect 14648 5559 14700 5568
rect 14648 5525 14657 5559
rect 14657 5525 14691 5559
rect 14691 5525 14700 5559
rect 14648 5516 14700 5525
rect 15476 5559 15528 5568
rect 15476 5525 15485 5559
rect 15485 5525 15519 5559
rect 15519 5525 15528 5559
rect 15476 5516 15528 5525
rect 17868 5559 17920 5568
rect 17868 5525 17877 5559
rect 17877 5525 17911 5559
rect 17911 5525 17920 5559
rect 17868 5516 17920 5525
rect 18788 5584 18840 5636
rect 19524 5720 19576 5772
rect 20628 5788 20680 5840
rect 23664 5788 23716 5840
rect 25044 5831 25096 5840
rect 25044 5797 25053 5831
rect 25053 5797 25087 5831
rect 25087 5797 25096 5831
rect 25044 5788 25096 5797
rect 20076 5720 20128 5772
rect 21272 5720 21324 5772
rect 23388 5695 23440 5704
rect 23388 5661 23397 5695
rect 23397 5661 23431 5695
rect 23431 5661 23440 5695
rect 23388 5652 23440 5661
rect 23572 5652 23624 5704
rect 24952 5695 25004 5704
rect 24952 5661 24961 5695
rect 24961 5661 24995 5695
rect 24995 5661 25004 5695
rect 24952 5652 25004 5661
rect 20260 5584 20312 5636
rect 22744 5584 22796 5636
rect 19156 5516 19208 5568
rect 19984 5559 20036 5568
rect 19984 5525 19993 5559
rect 19993 5525 20027 5559
rect 20027 5525 20036 5559
rect 19984 5516 20036 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 6000 5312 6052 5364
rect 6644 5355 6696 5364
rect 6644 5321 6653 5355
rect 6653 5321 6687 5355
rect 6687 5321 6696 5355
rect 6644 5312 6696 5321
rect 7012 5312 7064 5364
rect 7288 5312 7340 5364
rect 7472 5355 7524 5364
rect 7472 5321 7481 5355
rect 7481 5321 7515 5355
rect 7515 5321 7524 5355
rect 7472 5312 7524 5321
rect 8392 5355 8444 5364
rect 8392 5321 8401 5355
rect 8401 5321 8435 5355
rect 8435 5321 8444 5355
rect 8392 5312 8444 5321
rect 10692 5312 10744 5364
rect 11520 5312 11572 5364
rect 12164 5355 12216 5364
rect 12164 5321 12173 5355
rect 12173 5321 12207 5355
rect 12207 5321 12216 5355
rect 12164 5312 12216 5321
rect 12808 5312 12860 5364
rect 15384 5312 15436 5364
rect 15660 5355 15712 5364
rect 15660 5321 15669 5355
rect 15669 5321 15703 5355
rect 15703 5321 15712 5355
rect 15660 5312 15712 5321
rect 16120 5312 16172 5364
rect 17316 5355 17368 5364
rect 17316 5321 17325 5355
rect 17325 5321 17359 5355
rect 17359 5321 17368 5355
rect 17316 5312 17368 5321
rect 18328 5312 18380 5364
rect 21272 5355 21324 5364
rect 10048 5287 10100 5296
rect 10048 5253 10057 5287
rect 10057 5253 10091 5287
rect 10091 5253 10100 5287
rect 10048 5244 10100 5253
rect 10784 5244 10836 5296
rect 11152 5244 11204 5296
rect 14648 5244 14700 5296
rect 8116 5176 8168 5228
rect 9956 5176 10008 5228
rect 11244 5176 11296 5228
rect 4988 4972 5040 5024
rect 7656 5151 7708 5160
rect 7656 5117 7674 5151
rect 7674 5117 7708 5151
rect 7656 5108 7708 5117
rect 8024 5108 8076 5160
rect 8852 5151 8904 5160
rect 8852 5117 8861 5151
rect 8861 5117 8895 5151
rect 8895 5117 8904 5151
rect 8852 5108 8904 5117
rect 9680 5108 9732 5160
rect 13176 5151 13228 5160
rect 13176 5117 13185 5151
rect 13185 5117 13219 5151
rect 13219 5117 13228 5151
rect 13176 5108 13228 5117
rect 14188 5176 14240 5228
rect 14740 5176 14792 5228
rect 15568 5176 15620 5228
rect 16028 5176 16080 5228
rect 9404 5040 9456 5092
rect 5356 4972 5408 5024
rect 6276 5015 6328 5024
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 7840 4972 7892 5024
rect 8208 4972 8260 5024
rect 9864 4972 9916 5024
rect 10968 5040 11020 5092
rect 15660 5108 15712 5160
rect 17684 5108 17736 5160
rect 21272 5321 21281 5355
rect 21281 5321 21315 5355
rect 21315 5321 21324 5355
rect 21272 5312 21324 5321
rect 21456 5312 21508 5364
rect 23664 5312 23716 5364
rect 25044 5312 25096 5364
rect 19984 5176 20036 5228
rect 21732 5219 21784 5228
rect 21732 5185 21741 5219
rect 21741 5185 21775 5219
rect 21775 5185 21784 5219
rect 21732 5176 21784 5185
rect 19156 5108 19208 5160
rect 20076 5151 20128 5160
rect 14648 5083 14700 5092
rect 14648 5049 14657 5083
rect 14657 5049 14691 5083
rect 14691 5049 14700 5083
rect 14648 5040 14700 5049
rect 15844 5040 15896 5092
rect 20076 5117 20085 5151
rect 20085 5117 20119 5151
rect 20119 5117 20128 5151
rect 20076 5108 20128 5117
rect 25136 5108 25188 5160
rect 14188 5015 14240 5024
rect 14188 4981 14197 5015
rect 14197 4981 14231 5015
rect 14231 4981 14240 5015
rect 14188 4972 14240 4981
rect 14556 4972 14608 5024
rect 16028 5015 16080 5024
rect 16028 4981 16037 5015
rect 16037 4981 16071 5015
rect 16071 4981 16080 5015
rect 16028 4972 16080 4981
rect 18144 4972 18196 5024
rect 21456 5040 21508 5092
rect 23756 5083 23808 5092
rect 23756 5049 23765 5083
rect 23765 5049 23799 5083
rect 23799 5049 23808 5083
rect 23756 5040 23808 5049
rect 19064 4972 19116 5024
rect 20168 5015 20220 5024
rect 20168 4981 20177 5015
rect 20177 4981 20211 5015
rect 20211 4981 20220 5015
rect 20168 4972 20220 4981
rect 22652 5015 22704 5024
rect 22652 4981 22661 5015
rect 22661 4981 22695 5015
rect 22695 4981 22704 5015
rect 22652 4972 22704 4981
rect 23572 4972 23624 5024
rect 24952 5040 25004 5092
rect 25688 4972 25740 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 5080 4768 5132 4820
rect 6092 4768 6144 4820
rect 8484 4768 8536 4820
rect 8852 4768 8904 4820
rect 5172 4632 5224 4684
rect 6184 4632 6236 4684
rect 7288 4632 7340 4684
rect 8300 4675 8352 4684
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 8484 4632 8536 4684
rect 9680 4768 9732 4820
rect 9956 4768 10008 4820
rect 12716 4768 12768 4820
rect 9864 4743 9916 4752
rect 9864 4709 9873 4743
rect 9873 4709 9907 4743
rect 9907 4709 9916 4743
rect 9864 4700 9916 4709
rect 11060 4700 11112 4752
rect 11796 4700 11848 4752
rect 12624 4700 12676 4752
rect 14648 4811 14700 4820
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 15292 4768 15344 4820
rect 18420 4768 18472 4820
rect 18696 4768 18748 4820
rect 21732 4811 21784 4820
rect 21732 4777 21741 4811
rect 21741 4777 21775 4811
rect 21775 4777 21784 4811
rect 21732 4768 21784 4777
rect 23388 4811 23440 4820
rect 23388 4777 23397 4811
rect 23397 4777 23431 4811
rect 23431 4777 23440 4811
rect 23388 4768 23440 4777
rect 23756 4811 23808 4820
rect 23756 4777 23765 4811
rect 23765 4777 23799 4811
rect 23799 4777 23808 4811
rect 23756 4768 23808 4777
rect 24952 4811 25004 4820
rect 14372 4700 14424 4752
rect 18972 4700 19024 4752
rect 21456 4700 21508 4752
rect 24124 4743 24176 4752
rect 24124 4709 24133 4743
rect 24133 4709 24167 4743
rect 24167 4709 24176 4743
rect 24124 4700 24176 4709
rect 24952 4777 24961 4811
rect 24961 4777 24995 4811
rect 24995 4777 25004 4811
rect 24952 4768 25004 4777
rect 10692 4632 10744 4684
rect 13452 4632 13504 4684
rect 8760 4607 8812 4616
rect 8760 4573 8769 4607
rect 8769 4573 8803 4607
rect 8803 4573 8812 4607
rect 8760 4564 8812 4573
rect 11612 4564 11664 4616
rect 8576 4496 8628 4548
rect 12440 4564 12492 4616
rect 12532 4564 12584 4616
rect 13176 4564 13228 4616
rect 14004 4632 14056 4684
rect 14556 4632 14608 4684
rect 15292 4675 15344 4684
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 15384 4632 15436 4684
rect 16120 4632 16172 4684
rect 17132 4632 17184 4684
rect 20628 4632 20680 4684
rect 14648 4564 14700 4616
rect 15660 4607 15712 4616
rect 15660 4573 15669 4607
rect 15669 4573 15703 4607
rect 15703 4573 15712 4607
rect 15660 4564 15712 4573
rect 18052 4607 18104 4616
rect 18052 4573 18061 4607
rect 18061 4573 18095 4607
rect 18095 4573 18104 4607
rect 18052 4564 18104 4573
rect 19156 4607 19208 4616
rect 19156 4573 19165 4607
rect 19165 4573 19199 4607
rect 19199 4573 19208 4607
rect 19156 4564 19208 4573
rect 7656 4428 7708 4480
rect 12440 4428 12492 4480
rect 12716 4471 12768 4480
rect 12716 4437 12725 4471
rect 12725 4437 12759 4471
rect 12759 4437 12768 4471
rect 12716 4428 12768 4437
rect 14740 4428 14792 4480
rect 16028 4496 16080 4548
rect 17040 4496 17092 4548
rect 18236 4496 18288 4548
rect 20168 4564 20220 4616
rect 22192 4564 22244 4616
rect 22468 4564 22520 4616
rect 23020 4564 23072 4616
rect 16212 4428 16264 4480
rect 17500 4428 17552 4480
rect 20076 4428 20128 4480
rect 22376 4496 22428 4548
rect 25044 4496 25096 4548
rect 21548 4428 21600 4480
rect 22468 4428 22520 4480
rect 23756 4428 23808 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 4160 4224 4212 4276
rect 12440 4224 12492 4276
rect 13452 4224 13504 4276
rect 15660 4224 15712 4276
rect 17040 4224 17092 4276
rect 17776 4267 17828 4276
rect 17776 4233 17785 4267
rect 17785 4233 17819 4267
rect 17819 4233 17828 4267
rect 17776 4224 17828 4233
rect 18972 4267 19024 4276
rect 18972 4233 18981 4267
rect 18981 4233 19015 4267
rect 19015 4233 19024 4267
rect 18972 4224 19024 4233
rect 22192 4224 22244 4276
rect 22652 4224 22704 4276
rect 23480 4224 23532 4276
rect 24124 4224 24176 4276
rect 2964 4199 3016 4208
rect 2964 4165 2973 4199
rect 2973 4165 3007 4199
rect 3007 4165 3016 4199
rect 2964 4156 3016 4165
rect 8116 4156 8168 4208
rect 8300 4156 8352 4208
rect 6276 4088 6328 4140
rect 7104 4088 7156 4140
rect 8484 4088 8536 4140
rect 10692 4156 10744 4208
rect 11796 4199 11848 4208
rect 11796 4165 11805 4199
rect 11805 4165 11839 4199
rect 11839 4165 11848 4199
rect 11796 4156 11848 4165
rect 23020 4199 23072 4208
rect 23020 4165 23029 4199
rect 23029 4165 23063 4199
rect 23063 4165 23072 4199
rect 23020 4156 23072 4165
rect 12532 4131 12584 4140
rect 12532 4097 12541 4131
rect 12541 4097 12575 4131
rect 12575 4097 12584 4131
rect 12532 4088 12584 4097
rect 18052 4131 18104 4140
rect 1435 4063 1487 4072
rect 1435 4029 1444 4063
rect 1444 4029 1478 4063
rect 1478 4029 1487 4063
rect 1435 4020 1487 4029
rect 1400 3884 1452 3936
rect 3240 3927 3292 3936
rect 3240 3893 3249 3927
rect 3249 3893 3283 3927
rect 3283 3893 3292 3927
rect 3240 3884 3292 3893
rect 4160 3884 4212 3936
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 8116 4063 8168 4072
rect 8116 4029 8125 4063
rect 8125 4029 8159 4063
rect 8159 4029 8168 4063
rect 8116 4020 8168 4029
rect 9128 4063 9180 4072
rect 9128 4029 9137 4063
rect 9137 4029 9171 4063
rect 9171 4029 9180 4063
rect 9128 4020 9180 4029
rect 9404 4020 9456 4072
rect 6276 3952 6328 4004
rect 9220 3952 9272 4004
rect 9956 3952 10008 4004
rect 11336 4063 11388 4072
rect 11336 4029 11345 4063
rect 11345 4029 11379 4063
rect 11379 4029 11388 4063
rect 11336 4020 11388 4029
rect 11520 4063 11572 4072
rect 11520 4029 11529 4063
rect 11529 4029 11563 4063
rect 11563 4029 11572 4063
rect 11520 4020 11572 4029
rect 12716 4020 12768 4072
rect 13360 3995 13412 4004
rect 13360 3961 13369 3995
rect 13369 3961 13403 3995
rect 13403 3961 13412 3995
rect 13360 3952 13412 3961
rect 14280 3995 14332 4004
rect 14280 3961 14289 3995
rect 14289 3961 14323 3995
rect 14323 3961 14332 3995
rect 14280 3952 14332 3961
rect 14924 3995 14976 4004
rect 4436 3884 4488 3936
rect 5172 3927 5224 3936
rect 5172 3893 5181 3927
rect 5181 3893 5215 3927
rect 5215 3893 5224 3927
rect 5172 3884 5224 3893
rect 6000 3884 6052 3936
rect 6184 3927 6236 3936
rect 6184 3893 6193 3927
rect 6193 3893 6227 3927
rect 6227 3893 6236 3927
rect 6184 3884 6236 3893
rect 7288 3884 7340 3936
rect 9588 3884 9640 3936
rect 9864 3884 9916 3936
rect 13912 3884 13964 3936
rect 14924 3961 14933 3995
rect 14933 3961 14967 3995
rect 14967 3961 14976 3995
rect 14924 3952 14976 3961
rect 14648 3884 14700 3936
rect 16028 4020 16080 4072
rect 16212 4063 16264 4072
rect 16212 4029 16221 4063
rect 16221 4029 16255 4063
rect 16255 4029 16264 4063
rect 16212 4020 16264 4029
rect 18052 4097 18061 4131
rect 18061 4097 18095 4131
rect 18095 4097 18104 4131
rect 18052 4088 18104 4097
rect 23388 4088 23440 4140
rect 24124 4088 24176 4140
rect 22192 4020 22244 4072
rect 24400 4020 24452 4072
rect 25044 4020 25096 4072
rect 16120 3952 16172 4004
rect 17776 3952 17828 4004
rect 21456 3952 21508 4004
rect 15844 3927 15896 3936
rect 15844 3893 15853 3927
rect 15853 3893 15887 3927
rect 15887 3893 15896 3927
rect 15844 3884 15896 3893
rect 16028 3884 16080 3936
rect 16304 3884 16356 3936
rect 19156 3884 19208 3936
rect 19524 3884 19576 3936
rect 20168 3884 20220 3936
rect 20720 3927 20772 3936
rect 20720 3893 20729 3927
rect 20729 3893 20763 3927
rect 20763 3893 20772 3927
rect 20720 3884 20772 3893
rect 21732 3927 21784 3936
rect 21732 3893 21741 3927
rect 21741 3893 21775 3927
rect 21775 3893 21784 3927
rect 21732 3884 21784 3893
rect 25412 3884 25464 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 6736 3723 6788 3732
rect 6736 3689 6745 3723
rect 6745 3689 6779 3723
rect 6779 3689 6788 3723
rect 6736 3680 6788 3689
rect 9680 3680 9732 3732
rect 10876 3680 10928 3732
rect 5264 3655 5316 3664
rect 5264 3621 5273 3655
rect 5273 3621 5307 3655
rect 5307 3621 5316 3655
rect 5264 3612 5316 3621
rect 8024 3612 8076 3664
rect 3056 3544 3108 3596
rect 5080 3544 5132 3596
rect 6644 3587 6696 3596
rect 6644 3553 6653 3587
rect 6653 3553 6687 3587
rect 6687 3553 6696 3587
rect 6644 3544 6696 3553
rect 8668 3587 8720 3596
rect 8668 3553 8677 3587
rect 8677 3553 8711 3587
rect 8711 3553 8720 3587
rect 8668 3544 8720 3553
rect 10140 3544 10192 3596
rect 5448 3519 5500 3528
rect 5448 3485 5457 3519
rect 5457 3485 5491 3519
rect 5491 3485 5500 3519
rect 5448 3476 5500 3485
rect 10692 3476 10744 3528
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 11152 3476 11204 3528
rect 11612 3680 11664 3732
rect 14004 3723 14056 3732
rect 14004 3689 14013 3723
rect 14013 3689 14047 3723
rect 14047 3689 14056 3723
rect 14004 3680 14056 3689
rect 14188 3680 14240 3732
rect 15292 3680 15344 3732
rect 17132 3723 17184 3732
rect 17132 3689 17141 3723
rect 17141 3689 17175 3723
rect 17175 3689 17184 3723
rect 17132 3680 17184 3689
rect 17776 3680 17828 3732
rect 20168 3680 20220 3732
rect 23572 3723 23624 3732
rect 12624 3612 12676 3664
rect 11888 3544 11940 3596
rect 14924 3612 14976 3664
rect 16028 3655 16080 3664
rect 16028 3621 16037 3655
rect 16037 3621 16071 3655
rect 16071 3621 16080 3655
rect 16028 3612 16080 3621
rect 18788 3612 18840 3664
rect 19340 3612 19392 3664
rect 20720 3612 20772 3664
rect 23572 3689 23581 3723
rect 23581 3689 23615 3723
rect 23615 3689 23624 3723
rect 23572 3680 23624 3689
rect 24400 3723 24452 3732
rect 24400 3689 24409 3723
rect 24409 3689 24443 3723
rect 24443 3689 24452 3723
rect 24400 3680 24452 3689
rect 24860 3680 24912 3732
rect 24952 3655 25004 3664
rect 24952 3621 24961 3655
rect 24961 3621 24995 3655
rect 24995 3621 25004 3655
rect 24952 3612 25004 3621
rect 16764 3544 16816 3596
rect 10876 3408 10928 3460
rect 12532 3408 12584 3460
rect 16028 3476 16080 3528
rect 16948 3476 17000 3528
rect 17592 3476 17644 3528
rect 23480 3587 23532 3596
rect 23480 3553 23489 3587
rect 23489 3553 23523 3587
rect 23523 3553 23532 3587
rect 23480 3544 23532 3553
rect 19524 3476 19576 3528
rect 20904 3519 20956 3528
rect 20904 3485 20913 3519
rect 20913 3485 20947 3519
rect 20947 3485 20956 3519
rect 20904 3476 20956 3485
rect 25228 3519 25280 3528
rect 25228 3485 25237 3519
rect 25237 3485 25271 3519
rect 25271 3485 25280 3519
rect 25228 3476 25280 3485
rect 18328 3408 18380 3460
rect 20076 3408 20128 3460
rect 23756 3408 23808 3460
rect 7472 3340 7524 3392
rect 8024 3340 8076 3392
rect 10968 3340 11020 3392
rect 12624 3340 12676 3392
rect 14648 3383 14700 3392
rect 14648 3349 14657 3383
rect 14657 3349 14691 3383
rect 14691 3349 14700 3383
rect 14648 3340 14700 3349
rect 15568 3340 15620 3392
rect 16212 3340 16264 3392
rect 17592 3340 17644 3392
rect 18420 3383 18472 3392
rect 18420 3349 18429 3383
rect 18429 3349 18463 3383
rect 18463 3349 18472 3383
rect 18420 3340 18472 3349
rect 20260 3383 20312 3392
rect 20260 3349 20269 3383
rect 20269 3349 20303 3383
rect 20303 3349 20312 3383
rect 20260 3340 20312 3349
rect 20628 3383 20680 3392
rect 20628 3349 20637 3383
rect 20637 3349 20671 3383
rect 20671 3349 20680 3383
rect 20628 3340 20680 3349
rect 21364 3340 21416 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 2504 3136 2556 3188
rect 3056 3179 3108 3188
rect 3056 3145 3065 3179
rect 3065 3145 3099 3179
rect 3099 3145 3108 3179
rect 3056 3136 3108 3145
rect 8944 3136 8996 3188
rect 9312 3179 9364 3188
rect 9312 3145 9321 3179
rect 9321 3145 9355 3179
rect 9355 3145 9364 3179
rect 9312 3136 9364 3145
rect 9496 3136 9548 3188
rect 11428 3136 11480 3188
rect 11520 3136 11572 3188
rect 19340 3179 19392 3188
rect 3700 3111 3752 3120
rect 3700 3077 3709 3111
rect 3709 3077 3743 3111
rect 3743 3077 3752 3111
rect 3700 3068 3752 3077
rect 5264 3068 5316 3120
rect 8668 3111 8720 3120
rect 8668 3077 8677 3111
rect 8677 3077 8711 3111
rect 8711 3077 8720 3111
rect 8668 3068 8720 3077
rect 9128 3068 9180 3120
rect 11888 3111 11940 3120
rect 5356 2975 5408 2984
rect 5356 2941 5365 2975
rect 5365 2941 5399 2975
rect 5399 2941 5408 2975
rect 5356 2932 5408 2941
rect 8300 2975 8352 2984
rect 8300 2941 8309 2975
rect 8309 2941 8343 2975
rect 8343 2941 8352 2975
rect 8300 2932 8352 2941
rect 9496 2975 9548 2984
rect 9496 2941 9505 2975
rect 9505 2941 9539 2975
rect 9539 2941 9548 2975
rect 9496 2932 9548 2941
rect 9772 2975 9824 2984
rect 9772 2941 9781 2975
rect 9781 2941 9815 2975
rect 9815 2941 9824 2975
rect 9772 2932 9824 2941
rect 1860 2796 1912 2848
rect 8208 2864 8260 2916
rect 8392 2907 8444 2916
rect 8392 2873 8401 2907
rect 8401 2873 8435 2907
rect 8435 2873 8444 2907
rect 8392 2864 8444 2873
rect 8668 2864 8720 2916
rect 11888 3077 11897 3111
rect 11897 3077 11931 3111
rect 11931 3077 11940 3111
rect 11888 3068 11940 3077
rect 10876 3043 10928 3052
rect 10876 3009 10885 3043
rect 10885 3009 10919 3043
rect 10919 3009 10928 3043
rect 10876 3000 10928 3009
rect 11060 3000 11112 3052
rect 12532 3043 12584 3052
rect 12532 3009 12541 3043
rect 12541 3009 12575 3043
rect 12575 3009 12584 3043
rect 12532 3000 12584 3009
rect 12808 3043 12860 3052
rect 12808 3009 12817 3043
rect 12817 3009 12851 3043
rect 12851 3009 12860 3043
rect 12808 3000 12860 3009
rect 13360 3000 13412 3052
rect 14096 2975 14148 2984
rect 14096 2941 14105 2975
rect 14105 2941 14139 2975
rect 14139 2941 14148 2975
rect 14096 2932 14148 2941
rect 10968 2907 11020 2916
rect 4896 2796 4948 2848
rect 5080 2839 5132 2848
rect 5080 2805 5089 2839
rect 5089 2805 5123 2839
rect 5123 2805 5132 2839
rect 5080 2796 5132 2805
rect 6552 2839 6604 2848
rect 6552 2805 6561 2839
rect 6561 2805 6595 2839
rect 6595 2805 6604 2839
rect 6552 2796 6604 2805
rect 10140 2796 10192 2848
rect 10968 2873 10977 2907
rect 10977 2873 11011 2907
rect 11011 2873 11020 2907
rect 10968 2864 11020 2873
rect 12624 2907 12676 2916
rect 12624 2873 12633 2907
rect 12633 2873 12667 2907
rect 12667 2873 12676 2907
rect 15844 3043 15896 3052
rect 15844 3009 15853 3043
rect 15853 3009 15887 3043
rect 15887 3009 15896 3043
rect 15844 3000 15896 3009
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 18328 3000 18380 3052
rect 12624 2864 12676 2873
rect 16304 2932 16356 2984
rect 19340 3145 19349 3179
rect 19349 3145 19383 3179
rect 19383 3145 19392 3179
rect 19340 3136 19392 3145
rect 19064 3068 19116 3120
rect 20904 3136 20956 3188
rect 23480 3136 23532 3188
rect 23388 3068 23440 3120
rect 20260 3000 20312 3052
rect 23756 3043 23808 3052
rect 23756 3009 23765 3043
rect 23765 3009 23799 3043
rect 23799 3009 23808 3043
rect 23756 3000 23808 3009
rect 23940 3000 23992 3052
rect 19432 2932 19484 2984
rect 17776 2864 17828 2916
rect 14740 2796 14792 2848
rect 15292 2839 15344 2848
rect 15292 2805 15301 2839
rect 15301 2805 15335 2839
rect 15335 2805 15344 2839
rect 15292 2796 15344 2805
rect 18052 2796 18104 2848
rect 19340 2864 19392 2916
rect 23296 2932 23348 2984
rect 25136 2932 25188 2984
rect 19984 2796 20036 2848
rect 20720 2796 20772 2848
rect 20996 2796 21048 2848
rect 23848 2907 23900 2916
rect 23848 2873 23857 2907
rect 23857 2873 23891 2907
rect 23891 2873 23900 2907
rect 23848 2864 23900 2873
rect 21364 2796 21416 2848
rect 23664 2796 23716 2848
rect 24860 2839 24912 2848
rect 24860 2805 24869 2839
rect 24869 2805 24903 2839
rect 24903 2805 24912 2839
rect 24860 2796 24912 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1676 2592 1728 2644
rect 4252 2592 4304 2644
rect 4528 2592 4580 2644
rect 7932 2592 7984 2644
rect 9496 2592 9548 2644
rect 9864 2592 9916 2644
rect 11152 2635 11204 2644
rect 4896 2524 4948 2576
rect 10232 2567 10284 2576
rect 10232 2533 10241 2567
rect 10241 2533 10275 2567
rect 10275 2533 10284 2567
rect 10232 2524 10284 2533
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 11980 2635 12032 2644
rect 11980 2601 11989 2635
rect 11989 2601 12023 2635
rect 12023 2601 12032 2635
rect 11980 2592 12032 2601
rect 12716 2592 12768 2644
rect 14096 2635 14148 2644
rect 14096 2601 14105 2635
rect 14105 2601 14139 2635
rect 14139 2601 14148 2635
rect 14096 2592 14148 2601
rect 15844 2592 15896 2644
rect 16948 2635 17000 2644
rect 16948 2601 16957 2635
rect 16957 2601 16991 2635
rect 16991 2601 17000 2635
rect 16948 2592 17000 2601
rect 20076 2592 20128 2644
rect 21732 2592 21784 2644
rect 11060 2524 11112 2576
rect 664 2456 716 2508
rect 2872 2456 2924 2508
rect 2872 2295 2924 2304
rect 2872 2261 2881 2295
rect 2881 2261 2915 2295
rect 2915 2261 2924 2295
rect 2872 2252 2924 2261
rect 6092 2456 6144 2508
rect 6000 2431 6052 2440
rect 6000 2397 6009 2431
rect 6009 2397 6043 2431
rect 6043 2397 6052 2431
rect 6000 2388 6052 2397
rect 8760 2499 8812 2508
rect 8760 2465 8769 2499
rect 8769 2465 8803 2499
rect 8803 2465 8812 2499
rect 8760 2456 8812 2465
rect 10048 2456 10100 2508
rect 10232 2388 10284 2440
rect 8852 2320 8904 2372
rect 10692 2320 10744 2372
rect 13636 2456 13688 2508
rect 12716 2431 12768 2440
rect 12716 2397 12725 2431
rect 12725 2397 12759 2431
rect 12759 2397 12768 2431
rect 12716 2388 12768 2397
rect 12808 2388 12860 2440
rect 13544 2388 13596 2440
rect 14740 2388 14792 2440
rect 16212 2567 16264 2576
rect 16212 2533 16221 2567
rect 16221 2533 16255 2567
rect 16255 2533 16264 2567
rect 16212 2524 16264 2533
rect 17592 2524 17644 2576
rect 18420 2524 18472 2576
rect 19524 2524 19576 2576
rect 20904 2524 20956 2576
rect 23296 2524 23348 2576
rect 23940 2524 23992 2576
rect 25228 2524 25280 2576
rect 15568 2431 15620 2440
rect 15568 2397 15577 2431
rect 15577 2397 15611 2431
rect 15611 2397 15620 2431
rect 15568 2388 15620 2397
rect 19432 2456 19484 2508
rect 22468 2456 22520 2508
rect 23756 2456 23808 2508
rect 24952 2456 25004 2508
rect 18420 2388 18472 2440
rect 21548 2431 21600 2440
rect 18880 2320 18932 2372
rect 21548 2397 21557 2431
rect 21557 2397 21591 2431
rect 21591 2397 21600 2431
rect 21548 2388 21600 2397
rect 22284 2388 22336 2440
rect 11244 2252 11296 2304
rect 11428 2252 11480 2304
rect 13728 2252 13780 2304
rect 14464 2295 14516 2304
rect 14464 2261 14473 2295
rect 14473 2261 14507 2295
rect 14507 2261 14516 2295
rect 14464 2252 14516 2261
rect 17592 2252 17644 2304
rect 18052 2295 18104 2304
rect 18052 2261 18061 2295
rect 18061 2261 18095 2295
rect 18095 2261 18104 2295
rect 18052 2252 18104 2261
rect 20904 2295 20956 2304
rect 20904 2261 20913 2295
rect 20913 2261 20947 2295
rect 20947 2261 20956 2295
rect 20904 2252 20956 2261
rect 22468 2252 22520 2304
rect 22652 2252 22704 2304
rect 23940 2252 23992 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 10048 2048 10100 2100
rect 18052 2048 18104 2100
rect 6276 1980 6328 2032
rect 11980 1980 12032 2032
rect 15476 144 15528 196
rect 6920 76 6972 128
rect 8300 76 8352 128
rect 9772 76 9824 128
rect 14464 76 14516 128
rect 21088 76 21140 128
rect 21916 76 21968 128
rect 22376 76 22428 128
rect 24308 76 24360 128
rect 26240 76 26292 128
rect 27528 76 27580 128
rect 15568 8 15620 60
rect 19340 8 19392 60
<< metal2 >>
rect 24950 26888 25006 26897
rect 24950 26823 25006 26832
rect 24766 25800 24822 25809
rect 24766 25735 24822 25744
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 24780 24410 24808 25735
rect 24768 24404 24820 24410
rect 24768 24346 24820 24352
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24964 23866 24992 26823
rect 27618 25392 27674 25401
rect 27618 25327 27674 25336
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 25148 23866 25176 24210
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 24122 23760 24178 23769
rect 24122 23695 24178 23704
rect 23664 23520 23716 23526
rect 23664 23462 23716 23468
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 15568 23180 15620 23186
rect 15568 23122 15620 23128
rect 18972 23180 19024 23186
rect 18972 23122 19024 23128
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15580 22438 15608 23122
rect 16394 22672 16450 22681
rect 16394 22607 16450 22616
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16250 15332 16934
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15304 15960 15332 16186
rect 15384 15972 15436 15978
rect 15304 15932 15384 15960
rect 15384 15914 15436 15920
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 15488 15638 15516 17070
rect 13820 15632 13872 15638
rect 13820 15574 13872 15580
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6380 13734 6408 14418
rect 12714 14376 12770 14385
rect 12624 14340 12676 14346
rect 12676 14320 12714 14328
rect 12676 14311 12770 14320
rect 12676 14300 12756 14311
rect 12624 14282 12676 14288
rect 13096 14006 13124 14418
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 8022 13696 8078 13705
rect 6182 13288 6238 13297
rect 6182 13223 6238 13232
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6090 12200 6146 12209
rect 6090 12135 6146 12144
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 3054 11792 3110 11801
rect 3054 11727 3110 11736
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1435 4072 1487 4078
rect 1412 4020 1435 4060
rect 1412 4014 1487 4020
rect 1412 3942 1440 4014
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 664 2508 716 2514
rect 664 2450 716 2456
rect 386 82 442 480
rect 676 82 704 2450
rect 386 54 704 82
rect 1122 82 1178 480
rect 1412 82 1440 3878
rect 1688 2650 1716 7346
rect 2962 7032 3018 7041
rect 2962 6967 3018 6976
rect 2976 4214 3004 6967
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 2502 3768 2558 3777
rect 2502 3703 2558 3712
rect 2516 3194 2544 3703
rect 3068 3602 3096 11727
rect 4158 11248 4214 11257
rect 4158 11183 4214 11192
rect 5998 11248 6054 11257
rect 5998 11183 6054 11192
rect 4172 4282 4200 11183
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5078 10704 5134 10713
rect 5078 10639 5134 10648
rect 4526 8528 4582 8537
rect 4526 8463 4582 8472
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3068 3194 3096 3538
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 1122 54 1440 82
rect 1872 82 1900 2790
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2884 2310 2912 2450
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 1950 82 2006 480
rect 1872 54 2006 82
rect 386 0 442 54
rect 1122 0 1178 54
rect 1950 0 2006 54
rect 2778 82 2834 480
rect 2884 82 2912 2246
rect 2778 54 2912 82
rect 3252 82 3280 3878
rect 3698 3224 3754 3233
rect 3698 3159 3754 3168
rect 3712 3126 3740 3159
rect 3700 3120 3752 3126
rect 3700 3062 3752 3068
rect 3514 82 3570 480
rect 4172 241 4200 3878
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4264 2417 4292 2586
rect 4250 2408 4306 2417
rect 4250 2343 4306 2352
rect 4158 232 4214 241
rect 4158 167 4214 176
rect 3252 54 3570 82
rect 2778 0 2834 54
rect 3514 0 3570 54
rect 4342 82 4398 480
rect 4448 82 4476 3878
rect 4540 2650 4568 8463
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 4908 2582 4936 2790
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 5000 377 5028 4966
rect 5092 4826 5120 10639
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6012 5370 6040 11183
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 5368 4729 5396 4966
rect 6104 4826 6132 12135
rect 6196 5710 6224 13223
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 5354 4720 5410 4729
rect 5172 4684 5224 4690
rect 5354 4655 5410 4664
rect 6184 4684 6236 4690
rect 5172 4626 5224 4632
rect 6184 4626 6236 4632
rect 5184 3942 5212 4626
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6196 3942 6224 4626
rect 6288 4146 6316 4966
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6276 4004 6328 4010
rect 6276 3946 6328 3952
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 5092 2854 5120 3538
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 5092 513 5120 2790
rect 5184 785 5212 3878
rect 5262 3768 5318 3777
rect 5262 3703 5318 3712
rect 5276 3670 5304 3703
rect 5264 3664 5316 3670
rect 5316 3624 5396 3652
rect 5264 3606 5316 3612
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 5170 776 5226 785
rect 5170 711 5226 720
rect 5078 504 5134 513
rect 5078 439 5134 448
rect 4986 368 5042 377
rect 4986 303 5042 312
rect 4342 54 4476 82
rect 5170 82 5226 480
rect 5276 82 5304 3062
rect 5368 2990 5396 3624
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5356 2984 5408 2990
rect 5460 2961 5488 3470
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5356 2926 5408 2932
rect 5446 2952 5502 2961
rect 5446 2887 5502 2896
rect 6012 2689 6040 3878
rect 5998 2680 6054 2689
rect 5998 2615 6054 2624
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6012 1601 6040 2382
rect 6104 2281 6132 2450
rect 6090 2272 6146 2281
rect 6090 2207 6146 2216
rect 5998 1592 6054 1601
rect 5998 1527 6054 1536
rect 5170 54 5304 82
rect 5906 82 5962 480
rect 6196 82 6224 3878
rect 6288 2038 6316 3946
rect 6276 2032 6328 2038
rect 6276 1974 6328 1980
rect 5906 54 6224 82
rect 6380 82 6408 13670
rect 8022 13631 8078 13640
rect 6642 13016 6698 13025
rect 6642 12951 6698 12960
rect 6656 6866 6684 12951
rect 7010 12744 7066 12753
rect 7010 12679 7066 12688
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6734 10024 6790 10033
rect 6734 9959 6790 9968
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6656 6458 6684 6802
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6656 5370 6684 5714
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6564 3369 6592 4014
rect 6748 3738 6776 9959
rect 6826 8528 6882 8537
rect 6826 8463 6882 8472
rect 6840 7002 6868 8463
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6550 3360 6606 3369
rect 6550 3295 6606 3304
rect 6552 2848 6604 2854
rect 6656 2836 6684 3538
rect 6604 2808 6684 2836
rect 6552 2790 6604 2796
rect 6564 1329 6592 2790
rect 6550 1320 6606 1329
rect 6550 1255 6606 1264
rect 6734 82 6790 480
rect 6932 134 6960 11494
rect 7024 5370 7052 12679
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 7944 11558 7972 12242
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7576 10266 7604 10406
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7654 9208 7710 9217
rect 7654 9143 7710 9152
rect 7286 8664 7342 8673
rect 7286 8599 7342 8608
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7116 6254 7144 6598
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7116 5273 7144 6190
rect 7300 5778 7328 8599
rect 7668 7954 7696 9143
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7668 7546 7696 7890
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7576 6458 7604 6802
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7300 5370 7328 5714
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7102 5264 7158 5273
rect 7102 5199 7158 5208
rect 7392 5137 7420 6054
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7484 5370 7512 5578
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7668 5166 7696 5510
rect 7656 5160 7708 5166
rect 7378 5128 7434 5137
rect 7656 5102 7708 5108
rect 7378 5063 7434 5072
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 6380 54 6790 82
rect 6920 128 6972 134
rect 7116 105 7144 4082
rect 7300 3942 7328 4626
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7300 1057 7328 3878
rect 7668 3505 7696 4422
rect 7654 3496 7710 3505
rect 7654 3431 7710 3440
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7484 3233 7512 3334
rect 7470 3224 7526 3233
rect 7470 3159 7526 3168
rect 7286 1048 7342 1057
rect 7286 983 7342 992
rect 6920 70 6972 76
rect 7102 96 7158 105
rect 4342 0 4398 54
rect 5170 0 5226 54
rect 5906 0 5962 54
rect 6734 0 6790 54
rect 7102 31 7158 40
rect 7562 82 7618 480
rect 7760 82 7788 10406
rect 7838 9480 7894 9489
rect 7838 9415 7894 9424
rect 7852 8090 7880 9415
rect 8036 8956 8064 13631
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 8298 12880 8354 12889
rect 8298 12815 8354 12824
rect 8312 12442 8340 12815
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 12360 12306 12388 13806
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12636 12986 12664 13330
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12544 12374 12572 12854
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11900 11898 11928 12174
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 11888 11212 11940 11218
rect 11992 11200 12020 11766
rect 12360 11626 12388 12242
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11940 11172 12020 11200
rect 11888 11154 11940 11160
rect 11900 10810 11928 11154
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 12084 10198 12112 11290
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12072 10192 12124 10198
rect 12072 10134 12124 10140
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 10876 9920 10928 9926
rect 10782 9888 10838 9897
rect 10876 9862 10928 9868
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 10782 9823 10838 9832
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8114 9072 8170 9081
rect 8114 9007 8170 9016
rect 7944 8928 8064 8956
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7852 3233 7880 4966
rect 7838 3224 7894 3233
rect 7838 3159 7894 3168
rect 7944 2650 7972 8928
rect 8128 6866 8156 9007
rect 8390 7848 8446 7857
rect 8390 7783 8446 7792
rect 8298 7712 8354 7721
rect 8298 7647 8354 7656
rect 8312 7546 8340 7647
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8312 7342 8340 7482
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8312 6118 8340 6802
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8312 5574 8340 6054
rect 8404 5710 8432 7783
rect 8772 7002 8800 9522
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9310 8936 9366 8945
rect 9310 8871 9366 8880
rect 9680 8900 9732 8906
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8864 7206 8892 7890
rect 8956 7546 8984 8774
rect 9324 8634 9352 8871
rect 9680 8842 9732 8848
rect 9692 8634 9720 8842
rect 9954 8800 10010 8809
rect 9954 8735 10010 8744
rect 9968 8634 9996 8735
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9324 8430 9352 8570
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8944 7268 8996 7274
rect 8944 7210 8996 7216
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8864 6662 8892 7142
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8588 6322 8616 6598
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8300 5568 8352 5574
rect 8220 5528 8300 5556
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 8036 3670 8064 5102
rect 8128 4214 8156 5170
rect 8220 5030 8248 5528
rect 8300 5510 8352 5516
rect 8404 5370 8432 5646
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 8116 4072 8168 4078
rect 8220 4049 8248 4966
rect 8496 4826 8524 5714
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8312 4214 8340 4626
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8496 4146 8524 4626
rect 8588 4554 8616 6258
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8680 5137 8708 5510
rect 8852 5160 8904 5166
rect 8666 5128 8722 5137
rect 8852 5102 8904 5108
rect 8666 5063 8722 5072
rect 8864 4826 8892 5102
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8760 4616 8812 4622
rect 8956 4593 8984 7210
rect 9048 6186 9076 8298
rect 10060 7478 10088 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10704 9178 10732 9386
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 8129 10732 8298
rect 10690 8120 10746 8129
rect 10690 8055 10746 8064
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 10428 7818 10456 7890
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10152 7410 10180 7686
rect 10428 7546 10456 7754
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10612 7546 10640 7686
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9140 6866 9168 7142
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9140 6769 9168 6802
rect 9126 6760 9182 6769
rect 9126 6695 9182 6704
rect 9310 6760 9366 6769
rect 9310 6695 9366 6704
rect 9324 6390 9352 6695
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9416 6322 9444 7278
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9508 6633 9536 6666
rect 9494 6624 9550 6633
rect 9494 6559 9550 6568
rect 9508 6458 9536 6559
rect 10152 6458 10180 6802
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10506 6352 10562 6361
rect 9404 6316 9456 6322
rect 10506 6287 10562 6296
rect 10692 6316 10744 6322
rect 9404 6258 9456 6264
rect 9036 6180 9088 6186
rect 9036 6122 9088 6128
rect 9048 5914 9076 6122
rect 9416 5914 9444 6258
rect 10520 6254 10548 6287
rect 10692 6258 10744 6264
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9036 5908 9088 5914
rect 9404 5908 9456 5914
rect 9088 5868 9352 5896
rect 9036 5850 9088 5856
rect 9034 5808 9090 5817
rect 9034 5743 9090 5752
rect 9048 5710 9076 5743
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9220 5636 9272 5642
rect 9220 5578 9272 5584
rect 8760 4558 8812 4564
rect 8942 4584 8998 4593
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8116 4014 8168 4020
rect 8206 4040 8262 4049
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 8024 3392 8076 3398
rect 8128 3380 8156 4014
rect 8206 3975 8262 3984
rect 8772 3641 8800 4558
rect 8942 4519 8998 4528
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 8758 3632 8814 3641
rect 8668 3596 8720 3602
rect 8758 3567 8814 3576
rect 8668 3538 8720 3544
rect 8076 3352 8156 3380
rect 8024 3334 8076 3340
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8036 1737 8064 3334
rect 8680 3126 8708 3538
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 8668 3120 8720 3126
rect 8956 3097 8984 3130
rect 9140 3126 9168 4014
rect 9232 4010 9260 5578
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9324 3194 9352 5868
rect 9404 5850 9456 5856
rect 9692 5166 9720 6054
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10704 5914 10732 6258
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10796 5778 10824 9823
rect 10888 9518 10916 9862
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 11520 9444 11572 9450
rect 11520 9386 11572 9392
rect 11532 9110 11560 9386
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11716 8838 11744 9862
rect 11808 9722 11836 10066
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11900 9382 11928 9998
rect 11980 9444 12032 9450
rect 11980 9386 12032 9392
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11992 9042 12020 9386
rect 12084 9382 12112 10134
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11348 7750 11376 8366
rect 11520 8356 11572 8362
rect 11520 8298 11572 8304
rect 11532 7954 11560 8298
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10980 7274 11008 7482
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 11348 6934 11376 7346
rect 11532 7002 11560 7890
rect 11716 7546 11744 8774
rect 11808 8498 11836 8774
rect 11992 8634 12020 8978
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10980 6118 11008 6394
rect 10968 6112 11020 6118
rect 10888 6072 10968 6100
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10060 5302 10088 5714
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10048 5296 10100 5302
rect 10048 5238 10100 5244
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9416 4078 9444 5034
rect 9692 4826 9720 5102
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9876 4758 9904 4966
rect 9968 4826 9996 5170
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9864 4752 9916 4758
rect 9678 4720 9734 4729
rect 9864 4694 9916 4700
rect 9954 4720 10010 4729
rect 9678 4655 9734 4664
rect 10704 4690 10732 5306
rect 10784 5296 10836 5302
rect 10784 5238 10836 5244
rect 9954 4655 10010 4664
rect 10692 4684 10744 4690
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9128 3120 9180 3126
rect 8668 3062 8720 3068
rect 8942 3088 8998 3097
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 8022 1728 8078 1737
rect 8022 1663 8078 1672
rect 8220 921 8248 2858
rect 8312 2553 8340 2926
rect 8680 2922 8708 3062
rect 9128 3062 9180 3068
rect 8942 3023 8998 3032
rect 9508 2990 9536 3130
rect 9600 3097 9628 3878
rect 9692 3738 9720 4655
rect 9968 4010 9996 4655
rect 10692 4626 10744 4632
rect 10704 4214 10732 4626
rect 10692 4208 10744 4214
rect 10138 4176 10194 4185
rect 10692 4150 10744 4156
rect 10138 4111 10194 4120
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9586 3088 9642 3097
rect 9586 3023 9642 3032
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 8298 2544 8354 2553
rect 8298 2479 8354 2488
rect 8404 1193 8432 2858
rect 9508 2650 9536 2926
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 8772 1737 8800 2450
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 8758 1728 8814 1737
rect 8758 1663 8814 1672
rect 8390 1184 8446 1193
rect 8390 1119 8446 1128
rect 8206 912 8262 921
rect 8206 847 8262 856
rect 7562 54 7788 82
rect 8298 128 8354 480
rect 8298 76 8300 128
rect 8352 76 8354 128
rect 7562 0 7618 54
rect 8298 0 8354 76
rect 8864 82 8892 2314
rect 9126 82 9182 480
rect 9784 134 9812 2926
rect 9876 2650 9904 3878
rect 10152 3777 10180 4111
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10138 3768 10194 3777
rect 10289 3760 10585 3780
rect 10138 3703 10194 3712
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10152 2854 10180 3538
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 10060 2106 10088 2450
rect 10048 2100 10100 2106
rect 10048 2042 10100 2048
rect 8864 54 9182 82
rect 9772 128 9824 134
rect 9772 70 9824 76
rect 9954 82 10010 480
rect 10152 82 10180 2790
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10232 2576 10284 2582
rect 10232 2518 10284 2524
rect 10244 2446 10272 2518
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10704 2378 10732 3470
rect 10692 2372 10744 2378
rect 10692 2314 10744 2320
rect 9126 0 9182 54
rect 9954 54 10180 82
rect 10690 82 10746 480
rect 10796 82 10824 5238
rect 10888 3738 10916 6072
rect 10968 6054 11020 6060
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10980 3534 11008 5034
rect 11072 4758 11100 6734
rect 11900 6458 11928 6938
rect 11992 6458 12020 8570
rect 12084 8090 12112 9318
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12176 8430 12204 8910
rect 12268 8634 12296 10406
rect 12544 10130 12572 10746
rect 12636 10742 12664 12174
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12728 10198 12756 12718
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12820 10470 12848 11222
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12820 9994 12848 10066
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12728 9722 12756 9862
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12912 9518 12940 10542
rect 12992 10532 13044 10538
rect 12992 10474 13044 10480
rect 13004 10266 13032 10474
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12990 9752 13046 9761
rect 12990 9687 13046 9696
rect 13004 9654 13032 9687
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12268 8362 12296 8570
rect 12256 8356 12308 8362
rect 12256 8298 12308 8304
rect 12268 8090 12296 8298
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12268 7342 12296 8026
rect 12360 7750 12388 8978
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12544 8498 12572 8910
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 8090 12572 8434
rect 12728 8294 12756 9454
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12268 7002 12296 7278
rect 12820 7274 12848 7754
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 12820 7002 12848 7210
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11992 6254 12020 6394
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11532 5846 11560 6054
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 11164 5302 11192 5782
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 11256 5234 11284 5646
rect 11532 5370 11560 5782
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 11624 4622 11652 5510
rect 12176 5370 12204 6802
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12544 6118 12572 6734
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12544 5914 12572 6054
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 12728 5846 12756 6190
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11336 4072 11388 4078
rect 11520 4072 11572 4078
rect 11388 4032 11468 4060
rect 11336 4014 11388 4020
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10888 3058 10916 3402
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10980 2922 11008 3334
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 11072 2582 11100 2994
rect 11164 2650 11192 3470
rect 11440 3194 11468 4032
rect 11520 4014 11572 4020
rect 11532 3194 11560 4014
rect 11624 3738 11652 4558
rect 11808 4214 11836 4694
rect 12452 4622 12480 5578
rect 12728 4826 12756 5646
rect 12820 5370 12848 5782
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12452 4282 12480 4422
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 12544 4146 12572 4558
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 12636 3670 12664 4694
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12728 4078 12756 4422
rect 13096 4154 13124 13942
rect 13268 13796 13320 13802
rect 13268 13738 13320 13744
rect 13280 12782 13308 13738
rect 13372 13734 13400 14418
rect 13464 14006 13492 14894
rect 13740 14618 13768 15438
rect 13832 15162 13860 15574
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15488 15162 15516 15574
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 14292 14550 14320 14758
rect 14280 14544 14332 14550
rect 14280 14486 14332 14492
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14108 14074 14136 14418
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 14292 13870 14320 14486
rect 14384 14278 14412 14894
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13280 12306 13308 12582
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13280 11558 13308 12242
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 13188 10266 13216 10950
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13280 10198 13308 11494
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13280 9450 13308 10134
rect 13372 9761 13400 13670
rect 13740 13190 13768 13806
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13740 12850 13768 13126
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13544 12776 13596 12782
rect 13832 12730 13860 13670
rect 14384 13462 14412 14214
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14372 13456 14424 13462
rect 14372 13398 14424 13404
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 13544 12718 13596 12724
rect 13556 12442 13584 12718
rect 13740 12702 13860 12730
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13464 11082 13492 11630
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13358 9752 13414 9761
rect 13464 9722 13492 10066
rect 13358 9687 13414 9696
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 13464 9058 13492 9658
rect 13556 9625 13584 11562
rect 13648 10538 13676 11698
rect 13740 11558 13768 12702
rect 13924 12646 13952 13330
rect 14476 12782 14504 13330
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14568 12889 14596 13194
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14554 12880 14610 12889
rect 14554 12815 14610 12824
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14476 12646 14504 12718
rect 14740 12708 14792 12714
rect 14740 12650 14792 12656
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13832 11898 13860 12242
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13740 11286 13768 11494
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13636 10532 13688 10538
rect 13636 10474 13688 10480
rect 13832 10130 13860 11834
rect 14108 11694 14136 12174
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14292 9722 14320 9862
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 13542 9616 13598 9625
rect 13542 9551 13598 9560
rect 14278 9616 14334 9625
rect 14334 9586 14412 9602
rect 14334 9580 14424 9586
rect 14334 9574 14372 9580
rect 14278 9551 14334 9560
rect 14372 9522 14424 9528
rect 13912 9444 13964 9450
rect 13912 9386 13964 9392
rect 13924 9110 13952 9386
rect 13372 9030 13492 9058
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 13188 8090 13216 8842
rect 13372 8838 13400 9030
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13188 6322 13216 6938
rect 13372 6866 13400 8774
rect 13464 8634 13492 8910
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13740 8566 13768 9046
rect 13924 8809 13952 9046
rect 14004 8900 14056 8906
rect 14004 8842 14056 8848
rect 13910 8800 13966 8809
rect 13910 8735 13966 8744
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13464 8022 13492 8230
rect 13452 8016 13504 8022
rect 13452 7958 13504 7964
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13372 6458 13400 6802
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13556 6236 13584 8502
rect 14016 7886 14044 8842
rect 14476 8634 14504 12582
rect 14556 12096 14608 12102
rect 14752 12084 14780 12650
rect 14844 12102 14872 12786
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 14608 12056 14780 12084
rect 14832 12096 14884 12102
rect 14556 12038 14608 12044
rect 14832 12038 14884 12044
rect 14568 11830 14596 12038
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14844 11762 14872 12038
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14568 11354 14596 11630
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14844 10674 14872 11698
rect 15108 11620 15160 11626
rect 15108 11562 15160 11568
rect 15120 11354 15148 11562
rect 15304 11558 15332 12378
rect 15396 12238 15424 13262
rect 15580 12850 15608 22374
rect 16408 17882 16436 22607
rect 18984 22438 19012 23122
rect 20904 23112 20956 23118
rect 20994 23080 21050 23089
rect 20956 23060 20994 23066
rect 20904 23054 20994 23060
rect 20916 23038 20994 23054
rect 20994 23015 21050 23024
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 18328 22432 18380 22438
rect 18328 22374 18380 22380
rect 18972 22432 19024 22438
rect 18972 22374 19024 22380
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 16132 17338 16160 17682
rect 17788 17338 17816 17682
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 16120 17332 16172 17338
rect 16120 17274 16172 17280
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15672 15502 15700 16526
rect 16132 16114 16160 17274
rect 17040 17128 17092 17134
rect 17040 17070 17092 17076
rect 16396 17060 16448 17066
rect 16396 17002 16448 17008
rect 16212 16720 16264 16726
rect 16212 16662 16264 16668
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16132 15638 16160 16050
rect 16224 15910 16252 16662
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16120 15632 16172 15638
rect 16120 15574 16172 15580
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15672 14618 15700 15438
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 15948 14074 15976 14350
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15936 13864 15988 13870
rect 15856 13824 15936 13852
rect 15856 13190 15884 13824
rect 15936 13806 15988 13812
rect 16132 13734 16160 14350
rect 16224 14006 16252 15846
rect 16408 15162 16436 17002
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16684 15910 16712 16458
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16408 14822 16436 15098
rect 16500 14890 16528 15302
rect 16684 15065 16712 15846
rect 16670 15056 16726 15065
rect 16670 14991 16726 15000
rect 16488 14884 16540 14890
rect 16488 14826 16540 14832
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16500 14385 16528 14826
rect 17052 14822 17080 17070
rect 17788 15638 17816 17274
rect 18156 16726 18184 17478
rect 18144 16720 18196 16726
rect 18196 16680 18276 16708
rect 18144 16662 18196 16668
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18156 16114 18184 16526
rect 18248 16250 18276 16680
rect 18340 16590 18368 22374
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 23308 22001 23336 22918
rect 23676 22681 23704 23462
rect 23662 22672 23718 22681
rect 23662 22607 23718 22616
rect 23294 21992 23350 22001
rect 23294 21927 23350 21936
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 23572 18828 23624 18834
rect 23572 18770 23624 18776
rect 23584 18086 23612 18770
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 23572 18080 23624 18086
rect 23572 18022 23624 18028
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 21548 17740 21600 17746
rect 21548 17682 21600 17688
rect 21560 17338 21588 17682
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21548 17332 21600 17338
rect 21548 17274 21600 17280
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18144 16108 18196 16114
rect 18144 16050 18196 16056
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 17776 15632 17828 15638
rect 17776 15574 17828 15580
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17420 15026 17448 15438
rect 17788 15162 17816 15574
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 17052 14618 17080 14758
rect 17420 14618 17448 14962
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 16856 14544 16908 14550
rect 16856 14486 16908 14492
rect 16486 14376 16542 14385
rect 16486 14311 16542 14320
rect 16868 14006 16896 14486
rect 16212 14000 16264 14006
rect 16212 13942 16264 13948
rect 16856 14000 16908 14006
rect 16856 13942 16908 13948
rect 16120 13728 16172 13734
rect 16120 13670 16172 13676
rect 16132 13530 16160 13670
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16868 13462 16896 13942
rect 17788 13530 17816 15098
rect 18156 14890 18184 15642
rect 18340 15638 18368 16526
rect 18984 15638 19012 17070
rect 19064 16992 19116 16998
rect 19064 16934 19116 16940
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 19076 16250 19104 16934
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 19076 15910 19104 16186
rect 19260 16114 19288 16390
rect 19536 16114 19564 16594
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 18972 15632 19024 15638
rect 18972 15574 19024 15580
rect 18984 15162 19012 15574
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18144 14884 18196 14890
rect 18144 14826 18196 14832
rect 18984 14618 19012 15098
rect 19260 15026 19288 16050
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19444 15706 19472 15846
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 19444 14822 19472 15438
rect 19536 15434 19564 16050
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19524 15428 19576 15434
rect 19524 15370 19576 15376
rect 20732 15162 20760 16934
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20732 14822 20760 15098
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 18972 14612 19024 14618
rect 18972 14554 19024 14560
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17880 14074 17908 14350
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 18788 14000 18840 14006
rect 18788 13942 18840 13948
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15580 12238 15608 12786
rect 15856 12714 15884 13126
rect 16776 12850 16804 13262
rect 18340 13190 18368 13670
rect 18800 13326 18828 13942
rect 18892 13938 18920 14214
rect 19444 14006 19472 14758
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19168 13433 19196 13874
rect 19812 13802 19840 14010
rect 20180 13841 20208 14758
rect 20824 14482 20852 17070
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 21546 16552 21602 16561
rect 21546 16487 21602 16496
rect 21560 16250 21588 16487
rect 21548 16244 21600 16250
rect 21548 16186 21600 16192
rect 21560 16046 21588 16186
rect 21548 16040 21600 16046
rect 21548 15982 21600 15988
rect 21652 15706 21680 16594
rect 21836 16250 21864 17614
rect 21916 17332 21968 17338
rect 21916 17274 21968 17280
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21836 15910 21864 16186
rect 21824 15904 21876 15910
rect 21824 15846 21876 15852
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20536 14000 20588 14006
rect 20536 13942 20588 13948
rect 20166 13832 20222 13841
rect 19800 13796 19852 13802
rect 20166 13767 20222 13776
rect 19800 13738 19852 13744
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19248 13456 19300 13462
rect 19154 13424 19210 13433
rect 19248 13398 19300 13404
rect 19154 13359 19210 13368
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18340 12986 18368 13126
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 15844 12708 15896 12714
rect 15844 12650 15896 12656
rect 16040 12646 16068 12718
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15396 11898 15424 12174
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15764 11626 15792 12038
rect 15752 11620 15804 11626
rect 15752 11562 15804 11568
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15304 11218 15332 11494
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15764 11082 15792 11562
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14568 8514 14596 9862
rect 14646 9752 14702 9761
rect 14646 9687 14702 9696
rect 14660 9586 14688 9687
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14752 9110 14780 10202
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14844 9518 14872 9998
rect 15304 9926 15332 10542
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 14844 9382 14872 9454
rect 15292 9444 15344 9450
rect 15292 9386 15344 9392
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14740 9104 14792 9110
rect 14740 9046 14792 9052
rect 14844 8956 14872 9318
rect 15304 8974 15332 9386
rect 14752 8928 14872 8956
rect 15292 8968 15344 8974
rect 14646 8664 14702 8673
rect 14646 8599 14702 8608
rect 14476 8486 14596 8514
rect 14370 8120 14426 8129
rect 14370 8055 14426 8064
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 13740 7478 13768 7822
rect 14016 7721 14044 7822
rect 14002 7712 14058 7721
rect 14002 7647 14058 7656
rect 13728 7472 13780 7478
rect 13728 7414 13780 7420
rect 13556 6208 13676 6236
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13188 5166 13216 6054
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13188 4622 13216 5102
rect 13648 5080 13676 6208
rect 13740 5914 13768 7414
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13832 6390 13860 6870
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 14200 5234 14228 7346
rect 14384 7342 14412 8055
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14292 6798 14320 7142
rect 14384 7002 14412 7278
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14292 6458 14320 6734
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 13556 5052 13676 5080
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 13464 4282 13492 4626
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13096 4126 13216 4154
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11440 2310 11468 3130
rect 11900 3126 11928 3538
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 12544 3058 12572 3402
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12806 3360 12862 3369
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 11978 2952 12034 2961
rect 12636 2922 12664 3334
rect 12806 3295 12862 3304
rect 12820 3058 12848 3295
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 11978 2887 12034 2896
rect 12624 2916 12676 2922
rect 11992 2650 12020 2887
rect 12624 2858 12676 2864
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12728 2446 12756 2586
rect 12820 2446 12848 2994
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 11428 2304 11480 2310
rect 11428 2246 11480 2252
rect 10690 54 10824 82
rect 11256 82 11284 2246
rect 11980 2032 12032 2038
rect 11980 1974 12032 1980
rect 11518 82 11574 480
rect 11256 54 11574 82
rect 11992 82 12020 1974
rect 12346 82 12402 480
rect 11992 54 12402 82
rect 9954 0 10010 54
rect 10690 0 10746 54
rect 11518 0 11574 54
rect 12346 0 12402 54
rect 13082 82 13138 480
rect 13188 82 13216 4126
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13372 3058 13400 3946
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13556 2446 13584 5052
rect 14200 5030 14228 5170
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 13634 4584 13690 4593
rect 13634 4519 13690 4528
rect 13648 2514 13676 4519
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13082 54 13216 82
rect 13740 82 13768 2246
rect 13924 1601 13952 3878
rect 14016 3738 14044 4626
rect 14200 3738 14228 4966
rect 14292 4010 14320 5510
rect 14384 4758 14412 6938
rect 14476 6610 14504 8486
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14568 7410 14596 7686
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14554 6624 14610 6633
rect 14476 6582 14554 6610
rect 14554 6559 14610 6568
rect 14568 6458 14596 6559
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14660 6225 14688 8599
rect 14646 6216 14702 6225
rect 14646 6151 14702 6160
rect 14648 5568 14700 5574
rect 14752 5556 14780 8928
rect 15292 8910 15344 8916
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15304 8294 15332 8910
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 14832 7880 14884 7886
rect 14830 7848 14832 7857
rect 14884 7848 14886 7857
rect 14830 7783 14886 7792
rect 14844 7546 14872 7783
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14844 7410 14872 7482
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 15120 7002 15148 7414
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15304 6866 15332 8230
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 14844 6118 14872 6802
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15290 6352 15346 6361
rect 15290 6287 15346 6296
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14700 5528 14780 5556
rect 14648 5510 14700 5516
rect 14660 5302 14688 5510
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14648 5092 14700 5098
rect 14648 5034 14700 5040
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14372 4752 14424 4758
rect 14372 4694 14424 4700
rect 14568 4690 14596 4966
rect 14660 4826 14688 5034
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14108 2650 14136 2926
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 14292 2417 14320 3946
rect 14660 3942 14688 4558
rect 14752 4486 14780 5170
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14646 3496 14702 3505
rect 14646 3431 14702 3440
rect 14660 3398 14688 3431
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 14752 2446 14780 2790
rect 14740 2440 14792 2446
rect 14278 2408 14334 2417
rect 14740 2382 14792 2388
rect 14278 2343 14334 2352
rect 14464 2304 14516 2310
rect 14752 2281 14780 2382
rect 14464 2246 14516 2252
rect 14738 2272 14794 2281
rect 13910 1592 13966 1601
rect 13910 1527 13966 1536
rect 13910 82 13966 480
rect 14476 134 14504 2246
rect 14738 2207 14794 2216
rect 13740 54 13966 82
rect 14464 128 14516 134
rect 14464 70 14516 76
rect 14738 82 14794 480
rect 14844 82 14872 6054
rect 15120 5914 15148 6190
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15304 5778 15332 6287
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15304 4826 15332 5714
rect 15396 5370 15424 9454
rect 15488 8838 15516 10406
rect 15580 10062 15608 10950
rect 15936 10532 15988 10538
rect 15936 10474 15988 10480
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15488 8498 15516 8774
rect 15764 8566 15792 9590
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15488 7750 15516 8434
rect 15568 8356 15620 8362
rect 15568 8298 15620 8304
rect 15580 7954 15608 8298
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15488 7546 15516 7686
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15672 7478 15700 7686
rect 15764 7478 15792 8502
rect 15856 8498 15884 9454
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15856 8294 15884 8434
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15660 7472 15712 7478
rect 15660 7414 15712 7420
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 15764 7002 15792 7414
rect 15856 7410 15884 8230
rect 15948 7750 15976 10474
rect 16040 10198 16068 12582
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16224 10470 16252 11086
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 16224 9654 16252 10406
rect 16316 9994 16344 10950
rect 16592 10656 16620 11086
rect 16684 10810 16712 12718
rect 16776 12442 16804 12786
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 18432 12374 18460 13126
rect 19260 12986 19288 13398
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18602 12744 18658 12753
rect 18602 12679 18658 12688
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 16856 11824 16908 11830
rect 16856 11766 16908 11772
rect 16868 11286 16896 11766
rect 17236 11558 17264 12242
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 17880 11626 17908 12174
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17868 11620 17920 11626
rect 17868 11562 17920 11568
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16672 10668 16724 10674
rect 16592 10628 16672 10656
rect 16672 10610 16724 10616
rect 16488 10192 16540 10198
rect 16488 10134 16540 10140
rect 16304 9988 16356 9994
rect 16304 9930 16356 9936
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16224 7750 16252 7890
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 16224 7206 16252 7686
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15856 6798 15884 7142
rect 15844 6792 15896 6798
rect 16316 6769 16344 9386
rect 16408 7274 16436 9862
rect 16500 9042 16528 10134
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16592 9722 16620 10066
rect 16684 10062 16712 10610
rect 17052 10198 17080 11290
rect 17236 11014 17264 11494
rect 17880 11014 17908 11562
rect 17972 11082 18000 12038
rect 18064 11558 18092 12174
rect 18234 11792 18290 11801
rect 18234 11727 18290 11736
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18064 11150 18092 11494
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17236 10470 17264 10950
rect 17498 10704 17554 10713
rect 17498 10639 17554 10648
rect 17684 10668 17736 10674
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17236 10266 17264 10406
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17040 10192 17092 10198
rect 17040 10134 17092 10140
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 17052 9722 17080 10134
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16592 7886 16620 9658
rect 17420 9654 17448 9862
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 16960 8634 16988 8978
rect 17328 8634 17356 8978
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16592 7342 16620 7686
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 15844 6734 15896 6740
rect 16302 6760 16358 6769
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15488 6322 15516 6598
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15856 6118 15884 6734
rect 16302 6695 16358 6704
rect 16316 6458 16344 6695
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15658 5808 15714 5817
rect 15658 5743 15714 5752
rect 15672 5710 15700 5743
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15396 4690 15424 5306
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 14936 3670 14964 3946
rect 15304 3738 15332 4626
rect 15396 4049 15424 4626
rect 15382 4040 15438 4049
rect 15382 3975 15438 3984
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 14924 3664 14976 3670
rect 14924 3606 14976 3612
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15304 1737 15332 2790
rect 15290 1728 15346 1737
rect 15290 1663 15346 1672
rect 15488 202 15516 5510
rect 15672 5370 15700 5646
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15580 4604 15608 5170
rect 15672 5166 15700 5306
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15856 5098 15884 6054
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 15660 4616 15712 4622
rect 15580 4576 15660 4604
rect 15660 4558 15712 4564
rect 15672 4282 15700 4558
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15580 2446 15608 3334
rect 15856 3058 15884 3878
rect 15948 3516 15976 6122
rect 16132 5370 16160 6394
rect 16316 5914 16344 6394
rect 16408 6322 16436 7210
rect 16670 6896 16726 6905
rect 16670 6831 16726 6840
rect 16764 6860 16816 6866
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16040 5030 16068 5170
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 16040 4729 16068 4966
rect 16026 4720 16082 4729
rect 16026 4655 16082 4664
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16028 4548 16080 4554
rect 16028 4490 16080 4496
rect 16040 4078 16068 4490
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 16132 4010 16160 4626
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16224 4078 16252 4422
rect 16684 4154 16712 6831
rect 16764 6802 16816 6808
rect 16776 6458 16804 6802
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 16684 4126 16804 4154
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 16040 3670 16068 3878
rect 16028 3664 16080 3670
rect 16028 3606 16080 3612
rect 16028 3528 16080 3534
rect 15948 3488 16028 3516
rect 16028 3470 16080 3476
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15856 2650 15884 2994
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15476 196 15528 202
rect 15476 138 15528 144
rect 13082 0 13138 54
rect 13910 0 13966 54
rect 14738 54 14872 82
rect 15566 60 15622 480
rect 14738 0 14794 54
rect 15566 8 15568 60
rect 15620 8 15622 60
rect 16132 82 16160 3946
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 16224 2582 16252 3334
rect 16316 2990 16344 3878
rect 16776 3602 16804 4126
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 16302 82 16358 480
rect 16132 54 16358 82
rect 16868 82 16896 7822
rect 17328 7410 17356 8570
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 17328 7002 17356 7346
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17132 6180 17184 6186
rect 17132 6122 17184 6128
rect 17040 5636 17092 5642
rect 17040 5578 17092 5584
rect 17052 4554 17080 5578
rect 17144 4690 17172 6122
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17328 5370 17356 5646
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 17040 4548 17092 4554
rect 17040 4490 17092 4496
rect 17052 4282 17080 4490
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 17144 3738 17172 4626
rect 17512 4486 17540 10639
rect 17684 10610 17736 10616
rect 17696 10470 17724 10610
rect 17880 10606 17908 10950
rect 17972 10742 18000 11018
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 18064 10674 18092 11086
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17696 10062 17724 10406
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17696 9518 17724 9998
rect 17880 9994 17908 10542
rect 18052 10532 18104 10538
rect 18052 10474 18104 10480
rect 18064 10266 18092 10474
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17684 9512 17736 9518
rect 17684 9454 17736 9460
rect 17880 9110 17908 9930
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18064 9178 18092 9454
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17604 7954 17632 8910
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17604 7002 17632 7890
rect 17880 7342 17908 7958
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17776 7200 17828 7206
rect 17696 7160 17776 7188
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 17696 5166 17724 7160
rect 17776 7142 17828 7148
rect 17880 7018 17908 7278
rect 17788 6990 17908 7018
rect 17788 6186 17816 6990
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17132 3732 17184 3738
rect 17132 3674 17184 3680
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 16960 2650 16988 3470
rect 17604 3398 17632 3470
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 17604 2310 17632 2518
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17604 1329 17632 2246
rect 17590 1320 17646 1329
rect 17590 1255 17646 1264
rect 17130 82 17186 480
rect 16868 54 17186 82
rect 17696 82 17724 5102
rect 17788 4282 17816 6122
rect 17880 5574 17908 6802
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17880 5137 17908 5510
rect 17866 5128 17922 5137
rect 17866 5063 17922 5072
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17788 4010 17816 4218
rect 18064 4146 18092 4558
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 17776 4004 17828 4010
rect 17776 3946 17828 3952
rect 17788 3738 17816 3946
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 17788 2922 17816 3674
rect 18156 3058 18184 4966
rect 18248 4554 18276 11727
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18340 10742 18368 10950
rect 18328 10736 18380 10742
rect 18328 10678 18380 10684
rect 18340 9926 18368 10678
rect 18510 10024 18566 10033
rect 18510 9959 18566 9968
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18328 9716 18380 9722
rect 18328 9658 18380 9664
rect 18340 5778 18368 9658
rect 18432 9042 18460 9862
rect 18524 9636 18552 9959
rect 18616 9761 18644 12679
rect 18708 12442 18736 12786
rect 20272 12782 20300 13126
rect 20548 12850 20576 13942
rect 20732 13258 20760 14350
rect 20824 14074 20852 14418
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20720 13252 20772 13258
rect 20720 13194 20772 13200
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18972 12164 19024 12170
rect 18972 12106 19024 12112
rect 18984 11762 19012 12106
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18708 10130 18736 10542
rect 18800 10470 18828 11494
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18602 9752 18658 9761
rect 18602 9687 18658 9696
rect 18524 9608 18644 9636
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18432 5846 18460 6598
rect 18420 5840 18472 5846
rect 18420 5782 18472 5788
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18340 5370 18368 5714
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18432 4826 18460 5782
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18236 4548 18288 4554
rect 18236 4490 18288 4496
rect 18328 3460 18380 3466
rect 18328 3402 18380 3408
rect 18340 3058 18368 3402
rect 18420 3392 18472 3398
rect 18420 3334 18472 3340
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 18064 2310 18092 2790
rect 18432 2582 18460 3334
rect 18420 2576 18472 2582
rect 18420 2518 18472 2524
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 18064 2106 18092 2246
rect 18052 2100 18104 2106
rect 18052 2042 18104 2048
rect 17958 82 18014 480
rect 18432 377 18460 2382
rect 18418 368 18474 377
rect 18418 303 18474 312
rect 17696 54 18014 82
rect 18524 82 18552 5646
rect 18616 4154 18644 9608
rect 18800 8090 18828 10406
rect 18984 9042 19012 11698
rect 19076 11626 19104 12038
rect 19536 11694 19564 12582
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 20272 12442 20300 12718
rect 20824 12646 20852 13330
rect 20916 13190 20944 14350
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20824 12374 20852 12582
rect 20812 12368 20864 12374
rect 20812 12310 20864 12316
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20534 12200 20590 12209
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 19524 11688 19576 11694
rect 19524 11630 19576 11636
rect 19064 11620 19116 11626
rect 19064 11562 19116 11568
rect 19076 11286 19104 11562
rect 19168 11558 19196 11630
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19064 11280 19116 11286
rect 19064 11222 19116 11228
rect 19168 11218 19196 11494
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19996 11354 20024 12174
rect 20272 11762 20300 12174
rect 20824 12170 20852 12310
rect 20534 12135 20590 12144
rect 20812 12164 20864 12170
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19064 10532 19116 10538
rect 19064 10474 19116 10480
rect 18972 9036 19024 9042
rect 18972 8978 19024 8984
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18892 8498 18920 8774
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18708 7546 18736 8026
rect 18984 8022 19012 8978
rect 18972 8016 19024 8022
rect 18972 7958 19024 7964
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18880 7268 18932 7274
rect 18880 7210 18932 7216
rect 18696 6724 18748 6730
rect 18696 6666 18748 6672
rect 18708 5624 18736 6666
rect 18788 5636 18840 5642
rect 18708 5596 18788 5624
rect 18708 4826 18736 5596
rect 18788 5578 18840 5584
rect 18696 4820 18748 4826
rect 18696 4762 18748 4768
rect 18616 4126 18828 4154
rect 18800 3670 18828 4126
rect 18788 3664 18840 3670
rect 18788 3606 18840 3612
rect 18892 2378 18920 7210
rect 19076 6866 19104 10474
rect 19168 10470 19196 11154
rect 19352 10674 19380 11154
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19156 10464 19208 10470
rect 19156 10406 19208 10412
rect 19168 9586 19196 10406
rect 19352 10266 19380 10610
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19340 10260 19392 10266
rect 19340 10202 19392 10208
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19352 9518 19380 10066
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19904 9518 19932 9998
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19892 9512 19944 9518
rect 19944 9472 20024 9500
rect 19892 9454 19944 9460
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19156 7948 19208 7954
rect 19156 7890 19208 7896
rect 19168 7546 19196 7890
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 19076 6254 19104 6802
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 19168 5710 19196 7482
rect 19260 6866 19288 9318
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19996 9110 20024 9472
rect 19984 9104 20036 9110
rect 19984 9046 20036 9052
rect 19430 8936 19486 8945
rect 19430 8871 19486 8880
rect 19444 8566 19472 8871
rect 19996 8634 20024 9046
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 19444 7410 19472 8502
rect 20548 8362 20576 12135
rect 20812 12106 20864 12112
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20640 10470 20668 11494
rect 20824 11218 20852 12106
rect 21008 11898 21036 14758
rect 21652 13814 21680 15642
rect 21928 15638 21956 17274
rect 22008 17128 22060 17134
rect 22008 17070 22060 17076
rect 21916 15632 21968 15638
rect 21916 15574 21968 15580
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21836 14890 21864 15438
rect 21928 15162 21956 15574
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 21824 14884 21876 14890
rect 21824 14826 21876 14832
rect 21928 14618 21956 15098
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 21916 14272 21968 14278
rect 21916 14214 21968 14220
rect 21928 14006 21956 14214
rect 21916 14000 21968 14006
rect 21916 13942 21968 13948
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 21652 13786 21772 13814
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21284 12646 21312 13670
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21652 12850 21680 13262
rect 21640 12844 21692 12850
rect 21640 12786 21692 12792
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21284 12374 21312 12582
rect 21272 12368 21324 12374
rect 21272 12310 21324 12316
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 21088 11688 21140 11694
rect 21088 11630 21140 11636
rect 21100 11354 21128 11630
rect 21284 11626 21312 12310
rect 21272 11620 21324 11626
rect 21272 11562 21324 11568
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 20812 11212 20864 11218
rect 20812 11154 20864 11160
rect 20824 10810 20852 11154
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 21100 10674 21128 11086
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 21192 10062 21220 11290
rect 21284 10470 21312 11562
rect 21456 11212 21508 11218
rect 21456 11154 21508 11160
rect 21468 10810 21496 11154
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21284 10266 21312 10406
rect 21744 10266 21772 13786
rect 21836 12374 21864 13874
rect 21928 13870 21956 13942
rect 22020 13938 22048 17070
rect 22112 16114 22140 18022
rect 22836 17740 22888 17746
rect 22836 17682 22888 17688
rect 22744 17060 22796 17066
rect 22744 17002 22796 17008
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 22204 15994 22232 16934
rect 22560 16652 22612 16658
rect 22560 16594 22612 16600
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 22112 15966 22232 15994
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 21916 13864 21968 13870
rect 21916 13806 21968 13812
rect 22020 12986 22048 13874
rect 22008 12980 22060 12986
rect 22008 12922 22060 12928
rect 22112 12832 22140 15966
rect 22284 15904 22336 15910
rect 22020 12804 22140 12832
rect 22204 15864 22284 15892
rect 21824 12368 21876 12374
rect 21824 12310 21876 12316
rect 22020 11898 22048 12804
rect 22100 12708 22152 12714
rect 22100 12650 22152 12656
rect 22112 12442 22140 12650
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 22020 11286 22048 11834
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 22020 10742 22048 11222
rect 22008 10736 22060 10742
rect 22008 10678 22060 10684
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21732 10260 21784 10266
rect 21732 10202 21784 10208
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21192 9722 21220 9998
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 21100 9178 21128 9454
rect 21180 9376 21232 9382
rect 21284 9364 21312 10202
rect 21232 9336 21312 9364
rect 21180 9318 21232 9324
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21192 9110 21220 9318
rect 21744 9110 21772 10202
rect 22204 9178 22232 15864
rect 22284 15846 22336 15852
rect 22480 15638 22508 16050
rect 22468 15632 22520 15638
rect 22468 15574 22520 15580
rect 22282 11248 22338 11257
rect 22282 11183 22338 11192
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 21180 9104 21232 9110
rect 21180 9046 21232 9052
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 20812 8492 20864 8498
rect 20812 8434 20864 8440
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 20628 8356 20680 8362
rect 20628 8298 20680 8304
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 20548 8090 20576 8298
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19536 7206 19564 7890
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19156 5704 19208 5710
rect 19156 5646 19208 5652
rect 19156 5568 19208 5574
rect 19260 5556 19288 6802
rect 19904 6322 19932 6802
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19996 6322 20024 6598
rect 19892 6316 19944 6322
rect 19892 6258 19944 6264
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 19524 6248 19576 6254
rect 19524 6190 19576 6196
rect 19904 6202 19932 6258
rect 19536 5778 19564 6190
rect 19904 6174 20116 6202
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 20088 5778 20116 6174
rect 20640 5846 20668 8298
rect 20824 7410 20852 8434
rect 21192 8294 21220 9046
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21192 8022 21220 8230
rect 21284 8090 21312 8910
rect 21824 8288 21876 8294
rect 21824 8230 21876 8236
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 21180 8016 21232 8022
rect 21180 7958 21232 7964
rect 21192 7546 21220 7958
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 21192 7002 21220 7482
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 20916 6254 20944 6734
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 20916 5914 20944 6190
rect 21192 6186 21220 6938
rect 21836 6662 21864 8230
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 21928 6866 21956 7822
rect 22204 7546 22232 9114
rect 22296 8362 22324 11183
rect 22466 11112 22522 11121
rect 22466 11047 22522 11056
rect 22374 9480 22430 9489
rect 22374 9415 22430 9424
rect 22284 8356 22336 8362
rect 22284 8298 22336 8304
rect 22192 7540 22244 7546
rect 22192 7482 22244 7488
rect 22388 7410 22416 9415
rect 22284 7404 22336 7410
rect 22284 7346 22336 7352
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 21916 6860 21968 6866
rect 21916 6802 21968 6808
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21824 6656 21876 6662
rect 21824 6598 21876 6604
rect 21180 6180 21232 6186
rect 21180 6122 21232 6128
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 21284 5778 21312 6598
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 20076 5772 20128 5778
rect 20076 5714 20128 5720
rect 21272 5772 21324 5778
rect 21272 5714 21324 5720
rect 19208 5528 19288 5556
rect 19984 5568 20036 5574
rect 19156 5510 19208 5516
rect 19984 5510 20036 5516
rect 19168 5166 19196 5510
rect 19996 5234 20024 5510
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 20088 5166 20116 5714
rect 20260 5636 20312 5642
rect 20260 5578 20312 5584
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 20076 5160 20128 5166
rect 20076 5102 20128 5108
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 20168 5024 20220 5030
rect 20168 4966 20220 4972
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 18984 4282 19012 4694
rect 18972 4276 19024 4282
rect 18972 4218 19024 4224
rect 18984 4185 19012 4218
rect 18970 4176 19026 4185
rect 18970 4111 19026 4120
rect 19076 3126 19104 4966
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 20180 4622 20208 4966
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 19168 3942 19196 4558
rect 20076 4480 20128 4486
rect 20272 4457 20300 5578
rect 21284 5370 21312 5714
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 21468 5098 21496 5306
rect 21732 5228 21784 5234
rect 21732 5170 21784 5176
rect 21456 5092 21508 5098
rect 21456 5034 21508 5040
rect 21468 4758 21496 5034
rect 21744 4826 21772 5170
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 21456 4752 21508 4758
rect 21456 4694 21508 4700
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 20076 4422 20128 4428
rect 20258 4448 20314 4457
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19340 3664 19392 3670
rect 19340 3606 19392 3612
rect 19352 3194 19380 3606
rect 19536 3534 19564 3878
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19340 2916 19392 2922
rect 19340 2858 19392 2864
rect 18880 2372 18932 2378
rect 18880 2314 18932 2320
rect 18694 82 18750 480
rect 18524 54 18750 82
rect 19352 66 19380 2858
rect 19444 2514 19472 2926
rect 19536 2582 19564 3470
rect 20088 3466 20116 4422
rect 20258 4383 20314 4392
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20180 3738 20208 3878
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20076 3460 20128 3466
rect 20076 3402 20128 3408
rect 20640 3398 20668 4626
rect 21468 4010 21496 4694
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21456 4004 21508 4010
rect 21456 3946 21508 3952
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20732 3670 20760 3878
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20902 3632 20958 3641
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20272 3058 20300 3334
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19524 2576 19576 2582
rect 19524 2518 19576 2524
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19522 82 19578 480
rect 19996 82 20024 2790
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 15566 0 15622 8
rect 16302 0 16358 54
rect 17130 0 17186 54
rect 17958 0 18014 54
rect 18694 0 18750 54
rect 19340 60 19392 66
rect 19340 2 19392 8
rect 19522 54 20024 82
rect 20088 82 20116 2586
rect 20272 241 20300 2994
rect 20640 2417 20668 3334
rect 20732 2854 20760 3606
rect 20902 3567 20958 3576
rect 20916 3534 20944 3567
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20916 3194 20944 3470
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 20994 2952 21050 2961
rect 20994 2887 21050 2896
rect 21178 2952 21234 2961
rect 21178 2887 21234 2896
rect 21008 2854 21036 2887
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 20626 2408 20682 2417
rect 20626 2343 20682 2352
rect 20916 2310 20944 2518
rect 20904 2304 20956 2310
rect 20904 2246 20956 2252
rect 20916 921 20944 2246
rect 21192 1057 21220 2887
rect 21376 2854 21404 3334
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21376 1737 21404 2790
rect 21560 2446 21588 4422
rect 22112 4154 22140 7210
rect 22296 6662 22324 7346
rect 22284 6656 22336 6662
rect 22284 6598 22336 6604
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 22204 4282 22232 4558
rect 22192 4276 22244 4282
rect 22192 4218 22244 4224
rect 22112 4126 22232 4154
rect 22204 4078 22232 4126
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 21732 3936 21784 3942
rect 21732 3878 21784 3884
rect 21744 2650 21772 3878
rect 21732 2644 21784 2650
rect 21732 2586 21784 2592
rect 21744 2553 21772 2586
rect 21730 2544 21786 2553
rect 21730 2479 21786 2488
rect 22296 2446 22324 6598
rect 22480 4622 22508 11047
rect 22572 9518 22600 16594
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22664 9654 22692 16526
rect 22756 13462 22784 17002
rect 22848 16998 22876 17682
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 23204 17128 23256 17134
rect 23204 17070 23256 17076
rect 22836 16992 22888 16998
rect 22836 16934 22888 16940
rect 22928 15972 22980 15978
rect 22928 15914 22980 15920
rect 22836 14544 22888 14550
rect 22836 14486 22888 14492
rect 22848 14006 22876 14486
rect 22836 14000 22888 14006
rect 22836 13942 22888 13948
rect 22744 13456 22796 13462
rect 22744 13398 22796 13404
rect 22756 12986 22784 13398
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 22848 12646 22876 13262
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22848 11937 22876 12582
rect 22834 11928 22890 11937
rect 22834 11863 22890 11872
rect 22652 9648 22704 9654
rect 22652 9590 22704 9596
rect 22560 9512 22612 9518
rect 22560 9454 22612 9460
rect 22940 9382 22968 15914
rect 23110 15464 23166 15473
rect 23110 15399 23166 15408
rect 23124 15162 23152 15399
rect 23112 15156 23164 15162
rect 23112 15098 23164 15104
rect 23124 14958 23152 15098
rect 23112 14952 23164 14958
rect 23112 14894 23164 14900
rect 23216 14328 23244 17070
rect 23308 14396 23336 17478
rect 23480 17060 23532 17066
rect 23480 17002 23532 17008
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23400 15910 23428 16594
rect 23388 15904 23440 15910
rect 23388 15846 23440 15852
rect 23388 14884 23440 14890
rect 23388 14826 23440 14832
rect 23400 14550 23428 14826
rect 23388 14544 23440 14550
rect 23388 14486 23440 14492
rect 23308 14368 23428 14396
rect 23216 14300 23336 14328
rect 23204 13932 23256 13938
rect 23204 13874 23256 13880
rect 23216 13462 23244 13874
rect 23204 13456 23256 13462
rect 23204 13398 23256 13404
rect 23020 13184 23072 13190
rect 23020 13126 23072 13132
rect 23032 12442 23060 13126
rect 23020 12436 23072 12442
rect 23020 12378 23072 12384
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 23204 12300 23256 12306
rect 23204 12242 23256 12248
rect 23032 11558 23060 12242
rect 23216 12102 23244 12242
rect 23204 12096 23256 12102
rect 23204 12038 23256 12044
rect 23216 11830 23244 12038
rect 23204 11824 23256 11830
rect 23204 11766 23256 11772
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 23032 10810 23060 11086
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 23308 10606 23336 14300
rect 23400 11898 23428 14368
rect 23388 11892 23440 11898
rect 23388 11834 23440 11840
rect 23400 11558 23428 11834
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 23492 10742 23520 17002
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 23572 14408 23624 14414
rect 23572 14350 23624 14356
rect 23584 13190 23612 14350
rect 23572 13184 23624 13190
rect 23572 13126 23624 13132
rect 23584 11830 23612 13126
rect 23572 11824 23624 11830
rect 23572 11766 23624 11772
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23584 10742 23612 11086
rect 23480 10736 23532 10742
rect 23480 10678 23532 10684
rect 23572 10736 23624 10742
rect 23572 10678 23624 10684
rect 23296 10600 23348 10606
rect 23296 10542 23348 10548
rect 23308 10266 23336 10542
rect 23492 10538 23520 10678
rect 23480 10532 23532 10538
rect 23480 10474 23532 10480
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23308 9722 23336 10202
rect 23388 10056 23440 10062
rect 23388 9998 23440 10004
rect 23296 9716 23348 9722
rect 23296 9658 23348 9664
rect 23400 9586 23428 9998
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23296 9512 23348 9518
rect 23296 9454 23348 9460
rect 22928 9376 22980 9382
rect 22928 9318 22980 9324
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 22940 9178 22968 9318
rect 22928 9172 22980 9178
rect 22928 9114 22980 9120
rect 23124 8974 23152 9318
rect 23204 9104 23256 9110
rect 23204 9046 23256 9052
rect 23112 8968 23164 8974
rect 23112 8910 23164 8916
rect 22560 8832 22612 8838
rect 22560 8774 22612 8780
rect 22572 8498 22600 8774
rect 23020 8560 23072 8566
rect 23020 8502 23072 8508
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22744 7268 22796 7274
rect 22744 7210 22796 7216
rect 22756 5642 22784 7210
rect 23032 6798 23060 8502
rect 23124 8090 23152 8910
rect 23216 8634 23244 9046
rect 23308 8634 23336 9454
rect 23400 8974 23428 9522
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 23296 8628 23348 8634
rect 23296 8570 23348 8576
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 23676 7954 23704 15098
rect 23768 15026 23796 18702
rect 24136 18358 24164 23695
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24584 22432 24636 22438
rect 24688 22420 24716 23122
rect 25148 23089 25176 23802
rect 27632 23322 27660 25327
rect 27620 23316 27672 23322
rect 27620 23258 27672 23264
rect 25134 23080 25190 23089
rect 25134 23015 25190 23024
rect 24858 22672 24914 22681
rect 24858 22607 24914 22616
rect 24636 22392 24716 22420
rect 24584 22374 24636 22380
rect 24596 22001 24624 22374
rect 24582 21992 24638 22001
rect 24582 21927 24638 21936
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24766 21720 24822 21729
rect 24872 21690 24900 22607
rect 24766 21655 24822 21664
rect 24860 21684 24912 21690
rect 24780 21146 24808 21655
rect 24860 21626 24912 21632
rect 25320 21344 25372 21350
rect 25320 21286 25372 21292
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20534 24716 20946
rect 24766 20632 24822 20641
rect 24766 20567 24822 20576
rect 24676 20528 24728 20534
rect 24676 20470 24728 20476
rect 24780 20058 24808 20567
rect 24952 20256 25004 20262
rect 24952 20198 25004 20204
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24676 19916 24728 19922
rect 24676 19858 24728 19864
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24688 19446 24716 19858
rect 24766 19544 24822 19553
rect 24766 19479 24822 19488
rect 24676 19440 24728 19446
rect 24676 19382 24728 19388
rect 24780 18970 24808 19479
rect 24860 19168 24912 19174
rect 24860 19110 24912 19116
rect 24768 18964 24820 18970
rect 24768 18906 24820 18912
rect 24676 18828 24728 18834
rect 24676 18770 24728 18776
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 18426 24716 18770
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24124 18352 24176 18358
rect 24124 18294 24176 18300
rect 23940 18216 23992 18222
rect 23940 18158 23992 18164
rect 24216 18216 24268 18222
rect 24216 18158 24268 18164
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23768 14618 23796 14962
rect 23860 14890 23888 17614
rect 23848 14884 23900 14890
rect 23848 14826 23900 14832
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23768 13802 23796 14214
rect 23952 13814 23980 18158
rect 24228 16794 24256 18158
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24872 17354 24900 19110
rect 24688 17326 24900 17354
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 24124 16584 24176 16590
rect 24124 16526 24176 16532
rect 24032 14408 24084 14414
rect 24032 14350 24084 14356
rect 24044 13938 24072 14350
rect 24032 13932 24084 13938
rect 24032 13874 24084 13880
rect 24136 13814 24164 16526
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24216 15564 24268 15570
rect 24216 15506 24268 15512
rect 24228 15162 24256 15506
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24216 15156 24268 15162
rect 24216 15098 24268 15104
rect 24308 15088 24360 15094
rect 24214 15056 24270 15065
rect 24270 15036 24308 15042
rect 24270 15030 24360 15036
rect 24270 15014 24348 15030
rect 24214 14991 24270 15000
rect 24584 14884 24636 14890
rect 24584 14826 24636 14832
rect 24596 14414 24624 14826
rect 24584 14408 24636 14414
rect 24584 14350 24636 14356
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 23756 13796 23808 13802
rect 23952 13786 24072 13814
rect 24136 13786 24256 13814
rect 23756 13738 23808 13744
rect 23768 12918 23796 13738
rect 23940 13184 23992 13190
rect 23940 13126 23992 13132
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23952 12850 23980 13126
rect 23940 12844 23992 12850
rect 23940 12786 23992 12792
rect 23952 11762 23980 12786
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 23756 11620 23808 11626
rect 23756 11562 23808 11568
rect 23768 11014 23796 11562
rect 23952 11150 23980 11698
rect 23940 11144 23992 11150
rect 23940 11086 23992 11092
rect 23756 11008 23808 11014
rect 23756 10950 23808 10956
rect 23768 9897 23796 10950
rect 24044 10674 24072 13786
rect 24228 13462 24256 13786
rect 24308 13728 24360 13734
rect 24308 13670 24360 13676
rect 24216 13456 24268 13462
rect 24320 13433 24348 13670
rect 24216 13398 24268 13404
rect 24306 13424 24362 13433
rect 24306 13359 24362 13368
rect 24124 13320 24176 13326
rect 24124 13262 24176 13268
rect 24214 13288 24270 13297
rect 24136 12442 24164 13262
rect 24688 13258 24716 17326
rect 24964 17218 24992 20198
rect 25228 18624 25280 18630
rect 25228 18566 25280 18572
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 25056 17338 25084 17682
rect 25044 17332 25096 17338
rect 25096 17292 25176 17320
rect 25044 17274 25096 17280
rect 24872 17190 24992 17218
rect 24768 15496 24820 15502
rect 24768 15438 24820 15444
rect 24214 13223 24270 13232
rect 24676 13252 24728 13258
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 24228 12152 24256 13223
rect 24676 13194 24728 13200
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24688 12850 24716 13194
rect 24676 12844 24728 12850
rect 24676 12786 24728 12792
rect 24676 12300 24728 12306
rect 24676 12242 24728 12248
rect 24688 12170 24716 12242
rect 24136 12124 24256 12152
rect 24676 12164 24728 12170
rect 24032 10668 24084 10674
rect 24032 10610 24084 10616
rect 24044 10198 24072 10610
rect 24032 10192 24084 10198
rect 24032 10134 24084 10140
rect 23754 9888 23810 9897
rect 23754 9823 23810 9832
rect 23848 9648 23900 9654
rect 23848 9590 23900 9596
rect 23860 9450 23888 9590
rect 23756 9444 23808 9450
rect 23756 9386 23808 9392
rect 23848 9444 23900 9450
rect 23848 9386 23900 9392
rect 23768 8838 23796 9386
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 23848 8628 23900 8634
rect 23848 8570 23900 8576
rect 23860 8362 23888 8570
rect 24044 8537 24072 8774
rect 24030 8528 24086 8537
rect 24030 8463 24086 8472
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23848 8356 23900 8362
rect 23848 8298 23900 8304
rect 23768 8090 23796 8298
rect 23940 8288 23992 8294
rect 23940 8230 23992 8236
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 23676 7342 23704 7890
rect 23952 7886 23980 8230
rect 24032 8016 24084 8022
rect 24032 7958 24084 7964
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23664 7336 23716 7342
rect 23664 7278 23716 7284
rect 23952 7002 23980 7822
rect 24044 7546 24072 7958
rect 24032 7540 24084 7546
rect 24032 7482 24084 7488
rect 24136 7426 24164 12124
rect 24676 12106 24728 12112
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11898 24716 12106
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10742 24716 10950
rect 24676 10736 24728 10742
rect 24676 10678 24728 10684
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24780 9058 24808 15438
rect 24872 14890 24900 17190
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 24952 15972 25004 15978
rect 24952 15914 25004 15920
rect 24860 14884 24912 14890
rect 24860 14826 24912 14832
rect 24860 13456 24912 13462
rect 24860 13398 24912 13404
rect 24872 12986 24900 13398
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24964 10198 24992 15914
rect 25056 15910 25084 16594
rect 25044 15904 25096 15910
rect 25044 15846 25096 15852
rect 25056 12714 25084 15846
rect 25148 14550 25176 17292
rect 25240 17134 25268 18566
rect 25228 17128 25280 17134
rect 25228 17070 25280 17076
rect 25332 16250 25360 21286
rect 25410 18592 25466 18601
rect 25410 18527 25466 18536
rect 25424 17338 25452 18527
rect 25504 18080 25556 18086
rect 25504 18022 25556 18028
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25320 16244 25372 16250
rect 25320 16186 25372 16192
rect 25136 14544 25188 14550
rect 25136 14486 25188 14492
rect 25148 14074 25176 14486
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 25044 12708 25096 12714
rect 25044 12650 25096 12656
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 25056 11898 25084 12038
rect 25044 11892 25096 11898
rect 25044 11834 25096 11840
rect 25318 11384 25374 11393
rect 25318 11319 25374 11328
rect 25332 11286 25360 11319
rect 25320 11280 25372 11286
rect 25320 11222 25372 11228
rect 25332 10810 25360 11222
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25228 10464 25280 10470
rect 25228 10406 25280 10412
rect 24952 10192 25004 10198
rect 24952 10134 25004 10140
rect 24964 9722 24992 10134
rect 25240 10062 25268 10406
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 25516 9994 25544 18022
rect 25778 17504 25834 17513
rect 25778 17439 25834 17448
rect 25792 15162 25820 17439
rect 25780 15156 25832 15162
rect 25780 15098 25832 15104
rect 25792 14958 25820 15098
rect 25780 14952 25832 14958
rect 25780 14894 25832 14900
rect 25778 14376 25834 14385
rect 25778 14311 25834 14320
rect 25792 14074 25820 14311
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25792 13870 25820 14010
rect 25780 13864 25832 13870
rect 25780 13806 25832 13812
rect 25778 13696 25834 13705
rect 25778 13631 25834 13640
rect 25792 11898 25820 13631
rect 26238 12880 26294 12889
rect 26238 12815 26294 12824
rect 27618 12880 27674 12889
rect 27618 12815 27674 12824
rect 25780 11892 25832 11898
rect 25780 11834 25832 11840
rect 25792 11694 25820 11834
rect 25780 11688 25832 11694
rect 25780 11630 25832 11636
rect 25778 10296 25834 10305
rect 25778 10231 25834 10240
rect 25504 9988 25556 9994
rect 25504 9930 25556 9936
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 25318 9616 25374 9625
rect 25318 9551 25374 9560
rect 24688 9030 24808 9058
rect 24860 9104 24912 9110
rect 24860 9046 24912 9052
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24214 8392 24270 8401
rect 24214 8327 24270 8336
rect 24400 8356 24452 8362
rect 24044 7398 24164 7426
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 23112 6928 23164 6934
rect 23112 6870 23164 6876
rect 23020 6792 23072 6798
rect 23020 6734 23072 6740
rect 23032 5914 23060 6734
rect 23124 6390 23152 6870
rect 23572 6724 23624 6730
rect 23572 6666 23624 6672
rect 23112 6384 23164 6390
rect 23112 6326 23164 6332
rect 23020 5908 23072 5914
rect 23020 5850 23072 5856
rect 23584 5710 23612 6666
rect 23664 6180 23716 6186
rect 23664 6122 23716 6128
rect 23676 5846 23704 6122
rect 23664 5840 23716 5846
rect 23664 5782 23716 5788
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23572 5704 23624 5710
rect 23572 5646 23624 5652
rect 22744 5636 22796 5642
rect 22744 5578 22796 5584
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22468 4616 22520 4622
rect 22468 4558 22520 4564
rect 22376 4548 22428 4554
rect 22376 4490 22428 4496
rect 21548 2440 21600 2446
rect 21548 2382 21600 2388
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 21362 1728 21418 1737
rect 21362 1663 21418 1672
rect 21178 1048 21234 1057
rect 21178 983 21234 992
rect 20902 912 20958 921
rect 20902 847 20958 856
rect 20258 232 20314 241
rect 20258 167 20314 176
rect 20350 82 20406 480
rect 20088 54 20406 82
rect 19522 0 19578 54
rect 20350 0 20406 54
rect 21086 128 21142 480
rect 21086 76 21088 128
rect 21140 76 21142 128
rect 21086 0 21142 76
rect 21914 128 21970 480
rect 22388 134 22416 4490
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22480 3777 22508 4422
rect 22664 4282 22692 4966
rect 23400 4826 23428 5646
rect 23584 5273 23612 5646
rect 23676 5370 23704 5782
rect 23664 5364 23716 5370
rect 23664 5306 23716 5312
rect 23570 5264 23626 5273
rect 23570 5199 23626 5208
rect 23756 5092 23808 5098
rect 23756 5034 23808 5040
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 22652 4276 22704 4282
rect 22652 4218 22704 4224
rect 23032 4214 23060 4558
rect 23020 4208 23072 4214
rect 23020 4150 23072 4156
rect 23400 4146 23428 4762
rect 23480 4276 23532 4282
rect 23480 4218 23532 4224
rect 23388 4140 23440 4146
rect 23388 4082 23440 4088
rect 22466 3768 22522 3777
rect 22466 3703 22522 3712
rect 23492 3602 23520 4218
rect 23584 3738 23612 4966
rect 23768 4826 23796 5034
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 23768 4486 23796 4762
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 24044 4154 24072 7398
rect 24228 6798 24256 8327
rect 24400 8298 24452 8304
rect 24412 7886 24440 8298
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24400 7404 24452 7410
rect 24400 7346 24452 7352
rect 24412 7002 24440 7346
rect 24400 6996 24452 7002
rect 24400 6938 24452 6944
rect 24688 6934 24716 9030
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24780 8362 24808 8910
rect 24872 8634 24900 9046
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 25136 8492 25188 8498
rect 25136 8434 25188 8440
rect 24768 8356 24820 8362
rect 24768 8298 24820 8304
rect 25148 8022 25176 8434
rect 25136 8016 25188 8022
rect 25136 7958 25188 7964
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 24676 6928 24728 6934
rect 24676 6870 24728 6876
rect 24216 6792 24268 6798
rect 24216 6734 24268 6740
rect 24228 6390 24256 6734
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 6458 24716 6870
rect 24872 6798 24900 7346
rect 24860 6792 24912 6798
rect 24860 6734 24912 6740
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24216 6384 24268 6390
rect 24216 6326 24268 6332
rect 25228 6248 25280 6254
rect 25228 6190 25280 6196
rect 25044 5840 25096 5846
rect 25044 5782 25096 5788
rect 24952 5704 25004 5710
rect 24952 5646 25004 5652
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24964 5098 24992 5646
rect 25056 5370 25084 5782
rect 25044 5364 25096 5370
rect 25044 5306 25096 5312
rect 24952 5092 25004 5098
rect 24952 5034 25004 5040
rect 24964 4826 24992 5034
rect 24952 4820 25004 4826
rect 24952 4762 25004 4768
rect 24124 4752 24176 4758
rect 24124 4694 24176 4700
rect 24136 4282 24164 4694
rect 25056 4554 25084 5306
rect 25136 5160 25188 5166
rect 25240 5137 25268 6190
rect 25136 5102 25188 5108
rect 25226 5128 25282 5137
rect 25148 4865 25176 5102
rect 25226 5063 25282 5072
rect 25134 4856 25190 4865
rect 25134 4791 25190 4800
rect 25044 4548 25096 4554
rect 25044 4490 25096 4496
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24124 4276 24176 4282
rect 24124 4218 24176 4224
rect 24044 4146 24164 4154
rect 24044 4140 24176 4146
rect 24044 4126 24124 4140
rect 24124 4082 24176 4088
rect 25056 4078 25084 4490
rect 25332 4154 25360 9551
rect 25516 9110 25544 9930
rect 25792 9722 25820 10231
rect 26056 10056 26108 10062
rect 26056 9998 26108 10004
rect 26068 9722 26096 9998
rect 25780 9716 25832 9722
rect 25780 9658 25832 9664
rect 26056 9716 26108 9722
rect 26056 9658 26108 9664
rect 25792 9518 25820 9658
rect 25780 9512 25832 9518
rect 25780 9454 25832 9460
rect 25778 9208 25834 9217
rect 25778 9143 25834 9152
rect 25504 9104 25556 9110
rect 25504 9046 25556 9052
rect 25792 8634 25820 9143
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 25792 8430 25820 8570
rect 25780 8424 25832 8430
rect 25780 8366 25832 8372
rect 25686 8256 25742 8265
rect 25686 8191 25742 8200
rect 25700 7954 25728 8191
rect 25688 7948 25740 7954
rect 25688 7890 25740 7896
rect 25700 7546 25728 7890
rect 25688 7540 25740 7546
rect 25688 7482 25740 7488
rect 25688 5024 25740 5030
rect 25688 4966 25740 4972
rect 25240 4126 25360 4154
rect 24400 4072 24452 4078
rect 24400 4014 24452 4020
rect 25044 4072 25096 4078
rect 25044 4014 25096 4020
rect 24412 3738 24440 4014
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 24860 3732 24912 3738
rect 24860 3674 24912 3680
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 23492 3194 23520 3538
rect 23756 3460 23808 3466
rect 23756 3402 23808 3408
rect 23480 3188 23532 3194
rect 23480 3130 23532 3136
rect 23388 3120 23440 3126
rect 23388 3062 23440 3068
rect 23296 2984 23348 2990
rect 23296 2926 23348 2932
rect 23308 2582 23336 2926
rect 23296 2576 23348 2582
rect 23296 2518 23348 2524
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 22480 2310 22508 2450
rect 22468 2304 22520 2310
rect 22468 2246 22520 2252
rect 22652 2304 22704 2310
rect 22652 2246 22704 2252
rect 22480 1057 22508 2246
rect 22466 1048 22522 1057
rect 22466 983 22522 992
rect 21914 76 21916 128
rect 21968 76 21970 128
rect 21914 0 21970 76
rect 22376 128 22428 134
rect 22376 70 22428 76
rect 22664 82 22692 2246
rect 22742 82 22798 480
rect 22664 54 22798 82
rect 23400 82 23428 3062
rect 23768 3058 23796 3402
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 23664 2848 23716 2854
rect 23664 2790 23716 2796
rect 23676 2394 23704 2790
rect 23768 2514 23796 2994
rect 23848 2916 23900 2922
rect 23848 2858 23900 2864
rect 23756 2508 23808 2514
rect 23756 2450 23808 2456
rect 23860 2394 23888 2858
rect 23952 2582 23980 2994
rect 24872 2854 24900 3674
rect 24952 3664 25004 3670
rect 24952 3606 25004 3612
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 23940 2576 23992 2582
rect 23940 2518 23992 2524
rect 23676 2366 23888 2394
rect 23952 2310 23980 2518
rect 23940 2304 23992 2310
rect 23940 2246 23992 2252
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24872 1193 24900 2790
rect 24964 2514 24992 3606
rect 25240 3534 25268 4126
rect 25412 3936 25464 3942
rect 25412 3878 25464 3884
rect 25228 3528 25280 3534
rect 25228 3470 25280 3476
rect 25134 3088 25190 3097
rect 25134 3023 25190 3032
rect 25148 2990 25176 3023
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 25240 2582 25268 3470
rect 25228 2576 25280 2582
rect 25228 2518 25280 2524
rect 24952 2508 25004 2514
rect 24952 2450 25004 2456
rect 24858 1184 24914 1193
rect 24858 1119 24914 1128
rect 23478 82 23534 480
rect 23400 54 23534 82
rect 22742 0 22798 54
rect 23478 0 23534 54
rect 24306 128 24362 480
rect 24306 76 24308 128
rect 24360 76 24362 128
rect 24306 0 24362 76
rect 25134 82 25190 480
rect 25424 82 25452 3878
rect 25134 54 25452 82
rect 25700 82 25728 4966
rect 25870 82 25926 480
rect 26252 134 26280 12815
rect 27632 12782 27660 12815
rect 27620 12776 27672 12782
rect 27620 12718 27672 12724
rect 27618 9072 27674 9081
rect 27618 9007 27674 9016
rect 27632 6633 27660 9007
rect 27618 6624 27674 6633
rect 27618 6559 27674 6568
rect 26792 6384 26844 6390
rect 26792 6326 26844 6332
rect 25700 54 25926 82
rect 26240 128 26292 134
rect 26240 70 26292 76
rect 26698 82 26754 480
rect 26804 82 26832 6326
rect 27158 4040 27214 4049
rect 27158 3975 27214 3984
rect 27172 649 27200 3975
rect 27158 640 27214 649
rect 27158 575 27214 584
rect 25134 0 25190 54
rect 25870 0 25926 54
rect 26698 54 26832 82
rect 27526 128 27582 480
rect 27526 76 27528 128
rect 27580 76 27582 128
rect 26698 0 26754 54
rect 27526 0 27582 76
<< via2 >>
rect 24950 26832 25006 26888
rect 24766 25744 24822 25800
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 27618 25336 27674 25392
rect 24122 23704 24178 23760
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 16394 22616 16450 22672
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 12714 14320 12770 14376
rect 6182 13232 6238 13288
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 6090 12144 6146 12200
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 3054 11736 3110 11792
rect 2962 6976 3018 7032
rect 2502 3712 2558 3768
rect 4158 11192 4214 11248
rect 5998 11192 6054 11248
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5078 10648 5134 10704
rect 4526 8472 4582 8528
rect 3698 3168 3754 3224
rect 4250 2352 4306 2408
rect 4158 176 4214 232
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5354 4664 5410 4720
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5262 3712 5318 3768
rect 5170 720 5226 776
rect 5078 448 5134 504
rect 4986 312 5042 368
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5446 2896 5502 2952
rect 5998 2624 6054 2680
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6090 2216 6146 2272
rect 5998 1536 6054 1592
rect 8022 13640 8078 13696
rect 6642 12960 6698 13016
rect 7010 12688 7066 12744
rect 6734 9968 6790 10024
rect 6826 8472 6882 8528
rect 6550 3304 6606 3360
rect 6550 1264 6606 1320
rect 7654 9152 7710 9208
rect 7286 8608 7342 8664
rect 7102 5208 7158 5264
rect 7378 5072 7434 5128
rect 7654 3440 7710 3496
rect 7470 3168 7526 3224
rect 7286 992 7342 1048
rect 7102 40 7158 96
rect 7838 9424 7894 9480
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 8298 12824 8354 12880
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10782 9832 10838 9888
rect 8114 9016 8170 9072
rect 7838 3168 7894 3224
rect 8390 7792 8446 7848
rect 8298 7656 8354 7712
rect 9310 8880 9366 8936
rect 9954 8744 10010 8800
rect 8666 5072 8722 5128
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10690 8064 10746 8120
rect 9126 6704 9182 6760
rect 9310 6704 9366 6760
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 9494 6568 9550 6624
rect 10506 6296 10562 6352
rect 9034 5752 9090 5808
rect 8206 3984 8262 4040
rect 8942 4528 8998 4584
rect 8758 3576 8814 3632
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 9678 4664 9734 4720
rect 9954 4664 10010 4720
rect 8022 1672 8078 1728
rect 8942 3032 8998 3088
rect 10138 4120 10194 4176
rect 9586 3032 9642 3088
rect 8298 2488 8354 2544
rect 8758 1672 8814 1728
rect 8390 1128 8446 1184
rect 8206 856 8262 912
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10138 3712 10194 3768
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 12990 9696 13046 9752
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 13358 9696 13414 9752
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14554 12824 14610 12880
rect 13542 9560 13598 9616
rect 14278 9560 14334 9616
rect 13910 8744 13966 8800
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 20994 23024 21050 23080
rect 16670 15000 16726 15056
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 23662 22616 23718 22672
rect 23294 21936 23350 21992
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 16486 14320 16542 14376
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 21546 16496 21602 16552
rect 20166 13776 20222 13832
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19154 13368 19210 13424
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14646 9696 14702 9752
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14646 8608 14702 8664
rect 14370 8064 14426 8120
rect 14002 7656 14058 7712
rect 11978 2896 12034 2952
rect 12806 3304 12862 3360
rect 13634 4528 13690 4584
rect 14554 6568 14610 6624
rect 14646 6160 14702 6216
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14830 7828 14832 7848
rect 14832 7828 14884 7848
rect 14884 7828 14886 7848
rect 14830 7792 14886 7828
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15290 6296 15346 6352
rect 14646 3440 14702 3496
rect 14278 2352 14334 2408
rect 13910 1536 13966 1592
rect 14738 2216 14794 2272
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 18602 12688 18658 12744
rect 18234 11736 18290 11792
rect 17498 10648 17554 10704
rect 16302 6704 16358 6760
rect 15658 5752 15714 5808
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15382 3984 15438 4040
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15290 1672 15346 1728
rect 16670 6840 16726 6896
rect 16026 4664 16082 4720
rect 17590 1264 17646 1320
rect 17866 5072 17922 5128
rect 18510 9968 18566 10024
rect 18602 9696 18658 9752
rect 18418 312 18474 368
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 20534 12144 20590 12200
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19430 8880 19486 8936
rect 22282 11192 22338 11248
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 22466 11056 22522 11112
rect 22374 9424 22430 9480
rect 18970 4120 19026 4176
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20258 4392 20314 4448
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20902 3576 20958 3632
rect 20994 2896 21050 2952
rect 21178 2896 21234 2952
rect 20626 2352 20682 2408
rect 21730 2488 21786 2544
rect 22834 11872 22890 11928
rect 23110 15408 23166 15464
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 25134 23024 25190 23080
rect 24858 22616 24914 22672
rect 24582 21936 24638 21992
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24766 21664 24822 21720
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24766 20576 24822 20632
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24766 19488 24822 19544
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24214 15000 24270 15056
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24306 13368 24362 13424
rect 24214 13232 24270 13288
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 23754 9832 23810 9888
rect 24030 8472 24086 8528
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 25410 18536 25466 18592
rect 25318 11328 25374 11384
rect 25778 17448 25834 17504
rect 25778 14320 25834 14376
rect 25778 13640 25834 13696
rect 26238 12824 26294 12880
rect 27618 12824 27674 12880
rect 25778 10240 25834 10296
rect 25318 9560 25374 9616
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24214 8336 24270 8392
rect 21362 1672 21418 1728
rect 21178 992 21234 1048
rect 20902 856 20958 912
rect 20258 176 20314 232
rect 23570 5208 23626 5264
rect 22466 3712 22522 3768
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 25226 5072 25282 5128
rect 25134 4800 25190 4856
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 25778 9152 25834 9208
rect 25686 8200 25742 8256
rect 22466 992 22522 1048
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25134 3032 25190 3088
rect 24858 1128 24914 1184
rect 27618 9016 27674 9072
rect 27618 6568 27674 6624
rect 27158 3984 27214 4040
rect 27158 584 27214 640
<< metal3 >>
rect 27520 27344 28000 27464
rect 24945 26890 25011 26893
rect 27662 26890 27722 27344
rect 24945 26888 27722 26890
rect 24945 26832 24950 26888
rect 25006 26832 27722 26888
rect 24945 26830 27722 26832
rect 24945 26827 25011 26830
rect 27520 26256 28000 26376
rect 24761 25802 24827 25805
rect 27662 25802 27722 26256
rect 24761 25800 27722 25802
rect 24761 25744 24766 25800
rect 24822 25744 27722 25800
rect 24761 25742 27722 25744
rect 24761 25739 24827 25742
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 27520 25392 28000 25424
rect 27520 25336 27618 25392
rect 27674 25336 28000 25392
rect 27520 25304 28000 25336
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 27520 24308 28000 24336
rect 27520 24244 27660 24308
rect 27724 24244 28000 24308
rect 27520 24216 28000 24244
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 24117 23762 24183 23765
rect 27654 23762 27660 23764
rect 24117 23760 27660 23762
rect 24117 23704 24122 23760
rect 24178 23704 27660 23760
rect 24117 23702 27660 23704
rect 24117 23699 24183 23702
rect 27654 23700 27660 23702
rect 27724 23700 27730 23764
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 27520 23128 28000 23248
rect 20989 23082 21055 23085
rect 25129 23082 25195 23085
rect 20989 23080 25195 23082
rect 20989 23024 20994 23080
rect 21050 23024 25134 23080
rect 25190 23024 25195 23080
rect 20989 23022 25195 23024
rect 20989 23019 21055 23022
rect 25129 23019 25195 23022
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 16389 22674 16455 22677
rect 23657 22674 23723 22677
rect 16389 22672 23723 22674
rect 16389 22616 16394 22672
rect 16450 22616 23662 22672
rect 23718 22616 23723 22672
rect 16389 22614 23723 22616
rect 16389 22611 16455 22614
rect 23657 22611 23723 22614
rect 24853 22674 24919 22677
rect 27662 22674 27722 23128
rect 24853 22672 27722 22674
rect 24853 22616 24858 22672
rect 24914 22616 27722 22672
rect 24853 22614 27722 22616
rect 24853 22611 24919 22614
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 27520 22176 28000 22296
rect 23289 21994 23355 21997
rect 24577 21994 24643 21997
rect 23289 21992 24643 21994
rect 23289 21936 23294 21992
rect 23350 21936 24582 21992
rect 24638 21936 24643 21992
rect 23289 21934 24643 21936
rect 23289 21931 23355 21934
rect 24577 21931 24643 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 24761 21722 24827 21725
rect 27662 21722 27722 22176
rect 24761 21720 27722 21722
rect 24761 21664 24766 21720
rect 24822 21664 27722 21720
rect 24761 21662 27722 21664
rect 24761 21659 24827 21662
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 27520 21088 28000 21208
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 24761 20634 24827 20637
rect 27662 20634 27722 21088
rect 24761 20632 27722 20634
rect 24761 20576 24766 20632
rect 24822 20576 27722 20632
rect 24761 20574 27722 20576
rect 24761 20571 24827 20574
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 27520 20000 28000 20120
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 24761 19546 24827 19549
rect 27662 19546 27722 20000
rect 24761 19544 27722 19546
rect 24761 19488 24766 19544
rect 24822 19488 27722 19544
rect 24761 19486 27722 19488
rect 24761 19483 24827 19486
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19168
rect 19610 19007 19930 19008
rect 25405 18594 25471 18597
rect 27662 18594 27722 19048
rect 25405 18592 27722 18594
rect 25405 18536 25410 18592
rect 25466 18536 27722 18592
rect 25405 18534 27722 18536
rect 25405 18531 25471 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 18080
rect 19610 17919 19930 17920
rect 25773 17506 25839 17509
rect 27662 17506 27722 17960
rect 25773 17504 27722 17506
rect 25773 17448 25778 17504
rect 25834 17448 27722 17504
rect 25773 17446 27722 17448
rect 25773 17443 25839 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 27520 17008 28000 17128
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 21541 16554 21607 16557
rect 27662 16554 27722 17008
rect 21541 16552 27722 16554
rect 21541 16496 21546 16552
rect 21602 16496 27722 16552
rect 21541 16494 27722 16496
rect 21541 16491 21607 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 27520 15920 28000 16040
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 23105 15466 23171 15469
rect 27662 15466 27722 15920
rect 23105 15464 27722 15466
rect 23105 15408 23110 15464
rect 23166 15408 27722 15464
rect 23105 15406 27722 15408
rect 23105 15403 23171 15406
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 16665 15058 16731 15061
rect 24209 15058 24275 15061
rect 16665 15056 24275 15058
rect 16665 15000 16670 15056
rect 16726 15000 24214 15056
rect 24270 15000 24275 15056
rect 16665 14998 24275 15000
rect 16665 14995 16731 14998
rect 24209 14995 24275 14998
rect 27520 14832 28000 14952
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 12709 14378 12775 14381
rect 16481 14378 16547 14381
rect 12709 14376 16547 14378
rect 12709 14320 12714 14376
rect 12770 14320 16486 14376
rect 16542 14320 16547 14376
rect 12709 14318 16547 14320
rect 12709 14315 12775 14318
rect 16481 14315 16547 14318
rect 25773 14378 25839 14381
rect 27662 14378 27722 14832
rect 25773 14376 27722 14378
rect 25773 14320 25778 14376
rect 25834 14320 27722 14376
rect 25773 14318 27722 14320
rect 25773 14315 25839 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 27520 13880 28000 14000
rect 20161 13834 20227 13837
rect 9630 13832 20227 13834
rect 9630 13776 20166 13832
rect 20222 13776 20227 13832
rect 9630 13774 20227 13776
rect 8017 13698 8083 13701
rect 9630 13698 9690 13774
rect 20161 13771 20227 13774
rect 8017 13696 9690 13698
rect 8017 13640 8022 13696
rect 8078 13640 9690 13696
rect 8017 13638 9690 13640
rect 25773 13698 25839 13701
rect 27662 13698 27722 13880
rect 25773 13696 27722 13698
rect 25773 13640 25778 13696
rect 25834 13640 27722 13696
rect 25773 13638 27722 13640
rect 8017 13635 8083 13638
rect 25773 13635 25839 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 19149 13426 19215 13429
rect 24301 13426 24367 13429
rect 19149 13424 24367 13426
rect 19149 13368 19154 13424
rect 19210 13368 24306 13424
rect 24362 13368 24367 13424
rect 19149 13366 24367 13368
rect 19149 13363 19215 13366
rect 24301 13363 24367 13366
rect 6177 13290 6243 13293
rect 24209 13290 24275 13293
rect 6177 13288 24275 13290
rect 6177 13232 6182 13288
rect 6238 13232 24214 13288
rect 24270 13232 24275 13288
rect 6177 13230 24275 13232
rect 6177 13227 6243 13230
rect 24209 13227 24275 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 6637 13018 6703 13021
rect 6637 13016 14842 13018
rect 6637 12960 6642 13016
rect 6698 12960 14842 13016
rect 6637 12958 14842 12960
rect 6637 12955 6703 12958
rect 8293 12882 8359 12885
rect 14549 12882 14615 12885
rect 8293 12880 14615 12882
rect 8293 12824 8298 12880
rect 8354 12824 14554 12880
rect 14610 12824 14615 12880
rect 8293 12822 14615 12824
rect 14782 12882 14842 12958
rect 26233 12882 26299 12885
rect 14782 12880 26299 12882
rect 14782 12824 26238 12880
rect 26294 12824 26299 12880
rect 14782 12822 26299 12824
rect 8293 12819 8359 12822
rect 14549 12819 14615 12822
rect 26233 12819 26299 12822
rect 27520 12880 28000 12912
rect 27520 12824 27618 12880
rect 27674 12824 28000 12880
rect 27520 12792 28000 12824
rect 7005 12746 7071 12749
rect 18597 12746 18663 12749
rect 7005 12744 18663 12746
rect 7005 12688 7010 12744
rect 7066 12688 18602 12744
rect 18658 12688 18663 12744
rect 7005 12686 18663 12688
rect 7005 12683 7071 12686
rect 18597 12683 18663 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 6085 12202 6151 12205
rect 20529 12202 20595 12205
rect 6085 12200 20595 12202
rect 6085 12144 6090 12200
rect 6146 12144 20534 12200
rect 20590 12144 20595 12200
rect 6085 12142 20595 12144
rect 6085 12139 6151 12142
rect 20529 12139 20595 12142
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 22686 11868 22692 11932
rect 22756 11930 22762 11932
rect 22829 11930 22895 11933
rect 22756 11928 22895 11930
rect 22756 11872 22834 11928
rect 22890 11872 22895 11928
rect 22756 11870 22895 11872
rect 22756 11868 22762 11870
rect 22829 11867 22895 11870
rect 3049 11794 3115 11797
rect 18229 11794 18295 11797
rect 3049 11792 18295 11794
rect 3049 11736 3054 11792
rect 3110 11736 18234 11792
rect 18290 11736 18295 11792
rect 3049 11734 18295 11736
rect 3049 11731 3115 11734
rect 18229 11731 18295 11734
rect 27520 11704 28000 11824
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 25313 11386 25379 11389
rect 27662 11386 27722 11704
rect 25313 11384 27722 11386
rect 25313 11328 25318 11384
rect 25374 11328 27722 11384
rect 25313 11326 27722 11328
rect 25313 11323 25379 11326
rect 4153 11250 4219 11253
rect 4286 11250 4292 11252
rect 4153 11248 4292 11250
rect 4153 11192 4158 11248
rect 4214 11192 4292 11248
rect 4153 11190 4292 11192
rect 4153 11187 4219 11190
rect 4286 11188 4292 11190
rect 4356 11188 4362 11252
rect 5993 11250 6059 11253
rect 5993 11248 13830 11250
rect 5993 11192 5998 11248
rect 6054 11192 13830 11248
rect 5993 11190 13830 11192
rect 5993 11187 6059 11190
rect 13770 11114 13830 11190
rect 16430 11188 16436 11252
rect 16500 11250 16506 11252
rect 22277 11250 22343 11253
rect 16500 11248 22343 11250
rect 16500 11192 22282 11248
rect 22338 11192 22343 11248
rect 16500 11190 22343 11192
rect 16500 11188 16506 11190
rect 22277 11187 22343 11190
rect 22461 11114 22527 11117
rect 13770 11112 22527 11114
rect 13770 11056 22466 11112
rect 22522 11056 22527 11112
rect 13770 11054 22527 11056
rect 22461 11051 22527 11054
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 27520 10752 28000 10872
rect 5073 10706 5139 10709
rect 17493 10706 17559 10709
rect 5073 10704 17559 10706
rect 5073 10648 5078 10704
rect 5134 10648 17498 10704
rect 17554 10648 17559 10704
rect 5073 10646 17559 10648
rect 5073 10643 5139 10646
rect 17493 10643 17559 10646
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 25773 10298 25839 10301
rect 27662 10298 27722 10752
rect 25773 10296 27722 10298
rect 25773 10240 25778 10296
rect 25834 10240 27722 10296
rect 25773 10238 27722 10240
rect 25773 10235 25839 10238
rect 6729 10026 6795 10029
rect 18505 10026 18571 10029
rect 6729 10024 18571 10026
rect 6729 9968 6734 10024
rect 6790 9968 18510 10024
rect 18566 9968 18571 10024
rect 6729 9966 18571 9968
rect 6729 9963 6795 9966
rect 18505 9963 18571 9966
rect 10777 9890 10843 9893
rect 10910 9890 10916 9892
rect 10777 9888 10916 9890
rect 10777 9832 10782 9888
rect 10838 9832 10916 9888
rect 10777 9830 10916 9832
rect 10777 9827 10843 9830
rect 10910 9828 10916 9830
rect 10980 9828 10986 9892
rect 23422 9828 23428 9892
rect 23492 9890 23498 9892
rect 23749 9890 23815 9893
rect 23492 9888 23815 9890
rect 23492 9832 23754 9888
rect 23810 9832 23815 9888
rect 23492 9830 23815 9832
rect 23492 9828 23498 9830
rect 23749 9827 23815 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 12985 9754 13051 9757
rect 13353 9754 13419 9757
rect 14641 9754 14707 9757
rect 12985 9752 14707 9754
rect 12985 9696 12990 9752
rect 13046 9696 13358 9752
rect 13414 9696 14646 9752
rect 14702 9696 14707 9752
rect 12985 9694 14707 9696
rect 12985 9691 13051 9694
rect 13353 9691 13419 9694
rect 14641 9691 14707 9694
rect 18597 9754 18663 9757
rect 18597 9752 23490 9754
rect 18597 9696 18602 9752
rect 18658 9696 23490 9752
rect 18597 9694 23490 9696
rect 18597 9691 18663 9694
rect 13537 9618 13603 9621
rect 14273 9618 14339 9621
rect 13537 9616 14339 9618
rect 13537 9560 13542 9616
rect 13598 9560 14278 9616
rect 14334 9560 14339 9616
rect 13537 9558 14339 9560
rect 23430 9618 23490 9694
rect 27520 9664 28000 9784
rect 25313 9618 25379 9621
rect 23430 9616 25379 9618
rect 23430 9560 25318 9616
rect 25374 9560 25379 9616
rect 23430 9558 25379 9560
rect 13537 9555 13603 9558
rect 14273 9555 14339 9558
rect 25313 9555 25379 9558
rect 7833 9482 7899 9485
rect 22369 9482 22435 9485
rect 7833 9480 22435 9482
rect 7833 9424 7838 9480
rect 7894 9424 22374 9480
rect 22430 9424 22435 9480
rect 7833 9422 22435 9424
rect 7833 9419 7899 9422
rect 22369 9419 22435 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 7649 9210 7715 9213
rect 7782 9210 7788 9212
rect 7649 9208 7788 9210
rect 7649 9152 7654 9208
rect 7710 9152 7788 9208
rect 7649 9150 7788 9152
rect 7649 9147 7715 9150
rect 7782 9148 7788 9150
rect 7852 9148 7858 9212
rect 25773 9210 25839 9213
rect 27662 9210 27722 9664
rect 25773 9208 27722 9210
rect 25773 9152 25778 9208
rect 25834 9152 27722 9208
rect 25773 9150 27722 9152
rect 25773 9147 25839 9150
rect 8109 9074 8175 9077
rect 27613 9074 27679 9077
rect 8109 9072 27679 9074
rect 8109 9016 8114 9072
rect 8170 9016 27618 9072
rect 27674 9016 27679 9072
rect 8109 9014 27679 9016
rect 8109 9011 8175 9014
rect 27613 9011 27679 9014
rect 9305 8938 9371 8941
rect 19425 8938 19491 8941
rect 9305 8936 19491 8938
rect 9305 8880 9310 8936
rect 9366 8880 19430 8936
rect 19486 8880 19491 8936
rect 9305 8878 19491 8880
rect 9305 8875 9371 8878
rect 19425 8875 19491 8878
rect 9949 8802 10015 8805
rect 13905 8802 13971 8805
rect 9949 8800 13971 8802
rect 9949 8744 9954 8800
rect 10010 8744 13910 8800
rect 13966 8744 13971 8800
rect 9949 8742 13971 8744
rect 9949 8739 10015 8742
rect 13905 8739 13971 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 27520 8712 28000 8832
rect 24277 8671 24597 8672
rect 7281 8666 7347 8669
rect 14641 8666 14707 8669
rect 7281 8664 14707 8666
rect 7281 8608 7286 8664
rect 7342 8608 14646 8664
rect 14702 8608 14707 8664
rect 7281 8606 14707 8608
rect 7281 8603 7347 8606
rect 14641 8603 14707 8606
rect 4521 8530 4587 8533
rect 4654 8530 4660 8532
rect 4521 8528 4660 8530
rect 4521 8472 4526 8528
rect 4582 8472 4660 8528
rect 4521 8470 4660 8472
rect 4521 8467 4587 8470
rect 4654 8468 4660 8470
rect 4724 8468 4730 8532
rect 6821 8530 6887 8533
rect 6821 8528 13830 8530
rect 6821 8472 6826 8528
rect 6882 8472 13830 8528
rect 6821 8470 13830 8472
rect 6821 8467 6887 8470
rect 13770 8394 13830 8470
rect 23422 8468 23428 8532
rect 23492 8530 23498 8532
rect 24025 8530 24091 8533
rect 23492 8528 24091 8530
rect 23492 8472 24030 8528
rect 24086 8472 24091 8528
rect 23492 8470 24091 8472
rect 23492 8468 23498 8470
rect 24025 8467 24091 8470
rect 24209 8394 24275 8397
rect 13770 8392 24275 8394
rect 13770 8336 24214 8392
rect 24270 8336 24275 8392
rect 13770 8334 24275 8336
rect 24209 8331 24275 8334
rect 25681 8258 25747 8261
rect 27662 8258 27722 8712
rect 25681 8256 27722 8258
rect 25681 8200 25686 8256
rect 25742 8200 27722 8256
rect 25681 8198 27722 8200
rect 25681 8195 25747 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 10685 8122 10751 8125
rect 14365 8122 14431 8125
rect 10685 8120 14431 8122
rect 10685 8064 10690 8120
rect 10746 8064 14370 8120
rect 14426 8064 14431 8120
rect 10685 8062 14431 8064
rect 10685 8059 10751 8062
rect 14365 8059 14431 8062
rect 8385 7850 8451 7853
rect 14825 7850 14891 7853
rect 8385 7848 14891 7850
rect 8385 7792 8390 7848
rect 8446 7792 14830 7848
rect 14886 7792 14891 7848
rect 8385 7790 14891 7792
rect 8385 7787 8451 7790
rect 14825 7787 14891 7790
rect 8293 7714 8359 7717
rect 13997 7714 14063 7717
rect 8293 7712 14063 7714
rect 8293 7656 8298 7712
rect 8354 7656 14002 7712
rect 14058 7656 14063 7712
rect 8293 7654 14063 7656
rect 8293 7651 8359 7654
rect 13997 7651 14063 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27520 7624 28000 7744
rect 24277 7583 24597 7584
rect 18638 7244 18644 7308
rect 18708 7306 18714 7308
rect 27662 7306 27722 7624
rect 18708 7246 27722 7306
rect 18708 7244 18714 7246
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 2957 7034 3023 7037
rect 2957 7032 4170 7034
rect 2957 6976 2962 7032
rect 3018 6976 4170 7032
rect 2957 6974 4170 6976
rect 2957 6971 3023 6974
rect 4110 6898 4170 6974
rect 16665 6898 16731 6901
rect 4110 6896 16731 6898
rect 4110 6840 16670 6896
rect 16726 6840 16731 6896
rect 4110 6838 16731 6840
rect 16665 6835 16731 6838
rect 9121 6762 9187 6765
rect 9305 6762 9371 6765
rect 16297 6762 16363 6765
rect 9121 6760 16363 6762
rect 9121 6704 9126 6760
rect 9182 6704 9310 6760
rect 9366 6704 16302 6760
rect 16358 6704 16363 6760
rect 9121 6702 16363 6704
rect 9121 6699 9187 6702
rect 9305 6699 9371 6702
rect 16297 6699 16363 6702
rect 9489 6626 9555 6629
rect 14549 6626 14615 6629
rect 9489 6624 14615 6626
rect 9489 6568 9494 6624
rect 9550 6568 14554 6624
rect 14610 6568 14615 6624
rect 9489 6566 14615 6568
rect 9489 6563 9555 6566
rect 14549 6563 14615 6566
rect 27520 6624 28000 6656
rect 27520 6568 27618 6624
rect 27674 6568 28000 6624
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 27520 6536 28000 6568
rect 24277 6495 24597 6496
rect 10501 6354 10567 6357
rect 15285 6354 15351 6357
rect 10501 6352 15351 6354
rect 10501 6296 10506 6352
rect 10562 6296 15290 6352
rect 15346 6296 15351 6352
rect 10501 6294 15351 6296
rect 10501 6291 10567 6294
rect 15285 6291 15351 6294
rect 14641 6218 14707 6221
rect 14641 6216 27722 6218
rect 14641 6160 14646 6216
rect 14702 6160 27722 6216
rect 14641 6158 27722 6160
rect 14641 6155 14707 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 9029 5810 9095 5813
rect 15653 5810 15719 5813
rect 9029 5808 15719 5810
rect 9029 5752 9034 5808
rect 9090 5752 15658 5808
rect 15714 5752 15719 5808
rect 9029 5750 15719 5752
rect 9029 5747 9095 5750
rect 15653 5747 15719 5750
rect 27662 5704 27722 6158
rect 27520 5584 28000 5704
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 7097 5266 7163 5269
rect 23565 5266 23631 5269
rect 7097 5264 23631 5266
rect 7097 5208 7102 5264
rect 7158 5208 23570 5264
rect 23626 5208 23631 5264
rect 7097 5206 23631 5208
rect 7097 5203 7163 5206
rect 23565 5203 23631 5206
rect 7373 5130 7439 5133
rect 8518 5130 8524 5132
rect 7373 5128 8524 5130
rect 7373 5072 7378 5128
rect 7434 5072 8524 5128
rect 7373 5070 8524 5072
rect 7373 5067 7439 5070
rect 8518 5068 8524 5070
rect 8588 5068 8594 5132
rect 8661 5130 8727 5133
rect 17861 5130 17927 5133
rect 8661 5128 17927 5130
rect 8661 5072 8666 5128
rect 8722 5072 17866 5128
rect 17922 5072 17927 5128
rect 8661 5070 17927 5072
rect 8661 5067 8727 5070
rect 17861 5067 17927 5070
rect 23422 5068 23428 5132
rect 23492 5130 23498 5132
rect 25221 5130 25287 5133
rect 23492 5128 25287 5130
rect 23492 5072 25226 5128
rect 25282 5072 25287 5128
rect 23492 5070 25287 5072
rect 23492 5068 23498 5070
rect 25221 5067 25287 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 23606 4796 23612 4860
rect 23676 4858 23682 4860
rect 25129 4858 25195 4861
rect 23676 4856 25195 4858
rect 23676 4800 25134 4856
rect 25190 4800 25195 4856
rect 23676 4798 25195 4800
rect 23676 4796 23682 4798
rect 25129 4795 25195 4798
rect 5349 4722 5415 4725
rect 6862 4722 6868 4724
rect 5349 4720 6868 4722
rect 5349 4664 5354 4720
rect 5410 4664 6868 4720
rect 5349 4662 6868 4664
rect 5349 4659 5415 4662
rect 6862 4660 6868 4662
rect 6932 4660 6938 4724
rect 9673 4722 9739 4725
rect 9806 4722 9812 4724
rect 9673 4720 9812 4722
rect 9673 4664 9678 4720
rect 9734 4664 9812 4720
rect 9673 4662 9812 4664
rect 9673 4659 9739 4662
rect 9806 4660 9812 4662
rect 9876 4660 9882 4724
rect 9949 4722 10015 4725
rect 16021 4722 16087 4725
rect 9949 4720 16087 4722
rect 9949 4664 9954 4720
rect 10010 4664 16026 4720
rect 16082 4664 16087 4720
rect 9949 4662 16087 4664
rect 9949 4659 10015 4662
rect 16021 4659 16087 4662
rect 8937 4586 9003 4589
rect 13629 4586 13695 4589
rect 8937 4584 13695 4586
rect 8937 4528 8942 4584
rect 8998 4528 13634 4584
rect 13690 4528 13695 4584
rect 8937 4526 13695 4528
rect 8937 4523 9003 4526
rect 13629 4523 13695 4526
rect 27520 4496 28000 4616
rect 20110 4388 20116 4452
rect 20180 4450 20186 4452
rect 20253 4450 20319 4453
rect 20180 4448 20319 4450
rect 20180 4392 20258 4448
rect 20314 4392 20319 4448
rect 20180 4390 20319 4392
rect 20180 4388 20186 4390
rect 20253 4387 20319 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 10133 4178 10199 4181
rect 18965 4178 19031 4181
rect 10133 4176 19031 4178
rect 10133 4120 10138 4176
rect 10194 4120 18970 4176
rect 19026 4120 19031 4176
rect 10133 4118 19031 4120
rect 10133 4115 10199 4118
rect 18965 4115 19031 4118
rect 8201 4042 8267 4045
rect 15377 4042 15443 4045
rect 8201 4040 15443 4042
rect 8201 3984 8206 4040
rect 8262 3984 15382 4040
rect 15438 3984 15443 4040
rect 8201 3982 15443 3984
rect 8201 3979 8267 3982
rect 15377 3979 15443 3982
rect 27153 4042 27219 4045
rect 27662 4042 27722 4496
rect 27153 4040 27722 4042
rect 27153 3984 27158 4040
rect 27214 3984 27722 4040
rect 27153 3982 27722 3984
rect 27153 3979 27219 3982
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 2497 3770 2563 3773
rect 2630 3770 2636 3772
rect 2497 3768 2636 3770
rect 2497 3712 2502 3768
rect 2558 3712 2636 3768
rect 2497 3710 2636 3712
rect 2497 3707 2563 3710
rect 2630 3708 2636 3710
rect 2700 3708 2706 3772
rect 5257 3770 5323 3773
rect 10133 3770 10199 3773
rect 5257 3768 10199 3770
rect 5257 3712 5262 3768
rect 5318 3712 10138 3768
rect 10194 3712 10199 3768
rect 5257 3710 10199 3712
rect 5257 3707 5323 3710
rect 10133 3707 10199 3710
rect 20110 3708 20116 3772
rect 20180 3770 20186 3772
rect 22461 3770 22527 3773
rect 20180 3768 22527 3770
rect 20180 3712 22466 3768
rect 22522 3712 22527 3768
rect 20180 3710 22527 3712
rect 20180 3708 20186 3710
rect 22461 3707 22527 3710
rect 8753 3634 8819 3637
rect 20897 3634 20963 3637
rect 8753 3632 20963 3634
rect 8753 3576 8758 3632
rect 8814 3576 20902 3632
rect 20958 3576 20963 3632
rect 8753 3574 20963 3576
rect 8753 3571 8819 3574
rect 20897 3571 20963 3574
rect 7649 3498 7715 3501
rect 14641 3498 14707 3501
rect 7649 3496 14707 3498
rect 7649 3440 7654 3496
rect 7710 3440 14646 3496
rect 14702 3440 14707 3496
rect 7649 3438 14707 3440
rect 7649 3435 7715 3438
rect 14641 3435 14707 3438
rect 27520 3408 28000 3528
rect 6545 3362 6611 3365
rect 12801 3362 12867 3365
rect 6545 3360 12867 3362
rect 6545 3304 6550 3360
rect 6606 3304 12806 3360
rect 12862 3304 12867 3360
rect 6545 3302 12867 3304
rect 6545 3299 6611 3302
rect 12801 3299 12867 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 3693 3226 3759 3229
rect 3918 3226 3924 3228
rect 3693 3224 3924 3226
rect 3693 3168 3698 3224
rect 3754 3168 3924 3224
rect 3693 3166 3924 3168
rect 3693 3163 3759 3166
rect 3918 3164 3924 3166
rect 3988 3164 3994 3228
rect 7465 3226 7531 3229
rect 7598 3226 7604 3228
rect 7465 3224 7604 3226
rect 7465 3168 7470 3224
rect 7526 3168 7604 3224
rect 7465 3166 7604 3168
rect 7465 3163 7531 3166
rect 7598 3164 7604 3166
rect 7668 3164 7674 3228
rect 7833 3226 7899 3229
rect 7833 3224 14842 3226
rect 7833 3168 7838 3224
rect 7894 3168 14842 3224
rect 7833 3166 14842 3168
rect 7833 3163 7899 3166
rect 8937 3090 9003 3093
rect 9070 3090 9076 3092
rect 8937 3088 9076 3090
rect 8937 3032 8942 3088
rect 8998 3032 9076 3088
rect 8937 3030 9076 3032
rect 8937 3027 9003 3030
rect 9070 3028 9076 3030
rect 9140 3028 9146 3092
rect 9581 3090 9647 3093
rect 14782 3090 14842 3166
rect 25129 3090 25195 3093
rect 9581 3088 13830 3090
rect 9581 3032 9586 3088
rect 9642 3032 13830 3088
rect 9581 3030 13830 3032
rect 14782 3088 25195 3090
rect 14782 3032 25134 3088
rect 25190 3032 25195 3088
rect 14782 3030 25195 3032
rect 9581 3027 9647 3030
rect 5441 2954 5507 2957
rect 11973 2954 12039 2957
rect 5441 2952 12039 2954
rect 5441 2896 5446 2952
rect 5502 2896 11978 2952
rect 12034 2896 12039 2952
rect 5441 2894 12039 2896
rect 13770 2954 13830 3030
rect 25129 3027 25195 3030
rect 20989 2954 21055 2957
rect 13770 2952 21055 2954
rect 13770 2896 20994 2952
rect 21050 2896 21055 2952
rect 13770 2894 21055 2896
rect 5441 2891 5507 2894
rect 11973 2891 12039 2894
rect 20989 2891 21055 2894
rect 21173 2954 21239 2957
rect 27662 2954 27722 3408
rect 21173 2952 27722 2954
rect 21173 2896 21178 2952
rect 21234 2896 27722 2952
rect 21173 2894 27722 2896
rect 21173 2891 21239 2894
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 5993 2682 6059 2685
rect 9990 2682 9996 2684
rect 5993 2680 9996 2682
rect 5993 2624 5998 2680
rect 6054 2624 9996 2680
rect 5993 2622 9996 2624
rect 5993 2619 6059 2622
rect 9990 2620 9996 2622
rect 10060 2620 10066 2684
rect 8293 2546 8359 2549
rect 21725 2546 21791 2549
rect 8293 2544 21791 2546
rect 8293 2488 8298 2544
rect 8354 2488 21730 2544
rect 21786 2488 21791 2544
rect 8293 2486 21791 2488
rect 8293 2483 8359 2486
rect 21725 2483 21791 2486
rect 27520 2548 28000 2576
rect 27520 2484 27660 2548
rect 27724 2484 28000 2548
rect 27520 2456 28000 2484
rect 4245 2410 4311 2413
rect 14273 2410 14339 2413
rect 4245 2408 14339 2410
rect 4245 2352 4250 2408
rect 4306 2352 14278 2408
rect 14334 2352 14339 2408
rect 4245 2350 14339 2352
rect 4245 2347 4311 2350
rect 14273 2347 14339 2350
rect 20478 2348 20484 2412
rect 20548 2410 20554 2412
rect 20621 2410 20687 2413
rect 20548 2408 20687 2410
rect 20548 2352 20626 2408
rect 20682 2352 20687 2408
rect 20548 2350 20687 2352
rect 20548 2348 20554 2350
rect 20621 2347 20687 2350
rect 6085 2274 6151 2277
rect 14733 2274 14799 2277
rect 6085 2272 14799 2274
rect 6085 2216 6090 2272
rect 6146 2216 14738 2272
rect 14794 2216 14799 2272
rect 6085 2214 14799 2216
rect 6085 2211 6151 2214
rect 14733 2211 14799 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 8017 1730 8083 1733
rect 8150 1730 8156 1732
rect 8017 1728 8156 1730
rect 8017 1672 8022 1728
rect 8078 1672 8156 1728
rect 8017 1670 8156 1672
rect 8017 1667 8083 1670
rect 8150 1668 8156 1670
rect 8220 1668 8226 1732
rect 8753 1730 8819 1733
rect 15285 1730 15351 1733
rect 8753 1728 15351 1730
rect 8753 1672 8758 1728
rect 8814 1672 15290 1728
rect 15346 1672 15351 1728
rect 8753 1670 15351 1672
rect 8753 1667 8819 1670
rect 15285 1667 15351 1670
rect 21214 1668 21220 1732
rect 21284 1730 21290 1732
rect 21357 1730 21423 1733
rect 21284 1728 21423 1730
rect 21284 1672 21362 1728
rect 21418 1672 21423 1728
rect 21284 1670 21423 1672
rect 21284 1668 21290 1670
rect 21357 1667 21423 1670
rect 5993 1594 6059 1597
rect 13905 1594 13971 1597
rect 5993 1592 13971 1594
rect 5993 1536 5998 1592
rect 6054 1536 13910 1592
rect 13966 1536 13971 1592
rect 5993 1534 13971 1536
rect 5993 1531 6059 1534
rect 13905 1531 13971 1534
rect 27520 1368 28000 1488
rect 6545 1322 6611 1325
rect 17585 1322 17651 1325
rect 6545 1320 17651 1322
rect 6545 1264 6550 1320
rect 6606 1264 17590 1320
rect 17646 1264 17651 1320
rect 6545 1262 17651 1264
rect 6545 1259 6611 1262
rect 17585 1259 17651 1262
rect 8385 1186 8451 1189
rect 24853 1186 24919 1189
rect 8385 1184 24919 1186
rect 8385 1128 8390 1184
rect 8446 1128 24858 1184
rect 24914 1128 24919 1184
rect 8385 1126 24919 1128
rect 8385 1123 8451 1126
rect 24853 1123 24919 1126
rect 7281 1050 7347 1053
rect 21173 1050 21239 1053
rect 7281 1048 21239 1050
rect 7281 992 7286 1048
rect 7342 992 21178 1048
rect 21234 992 21239 1048
rect 7281 990 21239 992
rect 7281 987 7347 990
rect 21173 987 21239 990
rect 22318 988 22324 1052
rect 22388 1050 22394 1052
rect 22461 1050 22527 1053
rect 22388 1048 22527 1050
rect 22388 992 22466 1048
rect 22522 992 22527 1048
rect 22388 990 22527 992
rect 22388 988 22394 990
rect 22461 987 22527 990
rect 8201 914 8267 917
rect 20897 914 20963 917
rect 8201 912 20963 914
rect 8201 856 8206 912
rect 8262 856 20902 912
rect 20958 856 20963 912
rect 8201 854 20963 856
rect 8201 851 8267 854
rect 20897 851 20963 854
rect 5165 778 5231 781
rect 27662 778 27722 1368
rect 5165 776 27722 778
rect 5165 720 5170 776
rect 5226 720 27722 776
rect 5165 718 27722 720
rect 5165 715 5231 718
rect 27153 642 27219 645
rect 13770 640 27219 642
rect 13770 584 27158 640
rect 27214 584 27219 640
rect 13770 582 27219 584
rect 5073 506 5139 509
rect 13770 506 13830 582
rect 27153 579 27219 582
rect 5073 504 13830 506
rect 5073 448 5078 504
rect 5134 448 13830 504
rect 5073 446 13830 448
rect 5073 443 5139 446
rect 27520 416 28000 536
rect 4981 370 5047 373
rect 18413 370 18479 373
rect 4981 368 18479 370
rect 4981 312 4986 368
rect 5042 312 18418 368
rect 18474 312 18479 368
rect 4981 310 18479 312
rect 4981 307 5047 310
rect 18413 307 18479 310
rect 4153 234 4219 237
rect 20253 234 20319 237
rect 4153 232 20319 234
rect 4153 176 4158 232
rect 4214 176 20258 232
rect 20314 176 20319 232
rect 4153 174 20319 176
rect 4153 171 4219 174
rect 20253 171 20319 174
rect 7097 98 7163 101
rect 27662 98 27722 416
rect 7097 96 27722 98
rect 7097 40 7102 96
rect 7158 40 27722 96
rect 7097 38 27722 40
rect 7097 35 7163 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 27660 24244 27724 24308
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 27660 23700 27724 23764
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 22692 11868 22756 11932
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 4292 11188 4356 11252
rect 16436 11188 16500 11252
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 10916 9828 10980 9892
rect 23428 9828 23492 9892
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 7788 9148 7852 9212
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 4660 8468 4724 8532
rect 23428 8468 23492 8532
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 18644 7244 18708 7308
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 8524 5068 8588 5132
rect 23428 5068 23492 5132
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 23612 4796 23676 4860
rect 6868 4660 6932 4724
rect 9812 4660 9876 4724
rect 20116 4388 20180 4452
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 2636 3708 2700 3772
rect 20116 3708 20180 3772
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 3924 3164 3988 3228
rect 7604 3164 7668 3228
rect 9076 3028 9140 3092
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 9996 2620 10060 2684
rect 27660 2484 27724 2548
rect 20484 2348 20548 2412
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 8156 1668 8220 1732
rect 21220 1668 21284 1732
rect 22324 988 22388 1052
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 9814 4725 9874 11782
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 27659 24308 27725 24309
rect 27659 24244 27660 24308
rect 27724 24244 27725 24308
rect 27659 24243 27725 24244
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 27662 23765 27722 24243
rect 27659 23764 27725 23765
rect 27659 23700 27660 23764
rect 27724 23700 27725 23764
rect 27659 23699 27725 23700
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 6867 4724 6933 4725
rect 6867 4660 6868 4724
rect 6932 4660 6933 4724
rect 6867 4659 6933 4660
rect 9811 4724 9877 4725
rect 9811 4660 9812 4724
rect 9876 4660 9877 4724
rect 9811 4659 9877 4660
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 3926 3229 3986 4302
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 3923 3228 3989 3229
rect 3923 3164 3924 3228
rect 3988 3164 3989 3228
rect 3923 3163 3989 3164
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 6870 458 6930 4659
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 7603 3228 7669 3229
rect 7603 3164 7604 3228
rect 7668 3164 7669 3228
rect 7603 3163 7669 3164
rect 7606 2498 7666 3163
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 9995 2684 10061 2685
rect 9995 2620 9996 2684
rect 10060 2620 10061 2684
rect 9995 2619 10061 2620
rect 9998 1138 10058 2619
rect 10277 2128 10597 2688
rect 14944 8736 15264 9760
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 18646 7309 18706 9062
rect 19610 8192 19930 9216
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 18643 7308 18709 7309
rect 18643 7244 18644 7308
rect 18708 7244 18709 7308
rect 18643 7243 18709 7244
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 23611 4860 23677 4861
rect 23611 4796 23612 4860
rect 23676 4796 23677 4860
rect 23611 4795 23677 4796
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 23614 3178 23674 4795
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 2208 24597 3232
rect 27659 2548 27725 2549
rect 27659 2484 27660 2548
rect 27724 2484 27725 2548
rect 27659 2483 27725 2484
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 27662 458 27722 2483
<< via4 >>
rect 4206 11252 4442 11338
rect 4206 11188 4292 11252
rect 4292 11188 4356 11252
rect 4356 11188 4442 11252
rect 4206 11102 4442 11188
rect 9726 11782 9962 12018
rect 7702 9212 7938 9298
rect 7702 9148 7788 9212
rect 7788 9148 7852 9212
rect 7852 9148 7938 9212
rect 7702 9062 7938 9148
rect 4574 8532 4810 8618
rect 4574 8468 4660 8532
rect 4660 8468 4724 8532
rect 4724 8468 4810 8532
rect 4574 8382 4810 8468
rect 3838 4302 4074 4538
rect 8438 5132 8674 5218
rect 8438 5068 8524 5132
rect 8524 5068 8588 5132
rect 8588 5068 8674 5132
rect 8438 4982 8674 5068
rect 22606 11932 22842 12018
rect 22606 11868 22692 11932
rect 22692 11868 22756 11932
rect 22756 11868 22842 11932
rect 22606 11782 22842 11868
rect 16350 11252 16586 11338
rect 16350 11188 16436 11252
rect 16436 11188 16500 11252
rect 16500 11188 16586 11252
rect 16350 11102 16586 11188
rect 10830 9892 11066 9978
rect 10830 9828 10916 9892
rect 10916 9828 10980 9892
rect 10980 9828 11066 9892
rect 10830 9742 11066 9828
rect 2550 3772 2786 3858
rect 2550 3708 2636 3772
rect 2636 3708 2700 3772
rect 2700 3708 2786 3772
rect 2550 3622 2786 3708
rect 8990 3092 9226 3178
rect 8990 3028 9076 3092
rect 9076 3028 9140 3092
rect 9140 3028 9226 3092
rect 8990 2942 9226 3028
rect 7518 2262 7754 2498
rect 8070 1732 8306 1818
rect 8070 1668 8156 1732
rect 8156 1668 8220 1732
rect 8220 1668 8306 1732
rect 8070 1582 8306 1668
rect 18558 9062 18794 9298
rect 23342 9892 23578 9978
rect 23342 9828 23428 9892
rect 23428 9828 23492 9892
rect 23492 9828 23578 9892
rect 23342 9742 23578 9828
rect 23342 8532 23578 8618
rect 23342 8468 23428 8532
rect 23428 8468 23492 8532
rect 23492 8468 23578 8532
rect 23342 8382 23578 8468
rect 23342 5132 23578 5218
rect 23342 5068 23428 5132
rect 23428 5068 23492 5132
rect 23492 5068 23578 5132
rect 23342 4982 23578 5068
rect 20030 4452 20266 4538
rect 20030 4388 20116 4452
rect 20116 4388 20180 4452
rect 20180 4388 20266 4452
rect 20030 4302 20266 4388
rect 20030 3772 20266 3858
rect 20030 3708 20116 3772
rect 20116 3708 20180 3772
rect 20180 3708 20266 3772
rect 20030 3622 20266 3708
rect 23526 2942 23762 3178
rect 20398 2412 20634 2498
rect 20398 2348 20484 2412
rect 20484 2348 20548 2412
rect 20548 2348 20634 2412
rect 20398 2262 20634 2348
rect 21134 1732 21370 1818
rect 21134 1668 21220 1732
rect 21220 1668 21284 1732
rect 21284 1668 21370 1732
rect 21134 1582 21370 1668
rect 9910 902 10146 1138
rect 22238 1052 22474 1138
rect 22238 988 22324 1052
rect 22324 988 22388 1052
rect 22388 988 22474 1052
rect 22238 902 22474 988
rect 6782 222 7018 458
rect 27574 222 27810 458
<< metal5 >>
rect 9684 12018 22884 12060
rect 9684 11782 9726 12018
rect 9962 11782 22606 12018
rect 22842 11782 22884 12018
rect 9684 11740 22884 11782
rect 4164 11338 16628 11380
rect 4164 11102 4206 11338
rect 4442 11102 16350 11338
rect 16586 11102 16628 11338
rect 4164 11060 16628 11102
rect 10788 9978 23620 10020
rect 10788 9742 10830 9978
rect 11066 9742 23342 9978
rect 23578 9742 23620 9978
rect 10788 9700 23620 9742
rect 7660 9298 18836 9340
rect 7660 9062 7702 9298
rect 7938 9062 18558 9298
rect 18794 9062 18836 9298
rect 7660 9020 18836 9062
rect 4532 8618 23620 8660
rect 4532 8382 4574 8618
rect 4810 8382 23342 8618
rect 23578 8382 23620 8618
rect 4532 8340 23620 8382
rect 8396 5218 23620 5260
rect 8396 4982 8438 5218
rect 8674 4982 23342 5218
rect 23578 4982 23620 5218
rect 8396 4940 23620 4982
rect 3796 4538 20308 4580
rect 3796 4302 3838 4538
rect 4074 4302 20030 4538
rect 20266 4302 20308 4538
rect 3796 4260 20308 4302
rect 2508 3858 20308 3900
rect 2508 3622 2550 3858
rect 2786 3622 20030 3858
rect 20266 3622 20308 3858
rect 2508 3580 20308 3622
rect 8948 3178 23804 3220
rect 8948 2942 8990 3178
rect 9226 2942 23526 3178
rect 23762 2942 23804 3178
rect 8948 2900 23804 2942
rect 7476 2498 20676 2540
rect 7476 2262 7518 2498
rect 7754 2262 20398 2498
rect 20634 2262 20676 2498
rect 7476 2220 20676 2262
rect 8028 1818 21412 1860
rect 8028 1582 8070 1818
rect 8306 1582 21134 1818
rect 21370 1582 21412 1818
rect 8028 1540 21412 1582
rect 9868 1138 22516 1180
rect 9868 902 9910 1138
rect 10146 902 22238 1138
rect 22474 902 22516 1138
rect 9868 860 22516 902
rect 6740 458 27852 500
rect 6740 222 6782 458
rect 7018 222 27574 458
rect 27810 222 27852 458
rect 6740 180 27852 222
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_10 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_18
timestamp 1586364061
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_14
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_17
timestamp 1586364061
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_25
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_21
timestamp 1586364061
transform 1 0 3036 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_1_29
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_29
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _199_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_1_62 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_60 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_68
timestamp 1586364061
transform 1 0 7360 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_68
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_80
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_nand2_4  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_90
timestamp 1586364061
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_97
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_115
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_111
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _242_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_139
timestamp 1586364061
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_152
timestamp 1586364061
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_156
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_169
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_176
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_180
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 2720
box -38 -48 866 592
use scs8hd_or2_4  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_203
timestamp 1586364061
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_207
timestamp 1586364061
transform 1 0 20148 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_199
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_212
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_226
timestamp 1586364061
transform 1 0 21896 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_230
timestamp 1586364061
transform 1 0 22264 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_234
timestamp 1586364061
transform 1 0 22632 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_239
timestamp 1586364061
transform 1 0 23092 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_254
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_260
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use scs8hd_conb_1  _211_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_266
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_270
timestamp 1586364061
transform 1 0 25944 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_276
timestamp 1586364061
transform 1 0 26496 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_2_39
timestamp 1586364061
transform 1 0 4692 0 -1 3808
box -38 -48 406 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_43
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_46
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_50
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_4  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_73
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_96
timestamp 1586364061
transform 1 0 9936 0 -1 3808
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10948 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_104
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_118
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_122
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_2_137
timestamp 1586364061
transform 1 0 13708 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 13892 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_158
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_169
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_2_175
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_189
timestamp 1586364061
transform 1 0 18492 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_193
timestamp 1586364061
transform 1 0 18860 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_226
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 23276 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  FILLER_2_238
timestamp 1586364061
transform 1 0 23000 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 24288 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_250
timestamp 1586364061
transform 1 0 24104 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_254
timestamp 1586364061
transform 1 0 24472 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_267
timestamp 1586364061
transform 1 0 25668 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_6
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_10
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2668 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_16
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_20
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_24
timestamp 1586364061
transform 1 0 3312 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_35
timestamp 1586364061
transform 1 0 4324 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_42
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_46
timestamp 1586364061
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 314 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_80
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_84
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_97
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_101
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _159_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12604 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_134
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_151
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_168
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_172
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_180
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 130 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_195
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_199
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_206
timestamp 1586364061
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_210
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_225
timestamp 1586364061
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_229
timestamp 1586364061
transform 1 0 22172 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 23920 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_236
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 774 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 25484 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 26036 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_273
timestamp 1586364061
transform 1 0 26220 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_8  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_52
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_4_67
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 590 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_104
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_108
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_4  FILLER_4_121
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_127
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_132
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_or4_4  _157_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 17020 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_167
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_171
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_182
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_191
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_204
timestamp 1586364061
transform 1 0 19872 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_212
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_219
timestamp 1586364061
transform 1 0 21252 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_223
timestamp 1586364061
transform 1 0 21620 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_226
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23276 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_238
timestamp 1586364061
transform 1 0 23000 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_243
timestamp 1586364061
transform 1 0 23460 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24932 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_257
timestamp 1586364061
transform 1 0 24748 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_261
timestamp 1586364061
transform 1 0 25116 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_273
timestamp 1586364061
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_42
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_46
timestamp 1586364061
transform 1 0 5336 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_73
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_77
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_90
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_94
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_107
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_115
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_119
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 130 592
use scs8hd_or4_4  _153_
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_139
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use scs8hd_nand2_4  _138_
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_160
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_177
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 590 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 18492 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_187
timestamp 1586364061
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_191
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 222 592
use scs8hd_nor3_4  _168_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_212
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_216
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21712 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21528 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_235
timestamp 1586364061
transform 1 0 22724 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_260
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_266
timestamp 1586364061
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_270
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_276
timestamp 1586364061
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_52
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_67
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_67
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 314 592
use scs8hd_or4_4  _166_
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_72
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_72
timestamp 1586364061
transform 1 0 7728 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_78
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_83
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 314 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_100
timestamp 1586364061
transform 1 0 10304 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_121
timestamp 1586364061
transform 1 0 12236 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_134
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_138
timestamp 1586364061
transform 1 0 13800 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 866 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_140
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_158
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_154
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_164
timestamp 1586364061
transform 1 0 16192 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 16008 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__D
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_or4_4  _160_
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_175
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_184
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_181
timestamp 1586364061
transform 1 0 17756 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_190
timestamp 1586364061
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_189
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 18768 0 1 5984
box -38 -48 222 592
use scs8hd_nor3_4  _169_
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 1234 592
use scs8hd_nor3_4  _171_
timestamp 1586364061
transform 1 0 18952 0 1 5984
box -38 -48 1234 592
use scs8hd_decap_8  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_207
timestamp 1586364061
transform 1 0 20148 0 1 5984
box -38 -48 406 592
use scs8hd_inv_8  _207_
timestamp 1586364061
transform 1 0 21436 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_219
timestamp 1586364061
transform 1 0 21252 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_213
timestamp 1586364061
transform 1 0 20700 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_230
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_228
timestamp 1586364061
transform 1 0 22080 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_239
timestamp 1586364061
transform 1 0 23092 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_236
timestamp 1586364061
transform 1 0 22816 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22908 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22908 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23276 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_250
timestamp 1586364061
transform 1 0 24104 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_258
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_267
timestamp 1586364061
transform 1 0 25668 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_266
timestamp 1586364061
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_270
timestamp 1586364061
transform 1 0 25944 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_276
timestamp 1586364061
transform 1 0 26496 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_66
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 406 592
use scs8hd_buf_1  _098_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_73
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_77
timestamp 1586364061
transform 1 0 8188 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 9752 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_103
timestamp 1586364061
transform 1 0 10580 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_8_122
timestamp 1586364061
transform 1 0 12328 0 -1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_127
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_139
timestamp 1586364061
transform 1 0 13892 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_143
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_146
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_150
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 866 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_157
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_174
timestamp 1586364061
transform 1 0 17112 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 17848 0 -1 7072
box -38 -48 314 592
use scs8hd_nor3_4  _170_
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_185
timestamp 1586364061
transform 1 0 18124 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_189
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_226
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_230
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_234
timestamp 1586364061
transform 1 0 22632 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22908 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_246
timestamp 1586364061
transform 1 0 23736 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24472 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24288 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_250
timestamp 1586364061
transform 1 0 24104 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 774 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7728 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_90
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_97
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_101
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_119
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 406 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_140
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_or4_4  _143_
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_170
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_178
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 18216 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18676 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_189
timestamp 1586364061
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_206
timestamp 1586364061
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_210
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_223
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 590 592
use scs8hd_decap_4  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_249
timestamp 1586364061
transform 1 0 24012 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24288 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24104 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_261
timestamp 1586364061
transform 1 0 25116 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_266
timestamp 1586364061
transform 1 0 25576 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_9_274
timestamp 1586364061
transform 1 0 26312 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_73
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_4  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 10304 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_97
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_109
timestamp 1586364061
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 11684 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_113
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_128
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_132
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_171
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_179
timestamp 1586364061
transform 1 0 17572 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17664 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_10_191
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 590 592
use scs8hd_or2_4  _099_
timestamp 1586364061
transform 1 0 19412 0 -1 8160
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_212
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_4  FILLER_10_221
timestamp 1586364061
transform 1 0 21436 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21804 0 -1 8160
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_236
timestamp 1586364061
transform 1 0 22816 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_240
timestamp 1586364061
transform 1 0 23184 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_244
timestamp 1586364061
transform 1 0 23552 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_256
timestamp 1586364061
transform 1 0 24656 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_267
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_11_82
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 130 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_90
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_97
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12512 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_139
timestamp 1586364061
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_146
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_152
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use scs8hd_or4_4  _140_
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_165
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 16468 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_169
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_177
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_201
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_205
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_219
timestamp 1586364061
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_223
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_254
timestamp 1586364061
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_258
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_265
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 590 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_12_108
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 406 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 11776 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_112
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_115
timestamp 1586364061
transform 1 0 11684 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_132
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_142
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_146
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_12_167
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_180
timestamp 1586364061
transform 1 0 17664 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_184
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 774 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21252 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_230
timestamp 1586364061
transform 1 0 22264 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_234
timestamp 1586364061
transform 1 0 22632 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23000 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_247
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24564 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_264
timestamp 1586364061
transform 1 0 25392 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_272
timestamp 1586364061
transform 1 0 26128 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 590 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_122
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 590 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 13340 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 13708 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_131
timestamp 1586364061
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use scs8hd_or4_4  _126_
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_148
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_152
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_139
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_143
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _121_
timestamp 1586364061
transform 1 0 15732 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_165
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_169
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_172
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_176
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 17572 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_buf_1  _152_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_191
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_187
timestamp 1586364061
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use scs8hd_or4_4  _104_
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 866 592
use scs8hd_buf_1  _129_
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_195
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_194
timestamp 1586364061
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_201
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_212
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_227
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_231
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_226
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23276 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_238
timestamp 1586364061
transform 1 0 23000 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_260
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_250
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26036 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_265
timestamp 1586364061
transform 1 0 25484 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_273
timestamp 1586364061
transform 1 0 26220 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_267
timestamp 1586364061
transform 1 0 25668 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_70
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 590 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_126
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_130
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_151
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 130 592
use scs8hd_or4_4  _134_
timestamp 1586364061
transform 1 0 16284 0 1 10336
box -38 -48 866 592
use scs8hd_buf_1  _139_
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_157
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_161
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_174
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_178
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 222 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 17664 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_182
timestamp 1586364061
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 406 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_199
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_204
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 20516 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_213
timestamp 1586364061
transform 1 0 20700 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22632 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_228
timestamp 1586364061
transform 1 0 22080 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_258
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_265
timestamp 1586364061
transform 1 0 25484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  FILLER_16_113
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_148
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 314 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 15916 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 15548 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_159
timestamp 1586364061
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_172
timestamp 1586364061
transform 1 0 16928 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_176
timestamp 1586364061
transform 1 0 17296 0 -1 11424
box -38 -48 222 592
use scs8hd_or4_4  _115_
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_189
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_193
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use scs8hd_conb_1  _222_
timestamp 1586364061
transform 1 0 22448 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_228
timestamp 1586364061
transform 1 0 22080 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_235
timestamp 1586364061
transform 1 0 22724 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23460 0 -1 11424
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24472 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_252
timestamp 1586364061
transform 1 0 24288 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_256
timestamp 1586364061
transform 1 0 24656 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_77
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_89
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 1142 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_101
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_127
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_130
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_134
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_149
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_153
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_166
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__D
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_170
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_174
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_187
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_191
timestamp 1586364061
transform 1 0 18676 0 1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_209
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_213
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 22540 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_228
timestamp 1586364061
transform 1 0 22080 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_235
timestamp 1586364061
transform 1 0 22724 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 22908 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_239
timestamp 1586364061
transform 1 0 23092 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_258
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_265
timestamp 1586364061
transform 1 0 25484 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_74
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_78
timestamp 1586364061
transform 1 0 8280 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_90
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 774 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 11776 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_131
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_142
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_148
timestamp 1586364061
transform 1 0 14720 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_18_172
timestamp 1586364061
transform 1 0 16928 0 -1 12512
box -38 -48 590 592
use scs8hd_or4_4  _118_
timestamp 1586364061
transform 1 0 17664 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_189
timestamp 1586364061
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_193
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_229
timestamp 1586364061
transform 1 0 22172 0 -1 12512
box -38 -48 774 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 22908 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_246
timestamp 1586364061
transform 1 0 23736 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 24472 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 12052 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_121
timestamp 1586364061
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_128
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_142
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_157
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_155
timestamp 1586364061
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_162
timestamp 1586364061
transform 1 0 16008 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 15824 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_176
timestamp 1586364061
transform 1 0 17296 0 1 12512
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17940 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_181
timestamp 1586364061
transform 1 0 17756 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_185
timestamp 1586364061
transform 1 0 18124 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 19780 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_198
timestamp 1586364061
transform 1 0 19320 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_205
timestamp 1586364061
transform 1 0 19964 0 -1 13600
box -38 -48 590 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_212
timestamp 1586364061
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_216
timestamp 1586364061
transform 1 0 20976 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22540 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_231
timestamp 1586364061
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_235
timestamp 1586364061
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_228
timestamp 1586364061
transform 1 0 22080 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_241
timestamp 1586364061
transform 1 0 23276 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_239
timestamp 1586364061
transform 1 0 23092 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22908 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_245
timestamp 1586364061
transform 1 0 23644 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23460 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23828 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23828 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_256
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_260
timestamp 1586364061
transform 1 0 25024 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_258
timestamp 1586364061
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_267
timestamp 1586364061
transform 1 0 25668 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_271
timestamp 1586364061
transform 1 0 26036 0 1 12512
box -38 -48 590 592
use scs8hd_decap_4  FILLER_20_270
timestamp 1586364061
transform 1 0 25944 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_60
timestamp 1586364061
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_127
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_136
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_21_151
timestamp 1586364061
transform 1 0 14996 0 1 13600
box -38 -48 590 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_169
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_173
timestamp 1586364061
transform 1 0 17020 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19964 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19780 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_201
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_216
timestamp 1586364061
transform 1 0 20976 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21712 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_235
timestamp 1586364061
transform 1 0 22724 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22908 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_239
timestamp 1586364061
transform 1 0 23092 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_254
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_258
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_265
timestamp 1586364061
transform 1 0 25484 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_61
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_73
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_85
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_91
timestamp 1586364061
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_128
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_158
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_162
timestamp 1586364061
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_174
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17848 0 -1 14688
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_22_193
timestamp 1586364061
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use scs8hd_conb_1  _223_
timestamp 1586364061
transform 1 0 19780 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_197
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_8  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_226
timestamp 1586364061
transform 1 0 21896 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_230
timestamp 1586364061
transform 1 0 22264 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_243
timestamp 1586364061
transform 1 0 23460 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_247
timestamp 1586364061
transform 1 0 23828 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_12  FILLER_22_260
timestamp 1586364061
transform 1 0 25024 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_272
timestamp 1586364061
transform 1 0 26128 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_140
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_155
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_163
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_204
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20700 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_209
timestamp 1586364061
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_222
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_226
timestamp 1586364061
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_230
timestamp 1586364061
transform 1 0 22264 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_236
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_240
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_254
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_258
timestamp 1586364061
transform 1 0 24840 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_265
timestamp 1586364061
transform 1 0 25484 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_6  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17296 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_185
timestamp 1586364061
transform 1 0 18124 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_189
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_221
timestamp 1586364061
transform 1 0 21436 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 21528 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_233
timestamp 1586364061
transform 1 0 22540 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 24012 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_4  FILLER_24_245
timestamp 1586364061
transform 1 0 23644 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_258
timestamp 1586364061
transform 1 0 24840 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_270
timestamp 1586364061
transform 1 0 25944 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_274
timestamp 1586364061
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 590 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_141
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_145
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_149
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15180 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_162
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_166
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_170
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_25_178
timestamp 1586364061
transform 1 0 17480 0 1 15776
box -38 -48 314 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_187
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_191
timestamp 1586364061
transform 1 0 18676 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18952 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_205
timestamp 1586364061
transform 1 0 19964 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20976 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_209
timestamp 1586364061
transform 1 0 20332 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_215
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_219
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_223
timestamp 1586364061
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _172_
timestamp 1586364061
transform 1 0 24012 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 23828 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_258
timestamp 1586364061
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_262
timestamp 1586364061
transform 1 0 25208 0 1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_273
timestamp 1586364061
transform 1 0 26220 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_158
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_162
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_175
timestamp 1586364061
transform 1 0 17204 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 130 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 18768 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 18584 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 17664 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_183
timestamp 1586364061
transform 1 0 17940 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_193
timestamp 1586364061
transform 1 0 18860 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_182
timestamp 1586364061
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_198
timestamp 1586364061
transform 1 0 19320 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_206
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_6  FILLER_27_201
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_207
timestamp 1586364061
transform 1 0 20148 0 1 16864
box -38 -48 130 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_221
timestamp 1586364061
transform 1 0 21436 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_219
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 21528 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 21988 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_231
timestamp 1586364061
transform 1 0 22356 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_223
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_248
timestamp 1586364061
transform 1 0 23920 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_236
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 24656 0 -1 16864
box -38 -48 866 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 25208 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_254
timestamp 1586364061
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_258
timestamp 1586364061
transform 1 0 24840 0 1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 25760 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_265
timestamp 1586364061
transform 1 0 25484 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_273
timestamp 1586364061
transform 1 0 26220 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_266
timestamp 1586364061
transform 1 0 25576 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_270
timestamp 1586364061
transform 1 0 25944 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16192 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_162
timestamp 1586364061
transform 1 0 16008 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_167
timestamp 1586364061
transform 1 0 16468 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_179
timestamp 1586364061
transform 1 0 17572 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 17664 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_12  FILLER_28_189
timestamp 1586364061
transform 1 0 18492 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_201
timestamp 1586364061
transform 1 0 19596 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 21068 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_213
timestamp 1586364061
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 22632 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_226
timestamp 1586364061
transform 1 0 21896 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_28_243
timestamp 1586364061
transform 1 0 23460 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_12  FILLER_28_260
timestamp 1586364061
transform 1 0 25024 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_272
timestamp 1586364061
transform 1 0 26128 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _225_
timestamp 1586364061
transform 1 0 21528 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_225
timestamp 1586364061
transform 1 0 21804 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_236
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_249
timestamp 1586364061
transform 1 0 24012 0 1 17952
box -38 -48 406 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 24564 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_259
timestamp 1586364061
transform 1 0 24932 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_263
timestamp 1586364061
transform 1 0 25300 0 1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_29_275
timestamp 1586364061
transform 1 0 26404 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_conb_1  _224_
timestamp 1586364061
transform 1 0 22540 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_6  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_236
timestamp 1586364061
transform 1 0 22816 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_8  FILLER_30_247
timestamp 1586364061
transform 1 0 23828 0 -1 19040
box -38 -48 774 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 24564 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_259
timestamp 1586364061
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_271
timestamp 1586364061
transform 1 0 26036 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 25208 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_256
timestamp 1586364061
transform 1 0 24656 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_260
timestamp 1586364061
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_264
timestamp 1586364061
transform 1 0 25392 0 1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_31_276
timestamp 1586364061
transform 1 0 26496 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 24564 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_259
timestamp 1586364061
transform 1 0 24932 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_271
timestamp 1586364061
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 24564 0 -1 21216
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24196 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_254
timestamp 1586364061
transform 1 0 24472 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_258
timestamp 1586364061
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_262
timestamp 1586364061
transform 1 0 25208 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_259
timestamp 1586364061
transform 1 0 24932 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_274
timestamp 1586364061
transform 1 0 26312 0 1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_34_271
timestamp 1586364061
transform 1 0 26036 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_253
timestamp 1586364061
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_259
timestamp 1586364061
transform 1 0 24932 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_263
timestamp 1586364061
transform 1 0 25300 0 1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_35_275
timestamp 1586364061
transform 1 0 26404 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_155
timestamp 1586364061
transform 1 0 15364 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_160
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_172
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_180
timestamp 1586364061
transform 1 0 17664 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_37_192
timestamp 1586364061
transform 1 0 18768 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_197
timestamp 1586364061
transform 1 0 19228 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_209
timestamp 1586364061
transform 1 0 20332 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_221
timestamp 1586364061
transform 1 0 21436 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_233
timestamp 1586364061
transform 1 0 22540 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_241
timestamp 1586364061
transform 1 0 23276 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15640 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_161
timestamp 1586364061
transform 1 0 15916 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_173
timestamp 1586364061
transform 1 0 17020 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_185
timestamp 1586364061
transform 1 0 18124 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_193
timestamp 1586364061
transform 1 0 18860 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_198
timestamp 1586364061
transform 1 0 19320 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_210
timestamp 1586364061
transform 1 0 20424 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_259
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_271
timestamp 1586364061
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_171
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_259
timestamp 1586364061
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_271
timestamp 1586364061
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal2 s 14738 0 14794 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 15566 0 15622 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 16302 0 16358 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 17130 0 17186 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 17958 0 18014 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 18694 0 18750 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 4342 0 4398 480 6 bottom_left_grid_pin_11_
port 6 nsew default input
rlabel metal2 s 5170 0 5226 480 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal2 s 5906 0 5962 480 6 bottom_left_grid_pin_15_
port 8 nsew default input
rlabel metal2 s 386 0 442 480 6 bottom_left_grid_pin_1_
port 9 nsew default input
rlabel metal2 s 1122 0 1178 480 6 bottom_left_grid_pin_3_
port 10 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_5_
port 11 nsew default input
rlabel metal2 s 2778 0 2834 480 6 bottom_left_grid_pin_7_
port 12 nsew default input
rlabel metal2 s 3514 0 3570 480 6 bottom_left_grid_pin_9_
port 13 nsew default input
rlabel metal2 s 27526 0 27582 480 6 bottom_right_grid_pin_11_
port 14 nsew default input
rlabel metal3 s 27520 416 28000 536 6 chanx_right_in[0]
port 15 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 chanx_right_in[1]
port 16 nsew default input
rlabel metal3 s 27520 2456 28000 2576 6 chanx_right_in[2]
port 17 nsew default input
rlabel metal3 s 27520 3408 28000 3528 6 chanx_right_in[3]
port 18 nsew default input
rlabel metal3 s 27520 4496 28000 4616 6 chanx_right_in[4]
port 19 nsew default input
rlabel metal3 s 27520 5584 28000 5704 6 chanx_right_in[5]
port 20 nsew default input
rlabel metal3 s 27520 6536 28000 6656 6 chanx_right_in[6]
port 21 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_in[7]
port 22 nsew default input
rlabel metal3 s 27520 8712 28000 8832 6 chanx_right_in[8]
port 23 nsew default input
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_out[0]
port 24 nsew default tristate
rlabel metal3 s 27520 20000 28000 20120 6 chanx_right_out[1]
port 25 nsew default tristate
rlabel metal3 s 27520 21088 28000 21208 6 chanx_right_out[2]
port 26 nsew default tristate
rlabel metal3 s 27520 22176 28000 22296 6 chanx_right_out[3]
port 27 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_out[4]
port 28 nsew default tristate
rlabel metal3 s 27520 24216 28000 24336 6 chanx_right_out[5]
port 29 nsew default tristate
rlabel metal3 s 27520 25304 28000 25424 6 chanx_right_out[6]
port 30 nsew default tristate
rlabel metal3 s 27520 26256 28000 26376 6 chanx_right_out[7]
port 31 nsew default tristate
rlabel metal3 s 27520 27344 28000 27464 6 chanx_right_out[8]
port 32 nsew default tristate
rlabel metal2 s 6734 0 6790 480 6 chany_bottom_in[0]
port 33 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[1]
port 34 nsew default input
rlabel metal2 s 8298 0 8354 480 6 chany_bottom_in[2]
port 35 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[3]
port 36 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[4]
port 37 nsew default input
rlabel metal2 s 10690 0 10746 480 6 chany_bottom_in[5]
port 38 nsew default input
rlabel metal2 s 11518 0 11574 480 6 chany_bottom_in[6]
port 39 nsew default input
rlabel metal2 s 12346 0 12402 480 6 chany_bottom_in[7]
port 40 nsew default input
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_in[8]
port 41 nsew default input
rlabel metal2 s 20350 0 20406 480 6 chany_bottom_out[0]
port 42 nsew default tristate
rlabel metal2 s 21086 0 21142 480 6 chany_bottom_out[1]
port 43 nsew default tristate
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[2]
port 44 nsew default tristate
rlabel metal2 s 22742 0 22798 480 6 chany_bottom_out[3]
port 45 nsew default tristate
rlabel metal2 s 23478 0 23534 480 6 chany_bottom_out[4]
port 46 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[5]
port 47 nsew default tristate
rlabel metal2 s 25134 0 25190 480 6 chany_bottom_out[6]
port 48 nsew default tristate
rlabel metal2 s 25870 0 25926 480 6 chany_bottom_out[7]
port 49 nsew default tristate
rlabel metal2 s 26698 0 26754 480 6 chany_bottom_out[8]
port 50 nsew default tristate
rlabel metal2 s 19522 0 19578 480 6 data_in
port 51 nsew default input
rlabel metal2 s 13910 0 13966 480 6 enable
port 52 nsew default input
rlabel metal3 s 27520 17960 28000 18080 6 right_bottom_grid_pin_12_
port 53 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 right_top_grid_pin_11_
port 54 nsew default input
rlabel metal3 s 27520 15920 28000 16040 6 right_top_grid_pin_13_
port 55 nsew default input
rlabel metal3 s 27520 17008 28000 17128 6 right_top_grid_pin_15_
port 56 nsew default input
rlabel metal3 s 27520 9664 28000 9784 6 right_top_grid_pin_1_
port 57 nsew default input
rlabel metal3 s 27520 10752 28000 10872 6 right_top_grid_pin_3_
port 58 nsew default input
rlabel metal3 s 27520 11704 28000 11824 6 right_top_grid_pin_5_
port 59 nsew default input
rlabel metal3 s 27520 12792 28000 12912 6 right_top_grid_pin_7_
port 60 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 right_top_grid_pin_9_
port 61 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 63 nsew default input
<< end >>
