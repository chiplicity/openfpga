magic
tech sky130A
magscale 1 2
timestamp 1606228189
<< locali >>
rect 7205 18853 7297 18887
rect 7205 18683 7239 18853
rect 9965 18071 9999 18173
rect 6009 17527 6043 17697
rect 7021 17595 7055 17833
rect 9505 17527 9539 17765
rect 12081 17595 12115 17765
rect 7297 16575 7331 16677
rect 8585 16031 8619 16133
rect 6653 14807 6687 14909
rect 2881 14263 2915 14365
rect 13369 13923 13403 14025
rect 8861 12631 8895 12801
rect 12265 9435 12299 9605
rect 13369 9367 13403 9469
rect 8769 8823 8803 9129
rect 7757 7327 7791 7429
rect 10701 7259 10735 7429
rect 9137 6103 9171 6205
rect 9505 4539 9539 4709
rect 6837 3519 6871 3689
rect 11345 3587 11379 3689
rect 8125 2975 8159 3077
rect 10425 2839 10459 2941
rect 3801 2295 3835 2601
rect 10609 2295 10643 2601
<< viali >>
rect 3433 20009 3467 20043
rect 5825 20009 5859 20043
rect 12817 20009 12851 20043
rect 13369 20009 13403 20043
rect 16681 20009 16715 20043
rect 2513 19941 2547 19975
rect 3341 19941 3375 19975
rect 6377 19941 6411 19975
rect 9045 19941 9079 19975
rect 1685 19873 1719 19907
rect 2237 19873 2271 19907
rect 4629 19873 4663 19907
rect 5733 19873 5767 19907
rect 7185 19873 7219 19907
rect 9137 19873 9171 19907
rect 9781 19873 9815 19907
rect 10517 19873 10551 19907
rect 11345 19873 11379 19907
rect 11897 19873 11931 19907
rect 12633 19873 12667 19907
rect 13185 19873 13219 19907
rect 13737 19873 13771 19907
rect 16497 19873 16531 19907
rect 3525 19805 3559 19839
rect 4721 19805 4755 19839
rect 4905 19805 4939 19839
rect 6009 19805 6043 19839
rect 6929 19805 6963 19839
rect 9229 19805 9263 19839
rect 9965 19805 9999 19839
rect 10701 19805 10735 19839
rect 5365 19737 5399 19771
rect 8677 19737 8711 19771
rect 12081 19737 12115 19771
rect 1869 19669 1903 19703
rect 2973 19669 3007 19703
rect 4261 19669 4295 19703
rect 8309 19669 8343 19703
rect 11529 19669 11563 19703
rect 13921 19669 13955 19703
rect 6929 19465 6963 19499
rect 3525 19329 3559 19363
rect 7573 19329 7607 19363
rect 10057 19329 10091 19363
rect 1593 19261 1627 19295
rect 2145 19261 2179 19295
rect 4169 19261 4203 19295
rect 5825 19261 5859 19295
rect 7389 19261 7423 19295
rect 8401 19261 8435 19295
rect 11713 19261 11747 19295
rect 12449 19261 12483 19295
rect 14105 19261 14139 19295
rect 14657 19261 14691 19295
rect 15209 19261 15243 19295
rect 15761 19261 15795 19295
rect 16313 19261 16347 19295
rect 16865 19261 16899 19295
rect 17417 19261 17451 19295
rect 18061 19261 18095 19295
rect 18613 19261 18647 19295
rect 19165 19261 19199 19295
rect 19717 19261 19751 19295
rect 2421 19193 2455 19227
rect 3249 19193 3283 19227
rect 4436 19193 4470 19227
rect 7297 19193 7331 19227
rect 7941 19193 7975 19227
rect 8668 19193 8702 19227
rect 10302 19193 10336 19227
rect 12716 19193 12750 19227
rect 1777 19125 1811 19159
rect 2881 19125 2915 19159
rect 3341 19125 3375 19159
rect 5549 19125 5583 19159
rect 6009 19125 6043 19159
rect 9781 19125 9815 19159
rect 11437 19125 11471 19159
rect 11897 19125 11931 19159
rect 13829 19125 13863 19159
rect 14289 19125 14323 19159
rect 14841 19125 14875 19159
rect 15393 19125 15427 19159
rect 15945 19125 15979 19159
rect 16497 19125 16531 19159
rect 17049 19125 17083 19159
rect 17601 19125 17635 19159
rect 18245 19125 18279 19159
rect 18797 19125 18831 19159
rect 19349 19125 19383 19159
rect 19901 19125 19935 19159
rect 2973 18921 3007 18955
rect 3433 18921 3467 18955
rect 7113 18921 7147 18955
rect 8769 18921 8803 18955
rect 9229 18921 9263 18955
rect 9873 18921 9907 18955
rect 10333 18921 10367 18955
rect 13277 18921 13311 18955
rect 4322 18853 4356 18887
rect 6000 18853 6034 18887
rect 7297 18853 7331 18887
rect 7634 18853 7668 18887
rect 14105 18853 14139 18887
rect 15577 18853 15611 18887
rect 19073 18853 19107 18887
rect 1501 18785 1535 18819
rect 2237 18785 2271 18819
rect 3341 18785 3375 18819
rect 1777 18717 1811 18751
rect 2513 18717 2547 18751
rect 3617 18717 3651 18751
rect 4077 18717 4111 18751
rect 5733 18717 5767 18751
rect 9045 18785 9079 18819
rect 10241 18785 10275 18819
rect 11428 18785 11462 18819
rect 13185 18785 13219 18819
rect 13829 18785 13863 18819
rect 15301 18785 15335 18819
rect 18797 18785 18831 18819
rect 7389 18717 7423 18751
rect 10425 18717 10459 18751
rect 11161 18717 11195 18751
rect 13369 18717 13403 18751
rect 5457 18649 5491 18683
rect 7205 18649 7239 18683
rect 12541 18649 12575 18683
rect 12817 18581 12851 18615
rect 4169 18377 4203 18411
rect 6101 18377 6135 18411
rect 9873 18377 9907 18411
rect 10333 18377 10367 18411
rect 10793 18377 10827 18411
rect 7021 18309 7055 18343
rect 2329 18241 2363 18275
rect 8125 18241 8159 18275
rect 8493 18241 8527 18275
rect 11253 18241 11287 18275
rect 11437 18241 11471 18275
rect 11805 18241 11839 18275
rect 12633 18241 12667 18275
rect 13369 18241 13403 18275
rect 1777 18173 1811 18207
rect 2789 18173 2823 18207
rect 3056 18173 3090 18207
rect 4721 18173 4755 18207
rect 6837 18173 6871 18207
rect 8760 18173 8794 18207
rect 9965 18173 9999 18207
rect 10149 18173 10183 18207
rect 12449 18173 12483 18207
rect 13185 18173 13219 18207
rect 4966 18105 5000 18139
rect 7849 18105 7883 18139
rect 1961 18037 1995 18071
rect 7481 18037 7515 18071
rect 7941 18037 7975 18071
rect 9965 18037 9999 18071
rect 11161 18037 11195 18071
rect 4261 17833 4295 17867
rect 4813 17833 4847 17867
rect 5273 17833 5307 17867
rect 6101 17833 6135 17867
rect 7021 17833 7055 17867
rect 11989 17833 12023 17867
rect 14749 17833 14783 17867
rect 6561 17765 6595 17799
rect 1501 17697 1535 17731
rect 2053 17697 2087 17731
rect 2329 17697 2363 17731
rect 2789 17697 2823 17731
rect 4077 17697 4111 17731
rect 5181 17697 5215 17731
rect 6009 17697 6043 17731
rect 6469 17697 6503 17731
rect 2973 17629 3007 17663
rect 3525 17629 3559 17663
rect 5457 17629 5491 17663
rect 6745 17629 6779 17663
rect 9505 17765 9539 17799
rect 10876 17765 10910 17799
rect 12081 17765 12115 17799
rect 7113 17697 7147 17731
rect 7380 17697 7414 17731
rect 8769 17697 8803 17731
rect 7021 17561 7055 17595
rect 8493 17561 8527 17595
rect 9689 17697 9723 17731
rect 10609 17629 10643 17663
rect 12633 17697 12667 17731
rect 13277 17697 13311 17731
rect 14565 17697 14599 17731
rect 12725 17629 12759 17663
rect 12817 17629 12851 17663
rect 12081 17561 12115 17595
rect 12265 17561 12299 17595
rect 13461 17561 13495 17595
rect 1685 17493 1719 17527
rect 6009 17493 6043 17527
rect 8953 17493 8987 17527
rect 9505 17493 9539 17527
rect 9873 17493 9907 17527
rect 5733 17289 5767 17323
rect 8217 17289 8251 17323
rect 13645 17289 13679 17323
rect 3709 17221 3743 17255
rect 9873 17221 9907 17255
rect 1685 17153 1719 17187
rect 2421 17153 2455 17187
rect 3249 17153 3283 17187
rect 4261 17153 4295 17187
rect 5365 17153 5399 17187
rect 6377 17153 6411 17187
rect 10149 17153 10183 17187
rect 11805 17153 11839 17187
rect 1501 17085 1535 17119
rect 2237 17085 2271 17119
rect 2973 17085 3007 17119
rect 4169 17085 4203 17119
rect 6837 17085 6871 17119
rect 8493 17085 8527 17119
rect 13461 17085 13495 17119
rect 7104 17017 7138 17051
rect 8760 17017 8794 17051
rect 10394 17017 10428 17051
rect 4077 16949 4111 16983
rect 4721 16949 4755 16983
rect 5089 16949 5123 16983
rect 5181 16949 5215 16983
rect 6101 16949 6135 16983
rect 6193 16949 6227 16983
rect 11529 16949 11563 16983
rect 12449 16949 12483 16983
rect 2973 16745 3007 16779
rect 3433 16745 3467 16779
rect 7113 16745 7147 16779
rect 7389 16745 7423 16779
rect 8401 16745 8435 16779
rect 8861 16745 8895 16779
rect 10057 16745 10091 16779
rect 10885 16745 10919 16779
rect 11253 16745 11287 16779
rect 11897 16745 11931 16779
rect 12357 16745 12391 16779
rect 5978 16677 6012 16711
rect 7297 16677 7331 16711
rect 13185 16677 13219 16711
rect 1501 16609 1535 16643
rect 2053 16609 2087 16643
rect 3341 16609 3375 16643
rect 4333 16609 4367 16643
rect 7757 16609 7791 16643
rect 8769 16609 8803 16643
rect 11345 16609 11379 16643
rect 12265 16609 12299 16643
rect 12909 16609 12943 16643
rect 2237 16541 2271 16575
rect 3617 16541 3651 16575
rect 4077 16541 4111 16575
rect 5733 16541 5767 16575
rect 7297 16541 7331 16575
rect 7849 16541 7883 16575
rect 8033 16541 8067 16575
rect 8953 16541 8987 16575
rect 10149 16541 10183 16575
rect 10333 16541 10367 16575
rect 11437 16541 11471 16575
rect 12449 16541 12483 16575
rect 1685 16405 1719 16439
rect 5457 16405 5491 16439
rect 9689 16405 9723 16439
rect 3985 16201 4019 16235
rect 5641 16201 5675 16235
rect 6837 16201 6871 16235
rect 8769 16201 8803 16235
rect 13829 16201 13863 16235
rect 8585 16133 8619 16167
rect 7389 16065 7423 16099
rect 9413 16065 9447 16099
rect 11161 16065 11195 16099
rect 11805 16065 11839 16099
rect 1869 15997 1903 16031
rect 2605 15997 2639 16031
rect 4261 15997 4295 16031
rect 5917 15997 5951 16031
rect 6653 15997 6687 16031
rect 8585 15997 8619 16031
rect 9137 15997 9171 16031
rect 11621 15997 11655 16031
rect 12449 15997 12483 16031
rect 2145 15929 2179 15963
rect 2872 15929 2906 15963
rect 4528 15929 4562 15963
rect 7205 15929 7239 15963
rect 7849 15929 7883 15963
rect 8309 15929 8343 15963
rect 10977 15929 11011 15963
rect 12716 15929 12750 15963
rect 1409 15861 1443 15895
rect 6101 15861 6135 15895
rect 6469 15861 6503 15895
rect 7297 15861 7331 15895
rect 9229 15861 9263 15895
rect 10609 15861 10643 15895
rect 11069 15861 11103 15895
rect 14105 15861 14139 15895
rect 1593 15657 1627 15691
rect 2421 15657 2455 15691
rect 2973 15657 3007 15691
rect 3341 15657 3375 15691
rect 4813 15657 4847 15691
rect 5825 15657 5859 15691
rect 6285 15657 6319 15691
rect 6929 15657 6963 15691
rect 11345 15657 11379 15691
rect 11805 15657 11839 15691
rect 13737 15657 13771 15691
rect 14381 15657 14415 15691
rect 4353 15589 4387 15623
rect 6193 15589 6227 15623
rect 14473 15589 14507 15623
rect 1409 15521 1443 15555
rect 2329 15521 2363 15555
rect 4077 15521 4111 15555
rect 5181 15521 5215 15555
rect 7297 15521 7331 15555
rect 8208 15521 8242 15555
rect 9689 15521 9723 15555
rect 9945 15521 9979 15555
rect 11713 15521 11747 15555
rect 12357 15521 12391 15555
rect 12624 15521 12658 15555
rect 2513 15453 2547 15487
rect 3433 15453 3467 15487
rect 3617 15453 3651 15487
rect 5273 15453 5307 15487
rect 5457 15453 5491 15487
rect 6377 15453 6411 15487
rect 7389 15453 7423 15487
rect 7573 15453 7607 15487
rect 7941 15453 7975 15487
rect 11989 15453 12023 15487
rect 14565 15453 14599 15487
rect 14013 15385 14047 15419
rect 1961 15317 1995 15351
rect 9321 15317 9355 15351
rect 11069 15317 11103 15351
rect 1593 15113 1627 15147
rect 4353 15113 4387 15147
rect 5733 15113 5767 15147
rect 8217 15113 8251 15147
rect 9597 15113 9631 15147
rect 1961 15045 1995 15079
rect 2421 14977 2455 15011
rect 2605 14977 2639 15011
rect 5181 14977 5215 15011
rect 5365 14977 5399 15011
rect 6377 14977 6411 15011
rect 9137 14977 9171 15011
rect 10057 14977 10091 15011
rect 10241 14977 10275 15011
rect 14657 14977 14691 15011
rect 1409 14909 1443 14943
rect 2973 14909 3007 14943
rect 6193 14909 6227 14943
rect 6653 14909 6687 14943
rect 6837 14909 6871 14943
rect 10609 14909 10643 14943
rect 12449 14909 12483 14943
rect 2329 14841 2363 14875
rect 3240 14841 3274 14875
rect 6101 14841 6135 14875
rect 7104 14841 7138 14875
rect 9965 14841 9999 14875
rect 10876 14841 10910 14875
rect 12694 14841 12728 14875
rect 14473 14841 14507 14875
rect 4721 14773 4755 14807
rect 5089 14773 5123 14807
rect 6653 14773 6687 14807
rect 8585 14773 8619 14807
rect 8953 14773 8987 14807
rect 9045 14773 9079 14807
rect 11989 14773 12023 14807
rect 13829 14773 13863 14807
rect 14105 14773 14139 14807
rect 14565 14773 14599 14807
rect 2973 14569 3007 14603
rect 7021 14569 7055 14603
rect 7113 14569 7147 14603
rect 8125 14569 8159 14603
rect 9965 14569 9999 14603
rect 10977 14569 11011 14603
rect 11345 14569 11379 14603
rect 3341 14501 3375 14535
rect 6193 14501 6227 14535
rect 15669 14501 15703 14535
rect 1869 14433 1903 14467
rect 2329 14433 2363 14467
rect 4804 14433 4838 14467
rect 8033 14433 8067 14467
rect 9137 14433 9171 14467
rect 10333 14433 10367 14467
rect 10425 14433 10459 14467
rect 11161 14433 11195 14467
rect 11713 14433 11747 14467
rect 12817 14433 12851 14467
rect 12909 14433 12943 14467
rect 13176 14433 13210 14467
rect 2421 14365 2455 14399
rect 2605 14365 2639 14399
rect 2881 14365 2915 14399
rect 3433 14365 3467 14399
rect 3617 14365 3651 14399
rect 4537 14365 4571 14399
rect 7205 14365 7239 14399
rect 8309 14365 8343 14399
rect 10517 14365 10551 14399
rect 11805 14365 11839 14399
rect 11989 14365 12023 14399
rect 15761 14365 15795 14399
rect 15853 14365 15887 14399
rect 1961 14297 1995 14331
rect 6653 14297 6687 14331
rect 12633 14297 12667 14331
rect 14289 14297 14323 14331
rect 2881 14229 2915 14263
rect 5917 14229 5951 14263
rect 7665 14229 7699 14263
rect 15301 14229 15335 14263
rect 1409 14025 1443 14059
rect 7113 14025 7147 14059
rect 7757 14025 7791 14059
rect 9873 14025 9907 14059
rect 10885 14025 10919 14059
rect 12541 14025 12575 14059
rect 13369 14025 13403 14059
rect 8769 13957 8803 13991
rect 1869 13889 1903 13923
rect 2053 13889 2087 13923
rect 2421 13889 2455 13923
rect 8401 13889 8435 13923
rect 9321 13889 9355 13923
rect 10333 13889 10367 13923
rect 10517 13889 10551 13923
rect 11529 13889 11563 13923
rect 13185 13889 13219 13923
rect 13369 13889 13403 13923
rect 14105 13889 14139 13923
rect 15025 13889 15059 13923
rect 15209 13889 15243 13923
rect 1777 13821 1811 13855
rect 4445 13821 4479 13855
rect 4701 13821 4735 13855
rect 6285 13821 6319 13855
rect 7297 13821 7331 13855
rect 8125 13821 8159 13855
rect 11345 13821 11379 13855
rect 13921 13821 13955 13855
rect 2677 13753 2711 13787
rect 8217 13753 8251 13787
rect 10241 13753 10275 13787
rect 14933 13753 14967 13787
rect 3801 13685 3835 13719
rect 5825 13685 5859 13719
rect 6101 13685 6135 13719
rect 9137 13685 9171 13719
rect 9229 13685 9263 13719
rect 11253 13685 11287 13719
rect 12909 13685 12943 13719
rect 13001 13685 13035 13719
rect 13553 13685 13587 13719
rect 14013 13685 14047 13719
rect 14565 13685 14599 13719
rect 1593 13481 1627 13515
rect 2973 13481 3007 13515
rect 4537 13481 4571 13515
rect 9321 13481 9355 13515
rect 13461 13481 13495 13515
rect 14197 13481 14231 13515
rect 20545 13481 20579 13515
rect 3433 13413 3467 13447
rect 4445 13413 4479 13447
rect 5641 13413 5675 13447
rect 6438 13413 6472 13447
rect 9934 13413 9968 13447
rect 1409 13345 1443 13379
rect 2329 13345 2363 13379
rect 3341 13345 3375 13379
rect 5549 13345 5583 13379
rect 8208 13345 8242 13379
rect 11345 13345 11379 13379
rect 12081 13345 12115 13379
rect 12337 13345 12371 13379
rect 14105 13345 14139 13379
rect 19432 13345 19466 13379
rect 2421 13277 2455 13311
rect 2605 13277 2639 13311
rect 3617 13277 3651 13311
rect 4629 13277 4663 13311
rect 5825 13277 5859 13311
rect 6193 13277 6227 13311
rect 7941 13277 7975 13311
rect 9689 13277 9723 13311
rect 11621 13277 11655 13311
rect 14381 13277 14415 13311
rect 19165 13277 19199 13311
rect 4077 13209 4111 13243
rect 1961 13141 1995 13175
rect 5181 13141 5215 13175
rect 7573 13141 7607 13175
rect 11069 13141 11103 13175
rect 13737 13141 13771 13175
rect 1593 12937 1627 12971
rect 2421 12937 2455 12971
rect 3617 12937 3651 12971
rect 12081 12937 12115 12971
rect 12909 12937 12943 12971
rect 8769 12869 8803 12903
rect 2237 12801 2271 12835
rect 2973 12801 3007 12835
rect 4169 12801 4203 12835
rect 5089 12801 5123 12835
rect 5273 12801 5307 12835
rect 6193 12801 6227 12835
rect 7389 12801 7423 12835
rect 8861 12801 8895 12835
rect 9597 12801 9631 12835
rect 13277 12801 13311 12835
rect 17325 12801 17359 12835
rect 1961 12733 1995 12767
rect 6101 12733 6135 12767
rect 6837 12733 6871 12767
rect 7656 12733 7690 12767
rect 2789 12665 2823 12699
rect 4077 12665 4111 12699
rect 4997 12665 5031 12699
rect 6009 12665 6043 12699
rect 9505 12733 9539 12767
rect 10701 12733 10735 12767
rect 13093 12733 13127 12767
rect 13544 12733 13578 12767
rect 17049 12733 17083 12767
rect 10968 12665 11002 12699
rect 2053 12597 2087 12631
rect 2881 12597 2915 12631
rect 3525 12597 3559 12631
rect 3985 12597 4019 12631
rect 4629 12597 4663 12631
rect 5641 12597 5675 12631
rect 7021 12597 7055 12631
rect 8861 12597 8895 12631
rect 9045 12597 9079 12631
rect 9413 12597 9447 12631
rect 12449 12597 12483 12631
rect 14657 12597 14691 12631
rect 1501 12393 1535 12427
rect 2513 12393 2547 12427
rect 3525 12393 3559 12427
rect 6561 12393 6595 12427
rect 7573 12393 7607 12427
rect 7665 12393 7699 12427
rect 8585 12393 8619 12427
rect 9965 12393 9999 12427
rect 10977 12393 11011 12427
rect 11345 12393 11379 12427
rect 11989 12393 12023 12427
rect 12357 12393 12391 12427
rect 14933 12393 14967 12427
rect 15301 12393 15335 12427
rect 15761 12393 15795 12427
rect 2881 12325 2915 12359
rect 10333 12325 10367 12359
rect 12449 12325 12483 12359
rect 13820 12325 13854 12359
rect 1869 12257 1903 12291
rect 4445 12257 4479 12291
rect 4712 12257 4746 12291
rect 6469 12257 6503 12291
rect 8953 12257 8987 12291
rect 11437 12257 11471 12291
rect 13553 12257 13587 12291
rect 15669 12257 15703 12291
rect 1961 12189 1995 12223
rect 2145 12189 2179 12223
rect 2973 12189 3007 12223
rect 3157 12189 3191 12223
rect 6653 12189 6687 12223
rect 7757 12189 7791 12223
rect 9045 12189 9079 12223
rect 9137 12189 9171 12223
rect 10425 12189 10459 12223
rect 10609 12189 10643 12223
rect 11621 12189 11655 12223
rect 12541 12189 12575 12223
rect 15853 12189 15887 12223
rect 6101 12121 6135 12155
rect 5825 12053 5859 12087
rect 7205 12053 7239 12087
rect 1593 11849 1627 11883
rect 6193 11849 6227 11883
rect 8953 11849 8987 11883
rect 11989 11849 12023 11883
rect 14381 11849 14415 11883
rect 2513 11713 2547 11747
rect 3617 11713 3651 11747
rect 9505 11713 9539 11747
rect 13001 11713 13035 11747
rect 15209 11713 15243 11747
rect 1409 11645 1443 11679
rect 3433 11645 3467 11679
rect 3985 11645 4019 11679
rect 4813 11645 4847 11679
rect 5080 11645 5114 11679
rect 6837 11645 6871 11679
rect 7093 11645 7127 11679
rect 8677 11645 8711 11679
rect 10609 11645 10643 11679
rect 13268 11645 13302 11679
rect 2329 11577 2363 11611
rect 4261 11577 4295 11611
rect 9321 11577 9355 11611
rect 9965 11577 9999 11611
rect 10876 11577 10910 11611
rect 1961 11509 1995 11543
rect 2421 11509 2455 11543
rect 2973 11509 3007 11543
rect 3341 11509 3375 11543
rect 8217 11509 8251 11543
rect 8493 11509 8527 11543
rect 9413 11509 9447 11543
rect 14657 11509 14691 11543
rect 15025 11509 15059 11543
rect 15117 11509 15151 11543
rect 5089 11305 5123 11339
rect 5457 11305 5491 11339
rect 8585 11305 8619 11339
rect 11621 11305 11655 11339
rect 12173 11305 12207 11339
rect 13461 11305 13495 11339
rect 13829 11305 13863 11339
rect 14289 11305 14323 11339
rect 1869 11237 1903 11271
rect 4537 11237 4571 11271
rect 5549 11237 5583 11271
rect 13369 11237 13403 11271
rect 14197 11237 14231 11271
rect 1593 11169 1627 11203
rect 2596 11169 2630 11203
rect 4445 11169 4479 11203
rect 6469 11169 6503 11203
rect 6561 11169 6595 11203
rect 7297 11169 7331 11203
rect 7757 11169 7791 11203
rect 8953 11169 8987 11203
rect 9045 11169 9079 11203
rect 10333 11169 10367 11203
rect 12541 11169 12575 11203
rect 12633 11169 12667 11203
rect 2329 11101 2363 11135
rect 4629 11101 4663 11135
rect 5641 11101 5675 11135
rect 6745 11101 6779 11135
rect 7849 11101 7883 11135
rect 8033 11101 8067 11135
rect 9229 11101 9263 11135
rect 12725 11101 12759 11135
rect 13553 11101 13587 11135
rect 14381 11101 14415 11135
rect 14657 11101 14691 11135
rect 7113 11033 7147 11067
rect 13001 11033 13035 11067
rect 3709 10965 3743 10999
rect 4077 10965 4111 10999
rect 6101 10965 6135 10999
rect 7389 10965 7423 10999
rect 2789 10761 2823 10795
rect 3065 10761 3099 10795
rect 5089 10761 5123 10795
rect 9229 10761 9263 10795
rect 11069 10761 11103 10795
rect 11161 10761 11195 10795
rect 13185 10761 13219 10795
rect 6837 10693 6871 10727
rect 3617 10625 3651 10659
rect 4721 10625 4755 10659
rect 5549 10625 5583 10659
rect 5641 10625 5675 10659
rect 6101 10625 6135 10659
rect 7481 10625 7515 10659
rect 11713 10625 11747 10659
rect 13737 10625 13771 10659
rect 14749 10625 14783 10659
rect 1409 10557 1443 10591
rect 1676 10557 1710 10591
rect 3525 10557 3559 10591
rect 4537 10557 4571 10591
rect 7205 10557 7239 10591
rect 7849 10557 7883 10591
rect 8116 10557 8150 10591
rect 9413 10557 9447 10591
rect 9689 10557 9723 10591
rect 9945 10557 9979 10591
rect 11529 10557 11563 10591
rect 12817 10557 12851 10591
rect 13553 10557 13587 10591
rect 3433 10489 3467 10523
rect 14565 10489 14599 10523
rect 4077 10421 4111 10455
rect 4445 10421 4479 10455
rect 5457 10421 5491 10455
rect 7297 10421 7331 10455
rect 11621 10421 11655 10455
rect 12633 10421 12667 10455
rect 13645 10421 13679 10455
rect 14197 10421 14231 10455
rect 14657 10421 14691 10455
rect 1593 10217 1627 10251
rect 3433 10217 3467 10251
rect 4629 10217 4663 10251
rect 8861 10217 8895 10251
rect 11069 10217 11103 10251
rect 14381 10217 14415 10251
rect 5089 10149 5123 10183
rect 6070 10149 6104 10183
rect 9956 10149 9990 10183
rect 13246 10149 13280 10183
rect 1409 10081 1443 10115
rect 2044 10081 2078 10115
rect 4997 10081 5031 10115
rect 7748 10081 7782 10115
rect 11345 10081 11379 10115
rect 11601 10081 11635 10115
rect 13001 10081 13035 10115
rect 1777 10013 1811 10047
rect 5273 10013 5307 10047
rect 5825 10013 5859 10047
rect 7481 10013 7515 10047
rect 9689 10013 9723 10047
rect 7205 9945 7239 9979
rect 3157 9877 3191 9911
rect 12725 9877 12759 9911
rect 4169 9673 4203 9707
rect 6285 9673 6319 9707
rect 7849 9673 7883 9707
rect 1777 9605 1811 9639
rect 4629 9605 4663 9639
rect 6837 9605 6871 9639
rect 12265 9605 12299 9639
rect 12449 9605 12483 9639
rect 2329 9537 2363 9571
rect 7481 9537 7515 9571
rect 8401 9537 8435 9571
rect 10241 9537 10275 9571
rect 10977 9537 11011 9571
rect 11069 9537 11103 9571
rect 11805 9537 11839 9571
rect 11989 9537 12023 9571
rect 2789 9469 2823 9503
rect 4813 9469 4847 9503
rect 4905 9469 4939 9503
rect 12909 9537 12943 9571
rect 13001 9537 13035 9571
rect 14013 9537 14047 9571
rect 15025 9537 15059 9571
rect 2145 9401 2179 9435
rect 3056 9401 3090 9435
rect 5172 9401 5206 9435
rect 8217 9401 8251 9435
rect 10885 9401 10919 9435
rect 11713 9401 11747 9435
rect 12265 9401 12299 9435
rect 13369 9469 13403 9503
rect 14933 9401 14967 9435
rect 2237 9333 2271 9367
rect 7205 9333 7239 9367
rect 7297 9333 7331 9367
rect 8309 9333 8343 9367
rect 9689 9333 9723 9367
rect 10057 9333 10091 9367
rect 10149 9333 10183 9367
rect 10517 9333 10551 9367
rect 11345 9333 11379 9367
rect 12817 9333 12851 9367
rect 13369 9333 13403 9367
rect 13461 9333 13495 9367
rect 13829 9333 13863 9367
rect 13921 9333 13955 9367
rect 14473 9333 14507 9367
rect 14841 9333 14875 9367
rect 1869 9129 1903 9163
rect 4077 9129 4111 9163
rect 7113 9129 7147 9163
rect 7941 9129 7975 9163
rect 8401 9129 8435 9163
rect 8769 9129 8803 9163
rect 10977 9129 11011 9163
rect 12173 9129 12207 9163
rect 12725 9129 12759 9163
rect 13737 9129 13771 9163
rect 14105 9129 14139 9163
rect 2237 9061 2271 9095
rect 5457 9061 5491 9095
rect 6101 9061 6135 9095
rect 3249 8993 3283 9027
rect 4445 8993 4479 9027
rect 7205 8993 7239 9027
rect 8309 8993 8343 9027
rect 2329 8925 2363 8959
rect 2513 8925 2547 8959
rect 3341 8925 3375 8959
rect 3433 8925 3467 8959
rect 4537 8925 4571 8959
rect 4721 8925 4755 8959
rect 5549 8925 5583 8959
rect 5733 8925 5767 8959
rect 7389 8925 7423 8959
rect 8493 8925 8527 8959
rect 10149 9061 10183 9095
rect 13093 9061 13127 9095
rect 13185 9061 13219 9095
rect 9137 8993 9171 9027
rect 11069 8993 11103 9027
rect 12081 8993 12115 9027
rect 11161 8925 11195 8959
rect 12357 8925 12391 8959
rect 13277 8925 13311 8959
rect 14197 8925 14231 8959
rect 14289 8925 14323 8959
rect 10609 8857 10643 8891
rect 2881 8789 2915 8823
rect 5089 8789 5123 8823
rect 6745 8789 6779 8823
rect 7849 8789 7883 8823
rect 8769 8789 8803 8823
rect 8953 8789 8987 8823
rect 11713 8789 11747 8823
rect 3617 8585 3651 8619
rect 3893 8585 3927 8619
rect 6469 8585 6503 8619
rect 10057 8585 10091 8619
rect 14473 8585 14507 8619
rect 10425 8517 10459 8551
rect 12081 8517 12115 8551
rect 12449 8517 12483 8551
rect 13461 8517 13495 8551
rect 4445 8449 4479 8483
rect 5089 8449 5123 8483
rect 7021 8449 7055 8483
rect 10701 8449 10735 8483
rect 12909 8449 12943 8483
rect 13001 8449 13035 8483
rect 13921 8449 13955 8483
rect 14105 8449 14139 8483
rect 15025 8449 15059 8483
rect 1501 8381 1535 8415
rect 2237 8381 2271 8415
rect 2504 8381 2538 8415
rect 5356 8381 5390 8415
rect 8677 8381 8711 8415
rect 10609 8381 10643 8415
rect 12817 8381 12851 8415
rect 1777 8313 1811 8347
rect 4353 8313 4387 8347
rect 7288 8313 7322 8347
rect 8922 8313 8956 8347
rect 10968 8313 11002 8347
rect 4261 8245 4295 8279
rect 8401 8245 8435 8279
rect 13829 8245 13863 8279
rect 14841 8245 14875 8279
rect 14933 8245 14967 8279
rect 4077 8041 4111 8075
rect 5549 8041 5583 8075
rect 6193 8041 6227 8075
rect 6653 8041 6687 8075
rect 7757 8041 7791 8075
rect 1676 7973 1710 8007
rect 3065 7973 3099 8007
rect 4537 7973 4571 8007
rect 8125 7973 8159 8007
rect 9956 7973 9990 8007
rect 11704 7973 11738 8007
rect 4445 7905 4479 7939
rect 5641 7905 5675 7939
rect 6561 7905 6595 7939
rect 8217 7905 8251 7939
rect 11437 7905 11471 7939
rect 13093 7905 13127 7939
rect 13360 7905 13394 7939
rect 1409 7837 1443 7871
rect 4721 7837 4755 7871
rect 5825 7837 5859 7871
rect 6745 7837 6779 7871
rect 8309 7837 8343 7871
rect 8769 7837 8803 7871
rect 9689 7837 9723 7871
rect 2789 7701 2823 7735
rect 5181 7701 5215 7735
rect 11069 7701 11103 7735
rect 12817 7701 12851 7735
rect 14473 7701 14507 7735
rect 3525 7497 3559 7531
rect 6101 7497 6135 7531
rect 6837 7497 6871 7531
rect 10793 7497 10827 7531
rect 6377 7429 6411 7463
rect 7757 7429 7791 7463
rect 7849 7429 7883 7463
rect 9781 7429 9815 7463
rect 10701 7429 10735 7463
rect 3985 7361 4019 7395
rect 4077 7361 4111 7395
rect 7389 7361 7423 7395
rect 8401 7361 8435 7395
rect 10425 7361 10459 7395
rect 1869 7293 1903 7327
rect 2136 7293 2170 7327
rect 4721 7293 4755 7327
rect 6561 7293 6595 7327
rect 7297 7293 7331 7327
rect 7757 7293 7791 7327
rect 8217 7293 8251 7327
rect 10149 7293 10183 7327
rect 11437 7361 11471 7395
rect 11897 7361 11931 7395
rect 13001 7361 13035 7395
rect 14013 7361 14047 7395
rect 15025 7361 15059 7395
rect 16037 7361 16071 7395
rect 12817 7293 12851 7327
rect 13829 7293 13863 7327
rect 14841 7293 14875 7327
rect 3893 7225 3927 7259
rect 4988 7225 5022 7259
rect 8309 7225 8343 7259
rect 10701 7225 10735 7259
rect 13921 7225 13955 7259
rect 15853 7225 15887 7259
rect 15945 7225 15979 7259
rect 3249 7157 3283 7191
rect 7205 7157 7239 7191
rect 10241 7157 10275 7191
rect 11161 7157 11195 7191
rect 11253 7157 11287 7191
rect 12449 7157 12483 7191
rect 12909 7157 12943 7191
rect 13461 7157 13495 7191
rect 14473 7157 14507 7191
rect 14933 7157 14967 7191
rect 15485 7157 15519 7191
rect 3341 6953 3375 6987
rect 4445 6953 4479 6987
rect 7297 6953 7331 6987
rect 8401 6953 8435 6987
rect 11069 6953 11103 6987
rect 11805 6953 11839 6987
rect 12449 6953 12483 6987
rect 12817 6953 12851 6987
rect 6162 6885 6196 6919
rect 9956 6885 9990 6919
rect 11897 6885 11931 6919
rect 12909 6885 12943 6919
rect 2228 6817 2262 6851
rect 5181 6817 5215 6851
rect 8493 6817 8527 6851
rect 13829 6817 13863 6851
rect 13921 6817 13955 6851
rect 14749 6817 14783 6851
rect 15669 6817 15703 6851
rect 1961 6749 1995 6783
rect 4537 6749 4571 6783
rect 4721 6749 4755 6783
rect 5917 6749 5951 6783
rect 8585 6749 8619 6783
rect 9045 6749 9079 6783
rect 9689 6749 9723 6783
rect 12081 6749 12115 6783
rect 13093 6749 13127 6783
rect 14013 6749 14047 6783
rect 15761 6749 15795 6783
rect 15853 6749 15887 6783
rect 8033 6681 8067 6715
rect 4077 6613 4111 6647
rect 11437 6613 11471 6647
rect 13461 6613 13495 6647
rect 15301 6613 15335 6647
rect 3157 6409 3191 6443
rect 10885 6409 10919 6443
rect 13829 6409 13863 6443
rect 11345 6273 11379 6307
rect 11529 6273 11563 6307
rect 14105 6273 14139 6307
rect 16773 6273 16807 6307
rect 1777 6205 1811 6239
rect 4353 6205 4387 6239
rect 4620 6205 4654 6239
rect 7573 6205 7607 6239
rect 9137 6205 9171 6239
rect 9229 6205 9263 6239
rect 9496 6205 9530 6239
rect 12265 6205 12299 6239
rect 12449 6205 12483 6239
rect 14565 6205 14599 6239
rect 16681 6205 16715 6239
rect 2044 6137 2078 6171
rect 7840 6137 7874 6171
rect 12716 6137 12750 6171
rect 14832 6137 14866 6171
rect 16589 6137 16623 6171
rect 3433 6069 3467 6103
rect 5733 6069 5767 6103
rect 8953 6069 8987 6103
rect 9137 6069 9171 6103
rect 10609 6069 10643 6103
rect 11253 6069 11287 6103
rect 12081 6069 12115 6103
rect 15945 6069 15979 6103
rect 16221 6069 16255 6103
rect 2697 5865 2731 5899
rect 2789 5797 2823 5831
rect 10057 5797 10091 5831
rect 10149 5797 10183 5831
rect 4445 5729 4479 5763
rect 4537 5729 4571 5763
rect 5724 5729 5758 5763
rect 7380 5729 7414 5763
rect 11253 5729 11287 5763
rect 11509 5729 11543 5763
rect 12909 5729 12943 5763
rect 13553 5729 13587 5763
rect 13820 5729 13854 5763
rect 15301 5729 15335 5763
rect 15568 5729 15602 5763
rect 17141 5729 17175 5763
rect 18981 5729 19015 5763
rect 2973 5661 3007 5695
rect 4721 5661 4755 5695
rect 5457 5661 5491 5695
rect 7113 5661 7147 5695
rect 10333 5661 10367 5695
rect 17417 5661 17451 5695
rect 19257 5661 19291 5695
rect 6837 5593 6871 5627
rect 16681 5593 16715 5627
rect 2329 5525 2363 5559
rect 4077 5525 4111 5559
rect 8493 5525 8527 5559
rect 9689 5525 9723 5559
rect 12633 5525 12667 5559
rect 13093 5525 13127 5559
rect 14933 5525 14967 5559
rect 1869 5321 1903 5355
rect 6193 5321 6227 5355
rect 6837 5321 6871 5355
rect 13829 5321 13863 5355
rect 14841 5321 14875 5355
rect 11345 5253 11379 5287
rect 2421 5185 2455 5219
rect 3433 5185 3467 5219
rect 7389 5185 7423 5219
rect 8953 5185 8987 5219
rect 10517 5185 10551 5219
rect 10701 5185 10735 5219
rect 11805 5185 11839 5219
rect 11989 5185 12023 5219
rect 14473 5185 14507 5219
rect 15485 5185 15519 5219
rect 16313 5185 16347 5219
rect 16405 5185 16439 5219
rect 17417 5185 17451 5219
rect 2237 5117 2271 5151
rect 3249 5117 3283 5151
rect 4813 5117 4847 5151
rect 7205 5117 7239 5151
rect 8677 5117 8711 5151
rect 8769 5117 8803 5151
rect 12449 5117 12483 5151
rect 12705 5117 12739 5151
rect 13921 5117 13955 5151
rect 14289 5117 14323 5151
rect 15209 5117 15243 5151
rect 17233 5117 17267 5151
rect 19809 5117 19843 5151
rect 5080 5049 5114 5083
rect 7297 5049 7331 5083
rect 11713 5049 11747 5083
rect 17325 5049 17359 5083
rect 2329 4981 2363 5015
rect 2881 4981 2915 5015
rect 3341 4981 3375 5015
rect 8309 4981 8343 5015
rect 10057 4981 10091 5015
rect 10425 4981 10459 5015
rect 14105 4981 14139 5015
rect 15301 4981 15335 5015
rect 15853 4981 15887 5015
rect 16221 4981 16255 5015
rect 16865 4981 16899 5015
rect 19993 4981 20027 5015
rect 4077 4777 4111 4811
rect 5549 4777 5583 4811
rect 6561 4777 6595 4811
rect 7021 4777 7055 4811
rect 7573 4777 7607 4811
rect 10241 4777 10275 4811
rect 11621 4777 11655 4811
rect 11713 4777 11747 4811
rect 13921 4777 13955 4811
rect 14381 4777 14415 4811
rect 15301 4777 15335 4811
rect 15761 4777 15795 4811
rect 16313 4777 16347 4811
rect 5917 4709 5951 4743
rect 8953 4709 8987 4743
rect 9505 4709 9539 4743
rect 9781 4709 9815 4743
rect 16773 4709 16807 4743
rect 1593 4641 1627 4675
rect 1860 4641 1894 4675
rect 4445 4641 4479 4675
rect 6929 4641 6963 4675
rect 7941 4641 7975 4675
rect 9045 4641 9079 4675
rect 3341 4573 3375 4607
rect 3433 4573 3467 4607
rect 4537 4573 4571 4607
rect 4721 4573 4755 4607
rect 6009 4573 6043 4607
rect 6193 4573 6227 4607
rect 7113 4573 7147 4607
rect 8033 4573 8067 4607
rect 8217 4573 8251 4607
rect 9229 4573 9263 4607
rect 10609 4641 10643 4675
rect 10701 4641 10735 4675
rect 12541 4641 12575 4675
rect 12808 4641 12842 4675
rect 15669 4641 15703 4675
rect 16681 4641 16715 4675
rect 17969 4641 18003 4675
rect 10885 4573 10919 4607
rect 11897 4573 11931 4607
rect 14473 4573 14507 4607
rect 14657 4573 14691 4607
rect 15853 4573 15887 4607
rect 16865 4573 16899 4607
rect 9505 4505 9539 4539
rect 14013 4505 14047 4539
rect 2973 4437 3007 4471
rect 8585 4437 8619 4471
rect 11253 4437 11287 4471
rect 18153 4437 18187 4471
rect 6837 4233 6871 4267
rect 12449 4165 12483 4199
rect 16957 4165 16991 4199
rect 1777 4097 1811 4131
rect 4077 4097 4111 4131
rect 4261 4097 4295 4131
rect 7481 4097 7515 4131
rect 8493 4097 8527 4131
rect 10057 4097 10091 4131
rect 10977 4097 11011 4131
rect 13001 4097 13035 4131
rect 14013 4097 14047 4131
rect 14749 4097 14783 4131
rect 15761 4097 15795 4131
rect 2044 4029 2078 4063
rect 4629 4029 4663 4063
rect 7297 4029 7331 4063
rect 8217 4029 8251 4063
rect 9781 4029 9815 4063
rect 10793 4029 10827 4063
rect 10885 4029 10919 4063
rect 11621 4029 11655 4063
rect 11897 4029 11931 4063
rect 14565 4029 14599 4063
rect 15669 4029 15703 4063
rect 16221 4029 16255 4063
rect 16773 4029 16807 4063
rect 3985 3961 4019 3995
rect 4896 3961 4930 3995
rect 12817 3961 12851 3995
rect 14657 3961 14691 3995
rect 3157 3893 3191 3927
rect 3617 3893 3651 3927
rect 6009 3893 6043 3927
rect 6285 3893 6319 3927
rect 7205 3893 7239 3927
rect 7849 3893 7883 3927
rect 8309 3893 8343 3927
rect 9413 3893 9447 3927
rect 9873 3893 9907 3927
rect 10425 3893 10459 3927
rect 12909 3893 12943 3927
rect 14197 3893 14231 3927
rect 15209 3893 15243 3927
rect 15577 3893 15611 3927
rect 16405 3893 16439 3927
rect 1961 3689 1995 3723
rect 3341 3689 3375 3723
rect 6837 3689 6871 3723
rect 8401 3689 8435 3723
rect 11253 3689 11287 3723
rect 11345 3689 11379 3723
rect 12909 3689 12943 3723
rect 14197 3689 14231 3723
rect 14657 3689 14691 3723
rect 6377 3621 6411 3655
rect 2329 3553 2363 3587
rect 3433 3553 3467 3587
rect 4425 3553 4459 3587
rect 13553 3621 13587 3655
rect 13645 3621 13679 3655
rect 7288 3553 7322 3587
rect 9045 3553 9079 3587
rect 10129 3553 10163 3587
rect 11345 3553 11379 3587
rect 11785 3553 11819 3587
rect 14565 3553 14599 3587
rect 15301 3553 15335 3587
rect 15577 3553 15611 3587
rect 16037 3553 16071 3587
rect 16589 3553 16623 3587
rect 17141 3553 17175 3587
rect 2421 3485 2455 3519
rect 2605 3485 2639 3519
rect 3525 3485 3559 3519
rect 4169 3485 4203 3519
rect 6469 3485 6503 3519
rect 6653 3485 6687 3519
rect 6837 3485 6871 3519
rect 7021 3485 7055 3519
rect 9873 3485 9907 3519
rect 11529 3485 11563 3519
rect 13737 3485 13771 3519
rect 14749 3485 14783 3519
rect 5549 3417 5583 3451
rect 13185 3417 13219 3451
rect 16773 3417 16807 3451
rect 2973 3349 3007 3383
rect 6009 3349 6043 3383
rect 9229 3349 9263 3383
rect 16221 3349 16255 3383
rect 17325 3349 17359 3383
rect 4721 3145 4755 3179
rect 9689 3145 9723 3179
rect 10149 3145 10183 3179
rect 15669 3145 15703 3179
rect 8125 3077 8159 3111
rect 10517 3077 10551 3111
rect 12449 3077 12483 3111
rect 14473 3077 14507 3111
rect 16589 3077 16623 3111
rect 2421 3009 2455 3043
rect 2605 3009 2639 3043
rect 2973 3009 3007 3043
rect 5365 3009 5399 3043
rect 6377 3009 6411 3043
rect 7757 3009 7791 3043
rect 7941 3009 7975 3043
rect 10977 3009 11011 3043
rect 11161 3009 11195 3043
rect 13001 3009 13035 3043
rect 14105 3009 14139 3043
rect 15025 3009 15059 3043
rect 2329 2941 2363 2975
rect 3229 2941 3263 2975
rect 5089 2941 5123 2975
rect 6193 2941 6227 2975
rect 8125 2941 8159 2975
rect 8309 2941 8343 2975
rect 8565 2941 8599 2975
rect 9965 2941 9999 2975
rect 10425 2941 10459 2975
rect 10885 2941 10919 2975
rect 11621 2941 11655 2975
rect 13829 2941 13863 2975
rect 13921 2941 13955 2975
rect 15485 2941 15519 2975
rect 16405 2941 16439 2975
rect 16957 2941 16991 2975
rect 18429 2941 18463 2975
rect 7665 2873 7699 2907
rect 11897 2873 11931 2907
rect 12909 2873 12943 2907
rect 14933 2873 14967 2907
rect 1961 2805 1995 2839
rect 4353 2805 4387 2839
rect 5181 2805 5215 2839
rect 5733 2805 5767 2839
rect 6101 2805 6135 2839
rect 7297 2805 7331 2839
rect 10425 2805 10459 2839
rect 12817 2805 12851 2839
rect 13461 2805 13495 2839
rect 14841 2805 14875 2839
rect 17141 2805 17175 2839
rect 18613 2805 18647 2839
rect 1961 2601 1995 2635
rect 3433 2601 3467 2635
rect 3801 2601 3835 2635
rect 4077 2601 4111 2635
rect 5549 2601 5583 2635
rect 10241 2601 10275 2635
rect 10609 2601 10643 2635
rect 11161 2601 11195 2635
rect 11253 2601 11287 2635
rect 13001 2601 13035 2635
rect 14841 2601 14875 2635
rect 15669 2601 15703 2635
rect 2329 2465 2363 2499
rect 3341 2465 3375 2499
rect 2421 2397 2455 2431
rect 2605 2397 2639 2431
rect 3617 2397 3651 2431
rect 2973 2329 3007 2363
rect 4445 2533 4479 2567
rect 7481 2533 7515 2567
rect 9045 2533 9079 2567
rect 10149 2533 10183 2567
rect 5457 2465 5491 2499
rect 4537 2397 4571 2431
rect 4629 2397 4663 2431
rect 5641 2397 5675 2431
rect 7573 2397 7607 2431
rect 7757 2397 7791 2431
rect 9137 2397 9171 2431
rect 9321 2397 9355 2431
rect 10333 2397 10367 2431
rect 7113 2329 7147 2363
rect 8677 2329 8711 2363
rect 13093 2533 13127 2567
rect 11805 2465 11839 2499
rect 14013 2465 14047 2499
rect 14105 2465 14139 2499
rect 14657 2465 14691 2499
rect 15485 2465 15519 2499
rect 16037 2465 16071 2499
rect 16589 2465 16623 2499
rect 17509 2465 17543 2499
rect 11345 2397 11379 2431
rect 12081 2397 12115 2431
rect 13185 2397 13219 2431
rect 14197 2397 14231 2431
rect 10793 2329 10827 2363
rect 13645 2329 13679 2363
rect 16773 2329 16807 2363
rect 3801 2261 3835 2295
rect 5089 2261 5123 2295
rect 9781 2261 9815 2295
rect 10609 2261 10643 2295
rect 12633 2261 12667 2295
rect 16221 2261 16255 2295
rect 17693 2261 17727 2295
<< metal1 >>
rect 4062 21088 4068 21140
rect 4120 21128 4126 21140
rect 6270 21128 6276 21140
rect 4120 21100 6276 21128
rect 4120 21088 4126 21100
rect 6270 21088 6276 21100
rect 6328 21088 6334 21140
rect 3970 20952 3976 21004
rect 4028 20992 4034 21004
rect 8202 20992 8208 21004
rect 4028 20964 8208 20992
rect 4028 20952 4034 20964
rect 8202 20952 8208 20964
rect 8260 20952 8266 21004
rect 3510 20816 3516 20868
rect 3568 20856 3574 20868
rect 7374 20856 7380 20868
rect 3568 20828 7380 20856
rect 3568 20816 3574 20828
rect 7374 20816 7380 20828
rect 7432 20816 7438 20868
rect 8662 20816 8668 20868
rect 8720 20856 8726 20868
rect 9030 20856 9036 20868
rect 8720 20828 9036 20856
rect 8720 20816 8726 20828
rect 9030 20816 9036 20828
rect 9088 20816 9094 20868
rect 3326 20680 3332 20732
rect 3384 20720 3390 20732
rect 6454 20720 6460 20732
rect 3384 20692 6460 20720
rect 3384 20680 3390 20692
rect 6454 20680 6460 20692
rect 6512 20680 6518 20732
rect 3326 20408 3332 20460
rect 3384 20448 3390 20460
rect 4982 20448 4988 20460
rect 3384 20420 4988 20448
rect 3384 20408 3390 20420
rect 4982 20408 4988 20420
rect 5040 20408 5046 20460
rect 5718 20408 5724 20460
rect 5776 20448 5782 20460
rect 6822 20448 6828 20460
rect 5776 20420 6828 20448
rect 5776 20408 5782 20420
rect 6822 20408 6828 20420
rect 6880 20408 6886 20460
rect 2222 20340 2228 20392
rect 2280 20380 2286 20392
rect 6914 20380 6920 20392
rect 2280 20352 6920 20380
rect 2280 20340 2286 20352
rect 6914 20340 6920 20352
rect 6972 20340 6978 20392
rect 2866 20272 2872 20324
rect 2924 20312 2930 20324
rect 9766 20312 9772 20324
rect 2924 20284 9772 20312
rect 2924 20272 2930 20284
rect 9766 20272 9772 20284
rect 9824 20272 9830 20324
rect 4062 20204 4068 20256
rect 4120 20244 4126 20256
rect 8846 20244 8852 20256
rect 4120 20216 8852 20244
rect 4120 20204 4126 20216
rect 8846 20204 8852 20216
rect 8904 20204 8910 20256
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 3421 20043 3479 20049
rect 3421 20009 3433 20043
rect 3467 20040 3479 20043
rect 5166 20040 5172 20052
rect 3467 20012 5172 20040
rect 3467 20009 3479 20012
rect 3421 20003 3479 20009
rect 5166 20000 5172 20012
rect 5224 20000 5230 20052
rect 5258 20000 5264 20052
rect 5316 20040 5322 20052
rect 5813 20043 5871 20049
rect 5813 20040 5825 20043
rect 5316 20012 5825 20040
rect 5316 20000 5322 20012
rect 5813 20009 5825 20012
rect 5859 20009 5871 20043
rect 5813 20003 5871 20009
rect 8938 20000 8944 20052
rect 8996 20040 9002 20052
rect 12805 20043 12863 20049
rect 8996 20012 11928 20040
rect 8996 20000 9002 20012
rect 2501 19975 2559 19981
rect 2501 19941 2513 19975
rect 2547 19972 2559 19975
rect 2866 19972 2872 19984
rect 2547 19944 2872 19972
rect 2547 19941 2559 19944
rect 2501 19935 2559 19941
rect 2866 19932 2872 19944
rect 2924 19932 2930 19984
rect 3329 19975 3387 19981
rect 3329 19941 3341 19975
rect 3375 19972 3387 19975
rect 6365 19975 6423 19981
rect 6365 19972 6377 19975
rect 3375 19944 6377 19972
rect 3375 19941 3387 19944
rect 3329 19935 3387 19941
rect 6365 19941 6377 19944
rect 6411 19941 6423 19975
rect 6365 19935 6423 19941
rect 9033 19975 9091 19981
rect 9033 19941 9045 19975
rect 9079 19972 9091 19975
rect 11790 19972 11796 19984
rect 9079 19944 11796 19972
rect 9079 19941 9091 19944
rect 9033 19935 9091 19941
rect 11790 19932 11796 19944
rect 11848 19932 11854 19984
rect 1670 19904 1676 19916
rect 1631 19876 1676 19904
rect 1670 19864 1676 19876
rect 1728 19864 1734 19916
rect 2222 19904 2228 19916
rect 2183 19876 2228 19904
rect 2222 19864 2228 19876
rect 2280 19864 2286 19916
rect 3602 19864 3608 19916
rect 3660 19904 3666 19916
rect 4617 19907 4675 19913
rect 4617 19904 4629 19907
rect 3660 19876 4629 19904
rect 3660 19864 3666 19876
rect 4617 19873 4629 19876
rect 4663 19873 4675 19907
rect 4617 19867 4675 19873
rect 5626 19864 5632 19916
rect 5684 19904 5690 19916
rect 5721 19907 5779 19913
rect 5721 19904 5733 19907
rect 5684 19876 5733 19904
rect 5684 19864 5690 19876
rect 5721 19873 5733 19876
rect 5767 19873 5779 19907
rect 7006 19904 7012 19916
rect 5721 19867 5779 19873
rect 6840 19876 7012 19904
rect 3513 19839 3571 19845
rect 3513 19805 3525 19839
rect 3559 19836 3571 19839
rect 4706 19836 4712 19848
rect 3559 19808 4568 19836
rect 4667 19808 4712 19836
rect 3559 19805 3571 19808
rect 3513 19799 3571 19805
rect 1854 19700 1860 19712
rect 1815 19672 1860 19700
rect 1854 19660 1860 19672
rect 1912 19660 1918 19712
rect 2958 19700 2964 19712
rect 2919 19672 2964 19700
rect 2958 19660 2964 19672
rect 3016 19660 3022 19712
rect 4154 19660 4160 19712
rect 4212 19700 4218 19712
rect 4249 19703 4307 19709
rect 4249 19700 4261 19703
rect 4212 19672 4261 19700
rect 4212 19660 4218 19672
rect 4249 19669 4261 19672
rect 4295 19669 4307 19703
rect 4540 19700 4568 19808
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 4890 19836 4896 19848
rect 4851 19808 4896 19836
rect 4890 19796 4896 19808
rect 4948 19796 4954 19848
rect 5994 19836 6000 19848
rect 5955 19808 6000 19836
rect 5994 19796 6000 19808
rect 6052 19796 6058 19848
rect 5166 19728 5172 19780
rect 5224 19768 5230 19780
rect 5353 19771 5411 19777
rect 5353 19768 5365 19771
rect 5224 19740 5365 19768
rect 5224 19728 5230 19740
rect 5353 19737 5365 19740
rect 5399 19737 5411 19771
rect 5353 19731 5411 19737
rect 6840 19700 6868 19876
rect 7006 19864 7012 19876
rect 7064 19904 7070 19916
rect 7173 19907 7231 19913
rect 7173 19904 7185 19907
rect 7064 19876 7185 19904
rect 7064 19864 7070 19876
rect 7173 19873 7185 19876
rect 7219 19873 7231 19907
rect 7173 19867 7231 19873
rect 9125 19907 9183 19913
rect 9125 19873 9137 19907
rect 9171 19904 9183 19907
rect 9674 19904 9680 19916
rect 9171 19876 9680 19904
rect 9171 19873 9183 19876
rect 9125 19867 9183 19873
rect 9674 19864 9680 19876
rect 9732 19864 9738 19916
rect 9769 19907 9827 19913
rect 9769 19873 9781 19907
rect 9815 19873 9827 19907
rect 10502 19904 10508 19916
rect 10463 19876 10508 19904
rect 9769 19867 9827 19873
rect 6917 19839 6975 19845
rect 6917 19805 6929 19839
rect 6963 19805 6975 19839
rect 9214 19836 9220 19848
rect 9175 19808 9220 19836
rect 6917 19799 6975 19805
rect 4540 19672 6868 19700
rect 6932 19700 6960 19799
rect 9214 19796 9220 19808
rect 9272 19796 9278 19848
rect 8665 19771 8723 19777
rect 8665 19737 8677 19771
rect 8711 19768 8723 19771
rect 9784 19768 9812 19867
rect 10502 19864 10508 19876
rect 10560 19864 10566 19916
rect 11900 19913 11928 20012
rect 12805 20009 12817 20043
rect 12851 20040 12863 20043
rect 13170 20040 13176 20052
rect 12851 20012 13176 20040
rect 12851 20009 12863 20012
rect 12805 20003 12863 20009
rect 13170 20000 13176 20012
rect 13228 20000 13234 20052
rect 13357 20043 13415 20049
rect 13357 20009 13369 20043
rect 13403 20040 13415 20043
rect 13630 20040 13636 20052
rect 13403 20012 13636 20040
rect 13403 20009 13415 20012
rect 13357 20003 13415 20009
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 16669 20043 16727 20049
rect 16669 20009 16681 20043
rect 16715 20040 16727 20043
rect 17402 20040 17408 20052
rect 16715 20012 17408 20040
rect 16715 20009 16727 20012
rect 16669 20003 16727 20009
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 12158 19932 12164 19984
rect 12216 19972 12222 19984
rect 12216 19944 13768 19972
rect 12216 19932 12222 19944
rect 11333 19907 11391 19913
rect 11333 19873 11345 19907
rect 11379 19873 11391 19907
rect 11333 19867 11391 19873
rect 11885 19907 11943 19913
rect 11885 19873 11897 19907
rect 11931 19873 11943 19907
rect 12342 19904 12348 19916
rect 11885 19867 11943 19873
rect 11992 19876 12348 19904
rect 9953 19839 10011 19845
rect 9953 19805 9965 19839
rect 9999 19805 10011 19839
rect 9953 19799 10011 19805
rect 8711 19740 9812 19768
rect 8711 19737 8723 19740
rect 8665 19731 8723 19737
rect 7282 19700 7288 19712
rect 6932 19672 7288 19700
rect 4249 19663 4307 19669
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 7650 19660 7656 19712
rect 7708 19700 7714 19712
rect 8297 19703 8355 19709
rect 8297 19700 8309 19703
rect 7708 19672 8309 19700
rect 7708 19660 7714 19672
rect 8297 19669 8309 19672
rect 8343 19669 8355 19703
rect 8297 19663 8355 19669
rect 8386 19660 8392 19712
rect 8444 19700 8450 19712
rect 9968 19700 9996 19799
rect 10042 19796 10048 19848
rect 10100 19836 10106 19848
rect 10689 19839 10747 19845
rect 10689 19836 10701 19839
rect 10100 19808 10701 19836
rect 10100 19796 10106 19808
rect 10689 19805 10701 19808
rect 10735 19805 10747 19839
rect 11348 19836 11376 19867
rect 11992 19836 12020 19876
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 12618 19904 12624 19916
rect 12579 19876 12624 19904
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 13173 19907 13231 19913
rect 13173 19873 13185 19907
rect 13219 19904 13231 19907
rect 13354 19904 13360 19916
rect 13219 19876 13360 19904
rect 13219 19873 13231 19876
rect 13173 19867 13231 19873
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 13740 19913 13768 19944
rect 19334 19932 19340 19984
rect 19392 19972 19398 19984
rect 20162 19972 20168 19984
rect 19392 19944 20168 19972
rect 19392 19932 19398 19944
rect 20162 19932 20168 19944
rect 20220 19932 20226 19984
rect 13725 19907 13783 19913
rect 13725 19873 13737 19907
rect 13771 19873 13783 19907
rect 13725 19867 13783 19873
rect 16390 19864 16396 19916
rect 16448 19904 16454 19916
rect 16485 19907 16543 19913
rect 16485 19904 16497 19907
rect 16448 19876 16497 19904
rect 16448 19864 16454 19876
rect 16485 19873 16497 19876
rect 16531 19873 16543 19907
rect 16485 19867 16543 19873
rect 19702 19836 19708 19848
rect 11348 19808 12020 19836
rect 12084 19808 19708 19836
rect 10689 19799 10747 19805
rect 12084 19777 12112 19808
rect 19702 19796 19708 19808
rect 19760 19796 19766 19848
rect 12069 19771 12127 19777
rect 12069 19737 12081 19771
rect 12115 19737 12127 19771
rect 12069 19731 12127 19737
rect 12268 19740 19380 19768
rect 8444 19672 9996 19700
rect 11517 19703 11575 19709
rect 8444 19660 8450 19672
rect 11517 19669 11529 19703
rect 11563 19700 11575 19703
rect 12268 19700 12296 19740
rect 19352 19712 19380 19740
rect 11563 19672 12296 19700
rect 13909 19703 13967 19709
rect 11563 19669 11575 19672
rect 11517 19663 11575 19669
rect 13909 19669 13921 19703
rect 13955 19700 13967 19703
rect 18690 19700 18696 19712
rect 13955 19672 18696 19700
rect 13955 19669 13967 19672
rect 13909 19663 13967 19669
rect 18690 19660 18696 19672
rect 18748 19660 18754 19712
rect 19334 19660 19340 19712
rect 19392 19660 19398 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 4062 19456 4068 19508
rect 4120 19496 4126 19508
rect 5718 19496 5724 19508
rect 4120 19468 5724 19496
rect 4120 19456 4126 19468
rect 5718 19456 5724 19468
rect 5776 19456 5782 19508
rect 6914 19496 6920 19508
rect 6875 19468 6920 19496
rect 6914 19456 6920 19468
rect 6972 19456 6978 19508
rect 8404 19468 9444 19496
rect 3528 19400 4200 19428
rect 3528 19369 3556 19400
rect 3513 19363 3571 19369
rect 3513 19329 3525 19363
rect 3559 19329 3571 19363
rect 4172 19360 4200 19400
rect 5626 19388 5632 19440
rect 5684 19428 5690 19440
rect 6730 19428 6736 19440
rect 5684 19400 6736 19428
rect 5684 19388 5690 19400
rect 6730 19388 6736 19400
rect 6788 19388 6794 19440
rect 7742 19388 7748 19440
rect 7800 19428 7806 19440
rect 8404 19428 8432 19468
rect 7800 19400 8432 19428
rect 7800 19388 7806 19400
rect 7561 19363 7619 19369
rect 4172 19332 4292 19360
rect 3513 19323 3571 19329
rect 4264 19304 4292 19332
rect 7561 19329 7573 19363
rect 7607 19360 7619 19363
rect 8294 19360 8300 19372
rect 7607 19332 8300 19360
rect 7607 19329 7619 19332
rect 7561 19323 7619 19329
rect 8294 19320 8300 19332
rect 8352 19320 8358 19372
rect 1578 19292 1584 19304
rect 1539 19264 1584 19292
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 2133 19295 2191 19301
rect 2133 19261 2145 19295
rect 2179 19292 2191 19295
rect 3970 19292 3976 19304
rect 2179 19264 3976 19292
rect 2179 19261 2191 19264
rect 2133 19255 2191 19261
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 4157 19295 4215 19301
rect 4157 19292 4169 19295
rect 4080 19264 4169 19292
rect 2406 19224 2412 19236
rect 2367 19196 2412 19224
rect 2406 19184 2412 19196
rect 2464 19184 2470 19236
rect 3050 19184 3056 19236
rect 3108 19224 3114 19236
rect 3237 19227 3295 19233
rect 3237 19224 3249 19227
rect 3108 19196 3249 19224
rect 3108 19184 3114 19196
rect 3237 19193 3249 19196
rect 3283 19193 3295 19227
rect 3237 19187 3295 19193
rect 4080 19168 4108 19264
rect 4157 19261 4169 19264
rect 4203 19261 4215 19295
rect 4157 19255 4215 19261
rect 4246 19252 4252 19304
rect 4304 19252 4310 19304
rect 5810 19292 5816 19304
rect 4356 19264 5580 19292
rect 5771 19264 5816 19292
rect 1762 19156 1768 19168
rect 1723 19128 1768 19156
rect 1762 19116 1768 19128
rect 1820 19116 1826 19168
rect 2130 19116 2136 19168
rect 2188 19156 2194 19168
rect 2869 19159 2927 19165
rect 2869 19156 2881 19159
rect 2188 19128 2881 19156
rect 2188 19116 2194 19128
rect 2869 19125 2881 19128
rect 2915 19125 2927 19159
rect 3326 19156 3332 19168
rect 3287 19128 3332 19156
rect 2869 19119 2927 19125
rect 3326 19116 3332 19128
rect 3384 19116 3390 19168
rect 4062 19116 4068 19168
rect 4120 19116 4126 19168
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 4356 19156 4384 19264
rect 4424 19227 4482 19233
rect 4424 19193 4436 19227
rect 4470 19224 4482 19227
rect 5442 19224 5448 19236
rect 4470 19196 5448 19224
rect 4470 19193 4482 19196
rect 4424 19187 4482 19193
rect 5442 19184 5448 19196
rect 5500 19184 5506 19236
rect 5552 19224 5580 19264
rect 5810 19252 5816 19264
rect 5868 19252 5874 19304
rect 6914 19252 6920 19304
rect 6972 19292 6978 19304
rect 7377 19295 7435 19301
rect 7377 19292 7389 19295
rect 6972 19264 7389 19292
rect 6972 19252 6978 19264
rect 7377 19261 7389 19264
rect 7423 19261 7435 19295
rect 7377 19255 7435 19261
rect 7466 19252 7472 19304
rect 7524 19292 7530 19304
rect 8404 19301 8432 19400
rect 9416 19360 9444 19468
rect 10045 19363 10103 19369
rect 10045 19360 10057 19363
rect 9416 19332 10057 19360
rect 10045 19329 10057 19332
rect 10091 19329 10103 19363
rect 10045 19323 10103 19329
rect 8389 19295 8447 19301
rect 7524 19264 8340 19292
rect 7524 19252 7530 19264
rect 7285 19227 7343 19233
rect 5552 19196 6040 19224
rect 4212 19128 4384 19156
rect 4212 19116 4218 19128
rect 4890 19116 4896 19168
rect 4948 19156 4954 19168
rect 6012 19165 6040 19196
rect 7285 19193 7297 19227
rect 7331 19224 7343 19227
rect 7929 19227 7987 19233
rect 7929 19224 7941 19227
rect 7331 19196 7941 19224
rect 7331 19193 7343 19196
rect 7285 19187 7343 19193
rect 7929 19193 7941 19196
rect 7975 19193 7987 19227
rect 8312 19224 8340 19264
rect 8389 19261 8401 19295
rect 8435 19261 8447 19295
rect 11054 19292 11060 19304
rect 8389 19255 8447 19261
rect 8588 19264 11060 19292
rect 8588 19224 8616 19264
rect 11054 19252 11060 19264
rect 11112 19252 11118 19304
rect 11698 19292 11704 19304
rect 11659 19264 11704 19292
rect 11698 19252 11704 19264
rect 11756 19252 11762 19304
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 12526 19292 12532 19304
rect 12483 19264 12532 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 14093 19295 14151 19301
rect 14093 19261 14105 19295
rect 14139 19292 14151 19295
rect 14182 19292 14188 19304
rect 14139 19264 14188 19292
rect 14139 19261 14151 19264
rect 14093 19255 14151 19261
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 14645 19295 14703 19301
rect 14645 19292 14657 19295
rect 14332 19264 14657 19292
rect 14332 19252 14338 19264
rect 14645 19261 14657 19264
rect 14691 19261 14703 19295
rect 15194 19292 15200 19304
rect 15155 19264 15200 19292
rect 14645 19255 14703 19261
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 15746 19292 15752 19304
rect 15707 19264 15752 19292
rect 15746 19252 15752 19264
rect 15804 19252 15810 19304
rect 16298 19292 16304 19304
rect 16259 19264 16304 19292
rect 16298 19252 16304 19264
rect 16356 19252 16362 19304
rect 16850 19292 16856 19304
rect 16811 19264 16856 19292
rect 16850 19252 16856 19264
rect 16908 19252 16914 19304
rect 17405 19295 17463 19301
rect 17405 19292 17417 19295
rect 16960 19264 17417 19292
rect 8312 19196 8616 19224
rect 8656 19227 8714 19233
rect 7929 19187 7987 19193
rect 8656 19193 8668 19227
rect 8702 19224 8714 19227
rect 10134 19224 10140 19236
rect 8702 19196 10140 19224
rect 8702 19193 8714 19196
rect 8656 19187 8714 19193
rect 10134 19184 10140 19196
rect 10192 19184 10198 19236
rect 10226 19184 10232 19236
rect 10284 19233 10290 19236
rect 12710 19233 12716 19236
rect 10284 19227 10348 19233
rect 10284 19193 10302 19227
rect 10336 19193 10348 19227
rect 12704 19224 12716 19233
rect 12671 19196 12716 19224
rect 10284 19187 10348 19193
rect 12704 19187 12716 19196
rect 10284 19184 10290 19187
rect 12710 19184 12716 19187
rect 12768 19184 12774 19236
rect 13630 19184 13636 19236
rect 13688 19224 13694 19236
rect 16960 19224 16988 19264
rect 17405 19261 17417 19264
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 17494 19252 17500 19304
rect 17552 19292 17558 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17552 19264 18061 19292
rect 17552 19252 17558 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 18601 19295 18659 19301
rect 18601 19261 18613 19295
rect 18647 19261 18659 19295
rect 19150 19292 19156 19304
rect 19111 19264 19156 19292
rect 18601 19255 18659 19261
rect 13688 19196 16988 19224
rect 13688 19184 13694 19196
rect 17310 19184 17316 19236
rect 17368 19224 17374 19236
rect 18616 19224 18644 19255
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 19702 19292 19708 19304
rect 19663 19264 19708 19292
rect 19702 19252 19708 19264
rect 19760 19252 19766 19304
rect 17368 19196 18644 19224
rect 17368 19184 17374 19196
rect 18690 19184 18696 19236
rect 18748 19224 18754 19236
rect 21542 19224 21548 19236
rect 18748 19196 21548 19224
rect 18748 19184 18754 19196
rect 21542 19184 21548 19196
rect 21600 19184 21606 19236
rect 5537 19159 5595 19165
rect 5537 19156 5549 19159
rect 4948 19128 5549 19156
rect 4948 19116 4954 19128
rect 5537 19125 5549 19128
rect 5583 19125 5595 19159
rect 5537 19119 5595 19125
rect 5997 19159 6055 19165
rect 5997 19125 6009 19159
rect 6043 19125 6055 19159
rect 5997 19119 6055 19125
rect 6270 19116 6276 19168
rect 6328 19156 6334 19168
rect 8478 19156 8484 19168
rect 6328 19128 8484 19156
rect 6328 19116 6334 19128
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 8570 19116 8576 19168
rect 8628 19156 8634 19168
rect 8754 19156 8760 19168
rect 8628 19128 8760 19156
rect 8628 19116 8634 19128
rect 8754 19116 8760 19128
rect 8812 19116 8818 19168
rect 9214 19116 9220 19168
rect 9272 19156 9278 19168
rect 9769 19159 9827 19165
rect 9769 19156 9781 19159
rect 9272 19128 9781 19156
rect 9272 19116 9278 19128
rect 9769 19125 9781 19128
rect 9815 19125 9827 19159
rect 10152 19156 10180 19184
rect 11425 19159 11483 19165
rect 11425 19156 11437 19159
rect 10152 19128 11437 19156
rect 9769 19119 9827 19125
rect 11425 19125 11437 19128
rect 11471 19125 11483 19159
rect 11425 19119 11483 19125
rect 11885 19159 11943 19165
rect 11885 19125 11897 19159
rect 11931 19156 11943 19159
rect 12066 19156 12072 19168
rect 11931 19128 12072 19156
rect 11931 19125 11943 19128
rect 11885 19119 11943 19125
rect 12066 19116 12072 19128
rect 12124 19116 12130 19168
rect 13814 19116 13820 19168
rect 13872 19156 13878 19168
rect 14277 19159 14335 19165
rect 13872 19128 13917 19156
rect 13872 19116 13878 19128
rect 14277 19125 14289 19159
rect 14323 19156 14335 19159
rect 14550 19156 14556 19168
rect 14323 19128 14556 19156
rect 14323 19125 14335 19128
rect 14277 19119 14335 19125
rect 14550 19116 14556 19128
rect 14608 19116 14614 19168
rect 14829 19159 14887 19165
rect 14829 19125 14841 19159
rect 14875 19156 14887 19159
rect 15010 19156 15016 19168
rect 14875 19128 15016 19156
rect 14875 19125 14887 19128
rect 14829 19119 14887 19125
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 15381 19159 15439 19165
rect 15381 19125 15393 19159
rect 15427 19156 15439 19159
rect 15562 19156 15568 19168
rect 15427 19128 15568 19156
rect 15427 19125 15439 19128
rect 15381 19119 15439 19125
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 15933 19159 15991 19165
rect 15933 19125 15945 19159
rect 15979 19156 15991 19159
rect 16022 19156 16028 19168
rect 15979 19128 16028 19156
rect 15979 19125 15991 19128
rect 15933 19119 15991 19125
rect 16022 19116 16028 19128
rect 16080 19116 16086 19168
rect 16482 19156 16488 19168
rect 16443 19128 16488 19156
rect 16482 19116 16488 19128
rect 16540 19116 16546 19168
rect 16942 19116 16948 19168
rect 17000 19156 17006 19168
rect 17037 19159 17095 19165
rect 17037 19156 17049 19159
rect 17000 19128 17049 19156
rect 17000 19116 17006 19128
rect 17037 19125 17049 19128
rect 17083 19125 17095 19159
rect 17037 19119 17095 19125
rect 17589 19159 17647 19165
rect 17589 19125 17601 19159
rect 17635 19156 17647 19159
rect 17862 19156 17868 19168
rect 17635 19128 17868 19156
rect 17635 19125 17647 19128
rect 17589 19119 17647 19125
rect 17862 19116 17868 19128
rect 17920 19116 17926 19168
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18506 19156 18512 19168
rect 18279 19128 18512 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18506 19116 18512 19128
rect 18564 19116 18570 19168
rect 18782 19156 18788 19168
rect 18743 19128 18788 19156
rect 18782 19116 18788 19128
rect 18840 19116 18846 19168
rect 19242 19116 19248 19168
rect 19300 19156 19306 19168
rect 19337 19159 19395 19165
rect 19337 19156 19349 19159
rect 19300 19128 19349 19156
rect 19300 19116 19306 19128
rect 19337 19125 19349 19128
rect 19383 19125 19395 19159
rect 19337 19119 19395 19125
rect 19889 19159 19947 19165
rect 19889 19125 19901 19159
rect 19935 19156 19947 19159
rect 20622 19156 20628 19168
rect 19935 19128 20628 19156
rect 19935 19125 19947 19128
rect 19889 19119 19947 19125
rect 20622 19116 20628 19128
rect 20680 19116 20686 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 2961 18955 3019 18961
rect 2961 18921 2973 18955
rect 3007 18952 3019 18955
rect 3326 18952 3332 18964
rect 3007 18924 3332 18952
rect 3007 18921 3019 18924
rect 2961 18915 3019 18921
rect 3326 18912 3332 18924
rect 3384 18912 3390 18964
rect 3421 18955 3479 18961
rect 3421 18921 3433 18955
rect 3467 18952 3479 18955
rect 3467 18924 6132 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 3252 18856 3464 18884
rect 1489 18819 1547 18825
rect 1489 18785 1501 18819
rect 1535 18816 1547 18819
rect 2130 18816 2136 18828
rect 1535 18788 2136 18816
rect 1535 18785 1547 18788
rect 1489 18779 1547 18785
rect 2130 18776 2136 18788
rect 2188 18776 2194 18828
rect 2225 18819 2283 18825
rect 2225 18785 2237 18819
rect 2271 18816 2283 18819
rect 2958 18816 2964 18828
rect 2271 18788 2964 18816
rect 2271 18785 2283 18788
rect 2225 18779 2283 18785
rect 2958 18776 2964 18788
rect 3016 18776 3022 18828
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18717 1823 18751
rect 2498 18748 2504 18760
rect 2459 18720 2504 18748
rect 1765 18711 1823 18717
rect 1780 18612 1808 18711
rect 2498 18708 2504 18720
rect 2556 18708 2562 18760
rect 3252 18612 3280 18856
rect 3329 18819 3387 18825
rect 3329 18785 3341 18819
rect 3375 18785 3387 18819
rect 3436 18816 3464 18856
rect 4246 18844 4252 18896
rect 4304 18893 4310 18896
rect 4304 18887 4368 18893
rect 4304 18853 4322 18887
rect 4356 18853 4368 18887
rect 4304 18847 4368 18853
rect 4304 18844 4310 18847
rect 4430 18844 4436 18896
rect 4488 18884 4494 18896
rect 5810 18884 5816 18896
rect 4488 18856 5816 18884
rect 4488 18844 4494 18856
rect 5810 18844 5816 18856
rect 5868 18844 5874 18896
rect 5994 18893 6000 18896
rect 5988 18884 6000 18893
rect 5955 18856 6000 18884
rect 5988 18847 6000 18856
rect 5994 18844 6000 18847
rect 6052 18844 6058 18896
rect 6104 18884 6132 18924
rect 7006 18912 7012 18964
rect 7064 18952 7070 18964
rect 7101 18955 7159 18961
rect 7101 18952 7113 18955
rect 7064 18924 7113 18952
rect 7064 18912 7070 18924
rect 7101 18921 7113 18924
rect 7147 18921 7159 18955
rect 7101 18915 7159 18921
rect 7208 18924 7779 18952
rect 7208 18884 7236 18924
rect 7650 18893 7656 18896
rect 6104 18856 7236 18884
rect 7285 18887 7343 18893
rect 7285 18853 7297 18887
rect 7331 18884 7343 18887
rect 7622 18887 7656 18893
rect 7622 18884 7634 18887
rect 7331 18856 7634 18884
rect 7331 18853 7343 18856
rect 7285 18847 7343 18853
rect 7622 18853 7634 18856
rect 7622 18847 7656 18853
rect 7650 18844 7656 18847
rect 7708 18844 7714 18896
rect 7751 18884 7779 18924
rect 8294 18912 8300 18964
rect 8352 18952 8358 18964
rect 8757 18955 8815 18961
rect 8757 18952 8769 18955
rect 8352 18924 8769 18952
rect 8352 18912 8358 18924
rect 8757 18921 8769 18924
rect 8803 18921 8815 18955
rect 8757 18915 8815 18921
rect 8662 18884 8668 18896
rect 7751 18856 8668 18884
rect 8662 18844 8668 18856
rect 8720 18844 8726 18896
rect 8763 18884 8791 18915
rect 8846 18912 8852 18964
rect 8904 18952 8910 18964
rect 9217 18955 9275 18961
rect 9217 18952 9229 18955
rect 8904 18924 9229 18952
rect 8904 18912 8910 18924
rect 9217 18921 9229 18924
rect 9263 18921 9275 18955
rect 9217 18915 9275 18921
rect 9674 18912 9680 18964
rect 9732 18952 9738 18964
rect 9861 18955 9919 18961
rect 9861 18952 9873 18955
rect 9732 18924 9873 18952
rect 9732 18912 9738 18924
rect 9861 18921 9873 18924
rect 9907 18921 9919 18955
rect 9861 18915 9919 18921
rect 10321 18955 10379 18961
rect 10321 18921 10333 18955
rect 10367 18952 10379 18955
rect 10870 18952 10876 18964
rect 10367 18924 10876 18952
rect 10367 18921 10379 18924
rect 10321 18915 10379 18921
rect 10870 18912 10876 18924
rect 10928 18912 10934 18964
rect 11054 18912 11060 18964
rect 11112 18952 11118 18964
rect 11112 18924 12756 18952
rect 11112 18912 11118 18924
rect 12728 18884 12756 18924
rect 12802 18912 12808 18964
rect 12860 18952 12866 18964
rect 13265 18955 13323 18961
rect 13265 18952 13277 18955
rect 12860 18924 13277 18952
rect 12860 18912 12866 18924
rect 13265 18921 13277 18924
rect 13311 18921 13323 18955
rect 13265 18915 13323 18921
rect 12986 18884 12992 18896
rect 8763 18856 8984 18884
rect 12728 18856 12992 18884
rect 8754 18816 8760 18828
rect 3436 18788 8760 18816
rect 3329 18779 3387 18785
rect 3344 18748 3372 18779
rect 8754 18776 8760 18788
rect 8812 18776 8818 18828
rect 3418 18748 3424 18760
rect 3344 18720 3424 18748
rect 3418 18708 3424 18720
rect 3476 18708 3482 18760
rect 3510 18708 3516 18760
rect 3568 18748 3574 18760
rect 3605 18751 3663 18757
rect 3605 18748 3617 18751
rect 3568 18720 3617 18748
rect 3568 18708 3574 18720
rect 3605 18717 3617 18720
rect 3651 18748 3663 18751
rect 4062 18748 4068 18760
rect 3651 18720 3924 18748
rect 4023 18720 4068 18748
rect 3651 18717 3663 18720
rect 3605 18711 3663 18717
rect 1780 18584 3280 18612
rect 3896 18612 3924 18720
rect 4062 18708 4068 18720
rect 4120 18708 4126 18760
rect 5350 18708 5356 18760
rect 5408 18748 5414 18760
rect 5721 18751 5779 18757
rect 5721 18748 5733 18751
rect 5408 18720 5733 18748
rect 5408 18708 5414 18720
rect 5721 18717 5733 18720
rect 5767 18717 5779 18751
rect 5721 18711 5779 18717
rect 7282 18708 7288 18760
rect 7340 18748 7346 18760
rect 7377 18751 7435 18757
rect 7377 18748 7389 18751
rect 7340 18720 7389 18748
rect 7340 18708 7346 18720
rect 7377 18717 7389 18720
rect 7423 18717 7435 18751
rect 8956 18748 8984 18856
rect 12986 18844 12992 18856
rect 13044 18844 13050 18896
rect 14093 18887 14151 18893
rect 14093 18853 14105 18887
rect 14139 18884 14151 18887
rect 14274 18884 14280 18896
rect 14139 18856 14280 18884
rect 14139 18853 14151 18856
rect 14093 18847 14151 18853
rect 14274 18844 14280 18856
rect 14332 18844 14338 18896
rect 15565 18887 15623 18893
rect 15565 18853 15577 18887
rect 15611 18884 15623 18887
rect 16850 18884 16856 18896
rect 15611 18856 16856 18884
rect 15611 18853 15623 18856
rect 15565 18847 15623 18853
rect 16850 18844 16856 18856
rect 16908 18844 16914 18896
rect 19061 18887 19119 18893
rect 19061 18853 19073 18887
rect 19107 18884 19119 18887
rect 19702 18884 19708 18896
rect 19107 18856 19708 18884
rect 19107 18853 19119 18856
rect 19061 18847 19119 18853
rect 19702 18844 19708 18856
rect 19760 18844 19766 18896
rect 9033 18819 9091 18825
rect 9033 18785 9045 18819
rect 9079 18816 9091 18819
rect 10042 18816 10048 18828
rect 9079 18788 10048 18816
rect 9079 18785 9091 18788
rect 9033 18779 9091 18785
rect 10042 18776 10048 18788
rect 10100 18776 10106 18828
rect 10229 18819 10287 18825
rect 10229 18785 10241 18819
rect 10275 18816 10287 18819
rect 10686 18816 10692 18828
rect 10275 18788 10692 18816
rect 10275 18785 10287 18788
rect 10229 18779 10287 18785
rect 10686 18776 10692 18788
rect 10744 18776 10750 18828
rect 11416 18819 11474 18825
rect 11416 18785 11428 18819
rect 11462 18816 11474 18819
rect 11974 18816 11980 18828
rect 11462 18788 11980 18816
rect 11462 18785 11474 18788
rect 11416 18779 11474 18785
rect 11974 18776 11980 18788
rect 12032 18776 12038 18828
rect 13173 18819 13231 18825
rect 13173 18785 13185 18819
rect 13219 18816 13231 18819
rect 13262 18816 13268 18828
rect 13219 18788 13268 18816
rect 13219 18785 13231 18788
rect 13173 18779 13231 18785
rect 13262 18776 13268 18788
rect 13320 18776 13326 18828
rect 13814 18816 13820 18828
rect 13775 18788 13820 18816
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 15289 18819 15347 18825
rect 15289 18785 15301 18819
rect 15335 18816 15347 18819
rect 15378 18816 15384 18828
rect 15335 18788 15384 18816
rect 15335 18785 15347 18788
rect 15289 18779 15347 18785
rect 15378 18776 15384 18788
rect 15436 18776 15442 18828
rect 18782 18816 18788 18828
rect 18743 18788 18788 18816
rect 18782 18776 18788 18788
rect 18840 18776 18846 18828
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 21082 18816 21088 18828
rect 19392 18788 21088 18816
rect 19392 18776 19398 18788
rect 21082 18776 21088 18788
rect 21140 18776 21146 18828
rect 9858 18748 9864 18760
rect 8956 18720 9864 18748
rect 7377 18711 7435 18717
rect 9858 18708 9864 18720
rect 9916 18708 9922 18760
rect 10134 18708 10140 18760
rect 10192 18748 10198 18760
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 10192 18720 10425 18748
rect 10192 18708 10198 18720
rect 10413 18717 10425 18720
rect 10459 18717 10471 18751
rect 10413 18711 10471 18717
rect 10594 18708 10600 18760
rect 10652 18748 10658 18760
rect 11149 18751 11207 18757
rect 11149 18748 11161 18751
rect 10652 18720 11161 18748
rect 10652 18708 10658 18720
rect 11149 18717 11161 18720
rect 11195 18717 11207 18751
rect 11149 18711 11207 18717
rect 13357 18751 13415 18757
rect 13357 18717 13369 18751
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 5442 18680 5448 18692
rect 5403 18652 5448 18680
rect 5442 18640 5448 18652
rect 5500 18640 5506 18692
rect 7006 18640 7012 18692
rect 7064 18680 7070 18692
rect 7193 18683 7251 18689
rect 7193 18680 7205 18683
rect 7064 18652 7205 18680
rect 7064 18640 7070 18652
rect 7193 18649 7205 18652
rect 7239 18649 7251 18683
rect 7193 18643 7251 18649
rect 8478 18640 8484 18692
rect 8536 18680 8542 18692
rect 10318 18680 10324 18692
rect 8536 18652 10324 18680
rect 8536 18640 8542 18652
rect 10318 18640 10324 18652
rect 10376 18640 10382 18692
rect 12529 18683 12587 18689
rect 12529 18649 12541 18683
rect 12575 18680 12587 18683
rect 12710 18680 12716 18692
rect 12575 18652 12716 18680
rect 12575 18649 12587 18652
rect 12529 18643 12587 18649
rect 12710 18640 12716 18652
rect 12768 18680 12774 18692
rect 13372 18680 13400 18711
rect 12768 18652 13400 18680
rect 12768 18640 12774 18652
rect 6362 18612 6368 18624
rect 3896 18584 6368 18612
rect 6362 18572 6368 18584
rect 6420 18572 6426 18624
rect 6454 18572 6460 18624
rect 6512 18612 6518 18624
rect 12066 18612 12072 18624
rect 6512 18584 12072 18612
rect 6512 18572 6518 18584
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 12802 18612 12808 18624
rect 12763 18584 12808 18612
rect 12802 18572 12808 18584
rect 12860 18572 12866 18624
rect 12986 18572 12992 18624
rect 13044 18612 13050 18624
rect 15102 18612 15108 18624
rect 13044 18584 15108 18612
rect 13044 18572 13050 18584
rect 15102 18572 15108 18584
rect 15160 18572 15166 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 3050 18408 3056 18420
rect 2332 18380 3056 18408
rect 2332 18281 2360 18380
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 4157 18411 4215 18417
rect 4157 18377 4169 18411
rect 4203 18408 4215 18411
rect 4246 18408 4252 18420
rect 4203 18380 4252 18408
rect 4203 18377 4215 18380
rect 4157 18371 4215 18377
rect 4246 18368 4252 18380
rect 4304 18368 4310 18420
rect 5994 18368 6000 18420
rect 6052 18408 6058 18420
rect 6089 18411 6147 18417
rect 6089 18408 6101 18411
rect 6052 18380 6101 18408
rect 6052 18368 6058 18380
rect 6089 18377 6101 18380
rect 6135 18377 6147 18411
rect 6089 18371 6147 18377
rect 6362 18368 6368 18420
rect 6420 18408 6426 18420
rect 9861 18411 9919 18417
rect 9861 18408 9873 18411
rect 6420 18380 9873 18408
rect 6420 18368 6426 18380
rect 9861 18377 9873 18380
rect 9907 18377 9919 18411
rect 10318 18408 10324 18420
rect 10279 18380 10324 18408
rect 9861 18371 9919 18377
rect 10318 18368 10324 18380
rect 10376 18368 10382 18420
rect 10502 18368 10508 18420
rect 10560 18408 10566 18420
rect 10781 18411 10839 18417
rect 10781 18408 10793 18411
rect 10560 18380 10793 18408
rect 10560 18368 10566 18380
rect 10781 18377 10793 18380
rect 10827 18377 10839 18411
rect 13722 18408 13728 18420
rect 10781 18371 10839 18377
rect 11164 18380 13728 18408
rect 5718 18300 5724 18352
rect 5776 18340 5782 18352
rect 7009 18343 7067 18349
rect 7009 18340 7021 18343
rect 5776 18312 7021 18340
rect 5776 18300 5782 18312
rect 7009 18309 7021 18312
rect 7055 18309 7067 18343
rect 7009 18303 7067 18309
rect 7190 18300 7196 18352
rect 7248 18340 7254 18352
rect 7742 18340 7748 18352
rect 7248 18312 7748 18340
rect 7248 18300 7254 18312
rect 7742 18300 7748 18312
rect 7800 18340 7806 18352
rect 7800 18312 8524 18340
rect 7800 18300 7806 18312
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18241 2375 18275
rect 2317 18235 2375 18241
rect 7834 18232 7840 18284
rect 7892 18232 7898 18284
rect 8110 18272 8116 18284
rect 8071 18244 8116 18272
rect 8110 18232 8116 18244
rect 8168 18232 8174 18284
rect 8496 18281 8524 18312
rect 9490 18300 9496 18352
rect 9548 18340 9554 18352
rect 11164 18340 11192 18380
rect 13722 18368 13728 18380
rect 13780 18368 13786 18420
rect 12802 18340 12808 18352
rect 9548 18312 11192 18340
rect 11256 18312 12808 18340
rect 9548 18300 9554 18312
rect 11256 18281 11284 18312
rect 12802 18300 12808 18312
rect 12860 18300 12866 18352
rect 8481 18275 8539 18281
rect 8481 18241 8493 18275
rect 8527 18241 8539 18275
rect 8481 18235 8539 18241
rect 11241 18275 11299 18281
rect 11241 18241 11253 18275
rect 11287 18241 11299 18275
rect 11241 18235 11299 18241
rect 11425 18275 11483 18281
rect 11425 18241 11437 18275
rect 11471 18272 11483 18275
rect 11606 18272 11612 18284
rect 11471 18244 11612 18272
rect 11471 18241 11483 18244
rect 11425 18235 11483 18241
rect 11606 18232 11612 18244
rect 11664 18232 11670 18284
rect 11790 18272 11796 18284
rect 11751 18244 11796 18272
rect 11790 18232 11796 18244
rect 11848 18232 11854 18284
rect 12618 18272 12624 18284
rect 12579 18244 12624 18272
rect 12618 18232 12624 18244
rect 12676 18232 12682 18284
rect 13354 18272 13360 18284
rect 13315 18244 13360 18272
rect 13354 18232 13360 18244
rect 13412 18232 13418 18284
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 2682 18164 2688 18216
rect 2740 18204 2746 18216
rect 2777 18207 2835 18213
rect 2777 18204 2789 18207
rect 2740 18176 2789 18204
rect 2740 18164 2746 18176
rect 2777 18173 2789 18176
rect 2823 18204 2835 18207
rect 3044 18207 3102 18213
rect 2823 18176 3004 18204
rect 2823 18173 2835 18176
rect 2777 18167 2835 18173
rect 2976 18136 3004 18176
rect 3044 18173 3056 18207
rect 3090 18204 3102 18207
rect 3510 18204 3516 18216
rect 3090 18176 3516 18204
rect 3090 18173 3102 18176
rect 3044 18167 3102 18173
rect 3510 18164 3516 18176
rect 3568 18164 3574 18216
rect 4709 18207 4767 18213
rect 4709 18173 4721 18207
rect 4755 18204 4767 18207
rect 5350 18204 5356 18216
rect 4755 18176 5356 18204
rect 4755 18173 4767 18176
rect 4709 18167 4767 18173
rect 4062 18136 4068 18148
rect 2976 18108 4068 18136
rect 4062 18096 4068 18108
rect 4120 18136 4126 18148
rect 4724 18136 4752 18167
rect 5350 18164 5356 18176
rect 5408 18164 5414 18216
rect 6638 18164 6644 18216
rect 6696 18204 6702 18216
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6696 18176 6837 18204
rect 6696 18164 6702 18176
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 6825 18167 6883 18173
rect 4120 18108 4752 18136
rect 4120 18096 4126 18108
rect 4890 18096 4896 18148
rect 4948 18145 4954 18148
rect 4948 18139 5012 18145
rect 4948 18105 4966 18139
rect 5000 18105 5012 18139
rect 4948 18099 5012 18105
rect 4948 18096 4954 18099
rect 5534 18096 5540 18148
rect 5592 18136 5598 18148
rect 7098 18136 7104 18148
rect 5592 18108 7104 18136
rect 5592 18096 5598 18108
rect 7098 18096 7104 18108
rect 7156 18096 7162 18148
rect 7852 18145 7880 18232
rect 8748 18207 8806 18213
rect 8748 18173 8760 18207
rect 8794 18204 8806 18207
rect 9214 18204 9220 18216
rect 8794 18176 9220 18204
rect 8794 18173 8806 18176
rect 8748 18167 8806 18173
rect 9214 18164 9220 18176
rect 9272 18164 9278 18216
rect 9953 18207 10011 18213
rect 9953 18173 9965 18207
rect 9999 18204 10011 18207
rect 10137 18207 10195 18213
rect 10137 18204 10149 18207
rect 9999 18176 10149 18204
rect 9999 18173 10011 18176
rect 9953 18167 10011 18173
rect 10137 18173 10149 18176
rect 10183 18173 10195 18207
rect 10137 18167 10195 18173
rect 10410 18164 10416 18216
rect 10468 18204 10474 18216
rect 10468 18176 11836 18204
rect 10468 18164 10474 18176
rect 7837 18139 7895 18145
rect 7208 18108 7604 18136
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 2038 18028 2044 18080
rect 2096 18068 2102 18080
rect 7208 18068 7236 18108
rect 7466 18068 7472 18080
rect 2096 18040 7236 18068
rect 7427 18040 7472 18068
rect 2096 18028 2102 18040
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 7576 18068 7604 18108
rect 7837 18105 7849 18139
rect 7883 18105 7895 18139
rect 7837 18099 7895 18105
rect 8018 18096 8024 18148
rect 8076 18136 8082 18148
rect 11698 18136 11704 18148
rect 8076 18108 11704 18136
rect 8076 18096 8082 18108
rect 11698 18096 11704 18108
rect 11756 18096 11762 18148
rect 11808 18136 11836 18176
rect 12434 18164 12440 18216
rect 12492 18204 12498 18216
rect 13173 18207 13231 18213
rect 12492 18176 12537 18204
rect 12492 18164 12498 18176
rect 13173 18173 13185 18207
rect 13219 18173 13231 18207
rect 13173 18167 13231 18173
rect 13188 18136 13216 18167
rect 11808 18108 13216 18136
rect 7742 18068 7748 18080
rect 7576 18040 7748 18068
rect 7742 18028 7748 18040
rect 7800 18068 7806 18080
rect 7929 18071 7987 18077
rect 7929 18068 7941 18071
rect 7800 18040 7941 18068
rect 7800 18028 7806 18040
rect 7929 18037 7941 18040
rect 7975 18037 7987 18071
rect 7929 18031 7987 18037
rect 8294 18028 8300 18080
rect 8352 18068 8358 18080
rect 9953 18071 10011 18077
rect 9953 18068 9965 18071
rect 8352 18040 9965 18068
rect 8352 18028 8358 18040
rect 9953 18037 9965 18040
rect 9999 18037 10011 18071
rect 11146 18068 11152 18080
rect 11107 18040 11152 18068
rect 9953 18031 10011 18037
rect 11146 18028 11152 18040
rect 11204 18028 11210 18080
rect 12066 18028 12072 18080
rect 12124 18068 12130 18080
rect 12342 18068 12348 18080
rect 12124 18040 12348 18068
rect 12124 18028 12130 18040
rect 12342 18028 12348 18040
rect 12400 18028 12406 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 2958 17864 2964 17876
rect 1728 17836 2964 17864
rect 1728 17824 1734 17836
rect 2958 17824 2964 17836
rect 3016 17824 3022 17876
rect 3510 17824 3516 17876
rect 3568 17864 3574 17876
rect 4249 17867 4307 17873
rect 4249 17864 4261 17867
rect 3568 17836 4261 17864
rect 3568 17824 3574 17836
rect 4249 17833 4261 17836
rect 4295 17833 4307 17867
rect 4249 17827 4307 17833
rect 4706 17824 4712 17876
rect 4764 17864 4770 17876
rect 4801 17867 4859 17873
rect 4801 17864 4813 17867
rect 4764 17836 4813 17864
rect 4764 17824 4770 17836
rect 4801 17833 4813 17836
rect 4847 17833 4859 17867
rect 4801 17827 4859 17833
rect 5261 17867 5319 17873
rect 5261 17833 5273 17867
rect 5307 17864 5319 17867
rect 5534 17864 5540 17876
rect 5307 17836 5540 17864
rect 5307 17833 5319 17836
rect 5261 17827 5319 17833
rect 5534 17824 5540 17836
rect 5592 17824 5598 17876
rect 6089 17867 6147 17873
rect 6089 17833 6101 17867
rect 6135 17864 6147 17867
rect 6914 17864 6920 17876
rect 6135 17836 6920 17864
rect 6135 17833 6147 17836
rect 6089 17827 6147 17833
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 7009 17867 7067 17873
rect 7009 17833 7021 17867
rect 7055 17864 7067 17867
rect 11698 17864 11704 17876
rect 7055 17836 11704 17864
rect 7055 17833 7067 17836
rect 7009 17827 7067 17833
rect 11698 17824 11704 17836
rect 11756 17824 11762 17876
rect 11974 17864 11980 17876
rect 11935 17836 11980 17864
rect 11974 17824 11980 17836
rect 12032 17864 12038 17876
rect 14737 17867 14795 17873
rect 12032 17836 12848 17864
rect 12032 17824 12038 17836
rect 2056 17768 5764 17796
rect 2056 17737 2084 17768
rect 1489 17731 1547 17737
rect 1489 17697 1501 17731
rect 1535 17697 1547 17731
rect 1489 17691 1547 17697
rect 2041 17731 2099 17737
rect 2041 17697 2053 17731
rect 2087 17697 2099 17731
rect 2314 17728 2320 17740
rect 2275 17700 2320 17728
rect 2041 17691 2099 17697
rect 1504 17592 1532 17691
rect 2314 17688 2320 17700
rect 2372 17688 2378 17740
rect 2777 17731 2835 17737
rect 2777 17697 2789 17731
rect 2823 17697 2835 17731
rect 2777 17691 2835 17697
rect 2792 17592 2820 17691
rect 3234 17688 3240 17740
rect 3292 17728 3298 17740
rect 4065 17731 4123 17737
rect 4065 17728 4077 17731
rect 3292 17700 4077 17728
rect 3292 17688 3298 17700
rect 4065 17697 4077 17700
rect 4111 17697 4123 17731
rect 5166 17728 5172 17740
rect 5127 17700 5172 17728
rect 4065 17691 4123 17697
rect 5166 17688 5172 17700
rect 5224 17688 5230 17740
rect 5736 17728 5764 17768
rect 5810 17756 5816 17808
rect 5868 17796 5874 17808
rect 6549 17799 6607 17805
rect 6549 17796 6561 17799
rect 5868 17768 6561 17796
rect 5868 17756 5874 17768
rect 6549 17765 6561 17768
rect 6595 17765 6607 17799
rect 6549 17759 6607 17765
rect 7834 17756 7840 17808
rect 7892 17796 7898 17808
rect 9493 17799 9551 17805
rect 9493 17796 9505 17799
rect 7892 17768 9505 17796
rect 7892 17756 7898 17768
rect 9493 17765 9505 17768
rect 9539 17765 9551 17799
rect 9766 17796 9772 17808
rect 9493 17759 9551 17765
rect 9692 17768 9772 17796
rect 5997 17731 6055 17737
rect 5997 17728 6009 17731
rect 5736 17700 6009 17728
rect 5997 17697 6009 17700
rect 6043 17697 6055 17731
rect 5997 17691 6055 17697
rect 6362 17688 6368 17740
rect 6420 17728 6426 17740
rect 6457 17731 6515 17737
rect 6457 17728 6469 17731
rect 6420 17700 6469 17728
rect 6420 17688 6426 17700
rect 6457 17697 6469 17700
rect 6503 17697 6515 17731
rect 6457 17691 6515 17697
rect 7101 17731 7159 17737
rect 7101 17697 7113 17731
rect 7147 17728 7159 17731
rect 7190 17728 7196 17740
rect 7147 17700 7196 17728
rect 7147 17697 7159 17700
rect 7101 17691 7159 17697
rect 7190 17688 7196 17700
rect 7248 17688 7254 17740
rect 7368 17731 7426 17737
rect 7368 17697 7380 17731
rect 7414 17728 7426 17731
rect 8202 17728 8208 17740
rect 7414 17700 8208 17728
rect 7414 17697 7426 17700
rect 7368 17691 7426 17697
rect 8202 17688 8208 17700
rect 8260 17688 8266 17740
rect 8754 17728 8760 17740
rect 8715 17700 8760 17728
rect 8754 17688 8760 17700
rect 8812 17688 8818 17740
rect 9692 17737 9720 17768
rect 9766 17756 9772 17768
rect 9824 17756 9830 17808
rect 10864 17799 10922 17805
rect 10864 17765 10876 17799
rect 10910 17796 10922 17799
rect 11054 17796 11060 17808
rect 10910 17768 11060 17796
rect 10910 17765 10922 17768
rect 10864 17759 10922 17765
rect 11054 17756 11060 17768
rect 11112 17756 11118 17808
rect 12069 17799 12127 17805
rect 12069 17796 12081 17799
rect 11164 17768 12081 17796
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17697 9735 17731
rect 11164 17728 11192 17768
rect 12069 17765 12081 17768
rect 12115 17765 12127 17799
rect 12069 17759 12127 17765
rect 12621 17731 12679 17737
rect 12621 17728 12633 17731
rect 9677 17691 9735 17697
rect 9784 17700 11192 17728
rect 11604 17700 12633 17728
rect 2958 17660 2964 17672
rect 2919 17632 2964 17660
rect 2958 17620 2964 17632
rect 3016 17620 3022 17672
rect 3513 17663 3571 17669
rect 3513 17629 3525 17663
rect 3559 17660 3571 17663
rect 3602 17660 3608 17672
rect 3559 17632 3608 17660
rect 3559 17629 3571 17632
rect 3513 17623 3571 17629
rect 3602 17620 3608 17632
rect 3660 17620 3666 17672
rect 5442 17660 5448 17672
rect 5403 17632 5448 17660
rect 5442 17620 5448 17632
rect 5500 17620 5506 17672
rect 6733 17663 6791 17669
rect 6733 17629 6745 17663
rect 6779 17660 6791 17663
rect 6914 17660 6920 17672
rect 6779 17632 6920 17660
rect 6779 17629 6791 17632
rect 6733 17623 6791 17629
rect 6914 17620 6920 17632
rect 6972 17620 6978 17672
rect 9784 17660 9812 17700
rect 8119 17632 9812 17660
rect 3050 17592 3056 17604
rect 1504 17564 2728 17592
rect 2792 17564 3056 17592
rect 1670 17524 1676 17536
rect 1631 17496 1676 17524
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 2700 17524 2728 17564
rect 3050 17552 3056 17564
rect 3108 17552 3114 17604
rect 7009 17595 7067 17601
rect 7009 17592 7021 17595
rect 5920 17564 7021 17592
rect 5920 17524 5948 17564
rect 7009 17561 7021 17564
rect 7055 17561 7067 17595
rect 7009 17555 7067 17561
rect 2700 17496 5948 17524
rect 5997 17527 6055 17533
rect 5997 17493 6009 17527
rect 6043 17524 6055 17527
rect 8119 17524 8147 17632
rect 10134 17620 10140 17672
rect 10192 17660 10198 17672
rect 10594 17660 10600 17672
rect 10192 17632 10600 17660
rect 10192 17620 10198 17632
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 8481 17595 8539 17601
rect 8481 17561 8493 17595
rect 8527 17592 8539 17595
rect 9766 17592 9772 17604
rect 8527 17564 9772 17592
rect 8527 17561 8539 17564
rect 8481 17555 8539 17561
rect 9766 17552 9772 17564
rect 9824 17552 9830 17604
rect 6043 17496 8147 17524
rect 6043 17493 6055 17496
rect 5997 17487 6055 17493
rect 8294 17484 8300 17536
rect 8352 17524 8358 17536
rect 8941 17527 8999 17533
rect 8941 17524 8953 17527
rect 8352 17496 8953 17524
rect 8352 17484 8358 17496
rect 8941 17493 8953 17496
rect 8987 17493 8999 17527
rect 8941 17487 8999 17493
rect 9493 17527 9551 17533
rect 9493 17493 9505 17527
rect 9539 17524 9551 17527
rect 9861 17527 9919 17533
rect 9861 17524 9873 17527
rect 9539 17496 9873 17524
rect 9539 17493 9551 17496
rect 9493 17487 9551 17493
rect 9861 17493 9873 17496
rect 9907 17493 9919 17527
rect 9861 17487 9919 17493
rect 10870 17484 10876 17536
rect 10928 17524 10934 17536
rect 11604 17524 11632 17700
rect 12621 17697 12633 17700
rect 12667 17697 12679 17731
rect 12621 17691 12679 17697
rect 11882 17620 11888 17672
rect 11940 17660 11946 17672
rect 12820 17669 12848 17836
rect 14737 17833 14749 17867
rect 14783 17864 14795 17867
rect 19334 17864 19340 17876
rect 14783 17836 19340 17864
rect 14783 17833 14795 17836
rect 14737 17827 14795 17833
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 13265 17731 13323 17737
rect 13265 17697 13277 17731
rect 13311 17697 13323 17731
rect 13265 17691 13323 17697
rect 12713 17663 12771 17669
rect 12713 17660 12725 17663
rect 11940 17632 12725 17660
rect 11940 17620 11946 17632
rect 12713 17629 12725 17632
rect 12759 17629 12771 17663
rect 12713 17623 12771 17629
rect 12805 17663 12863 17669
rect 12805 17629 12817 17663
rect 12851 17629 12863 17663
rect 12805 17623 12863 17629
rect 12069 17595 12127 17601
rect 12069 17561 12081 17595
rect 12115 17592 12127 17595
rect 12253 17595 12311 17601
rect 12253 17592 12265 17595
rect 12115 17564 12265 17592
rect 12115 17561 12127 17564
rect 12069 17555 12127 17561
rect 12253 17561 12265 17564
rect 12299 17561 12311 17595
rect 12253 17555 12311 17561
rect 12342 17552 12348 17604
rect 12400 17592 12406 17604
rect 13280 17592 13308 17691
rect 14458 17688 14464 17740
rect 14516 17728 14522 17740
rect 14553 17731 14611 17737
rect 14553 17728 14565 17731
rect 14516 17700 14565 17728
rect 14516 17688 14522 17700
rect 14553 17697 14565 17700
rect 14599 17697 14611 17731
rect 14553 17691 14611 17697
rect 12400 17564 13308 17592
rect 13449 17595 13507 17601
rect 12400 17552 12406 17564
rect 13449 17561 13461 17595
rect 13495 17592 13507 17595
rect 22002 17592 22008 17604
rect 13495 17564 22008 17592
rect 13495 17561 13507 17564
rect 13449 17555 13507 17561
rect 22002 17552 22008 17564
rect 22060 17552 22066 17604
rect 10928 17496 11632 17524
rect 10928 17484 10934 17496
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 5721 17323 5779 17329
rect 5721 17320 5733 17323
rect 1504 17292 5733 17320
rect 1504 17125 1532 17292
rect 5721 17289 5733 17292
rect 5767 17289 5779 17323
rect 8202 17320 8208 17332
rect 5721 17283 5779 17289
rect 6380 17292 8208 17320
rect 3697 17255 3755 17261
rect 3697 17221 3709 17255
rect 3743 17252 3755 17255
rect 3743 17224 6316 17252
rect 3743 17221 3755 17224
rect 3697 17215 3755 17221
rect 1578 17144 1584 17196
rect 1636 17184 1642 17196
rect 1673 17187 1731 17193
rect 1673 17184 1685 17187
rect 1636 17156 1685 17184
rect 1636 17144 1642 17156
rect 1673 17153 1685 17156
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 1762 17144 1768 17196
rect 1820 17184 1826 17196
rect 2409 17187 2467 17193
rect 2409 17184 2421 17187
rect 1820 17156 2421 17184
rect 1820 17144 1826 17156
rect 2409 17153 2421 17156
rect 2455 17153 2467 17187
rect 3234 17184 3240 17196
rect 3195 17156 3240 17184
rect 2409 17147 2467 17153
rect 3234 17144 3240 17156
rect 3292 17144 3298 17196
rect 4246 17184 4252 17196
rect 4207 17156 4252 17184
rect 4246 17144 4252 17156
rect 4304 17144 4310 17196
rect 5353 17187 5411 17193
rect 5353 17153 5365 17187
rect 5399 17184 5411 17187
rect 5902 17184 5908 17196
rect 5399 17156 5908 17184
rect 5399 17153 5411 17156
rect 5353 17147 5411 17153
rect 5902 17144 5908 17156
rect 5960 17144 5966 17196
rect 1489 17119 1547 17125
rect 1489 17085 1501 17119
rect 1535 17085 1547 17119
rect 2222 17116 2228 17128
rect 2183 17088 2228 17116
rect 1489 17079 1547 17085
rect 2222 17076 2228 17088
rect 2280 17076 2286 17128
rect 2961 17119 3019 17125
rect 2961 17085 2973 17119
rect 3007 17085 3019 17119
rect 2961 17079 3019 17085
rect 2976 17048 3004 17079
rect 4062 17076 4068 17128
rect 4120 17116 4126 17128
rect 4157 17119 4215 17125
rect 4157 17116 4169 17119
rect 4120 17088 4169 17116
rect 4120 17076 4126 17088
rect 4157 17085 4169 17088
rect 4203 17085 4215 17119
rect 4157 17079 4215 17085
rect 6288 17048 6316 17224
rect 6380 17193 6408 17292
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 13633 17323 13691 17329
rect 8496 17292 11100 17320
rect 8496 17252 8524 17292
rect 8036 17224 8524 17252
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17153 6423 17187
rect 6365 17147 6423 17153
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 6914 17116 6920 17128
rect 6871 17088 6920 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 6914 17076 6920 17088
rect 6972 17076 6978 17128
rect 8036 17116 8064 17224
rect 9674 17212 9680 17264
rect 9732 17252 9738 17264
rect 9861 17255 9919 17261
rect 9861 17252 9873 17255
rect 9732 17224 9873 17252
rect 9732 17212 9738 17224
rect 9861 17221 9873 17224
rect 9907 17221 9919 17255
rect 11072 17252 11100 17292
rect 13633 17289 13645 17323
rect 13679 17320 13691 17323
rect 14090 17320 14096 17332
rect 13679 17292 14096 17320
rect 13679 17289 13691 17292
rect 13633 17283 13691 17289
rect 14090 17280 14096 17292
rect 14148 17280 14154 17332
rect 12434 17252 12440 17264
rect 11072 17224 12440 17252
rect 9861 17215 9919 17221
rect 7024 17088 8064 17116
rect 8481 17119 8539 17125
rect 7024 17048 7052 17088
rect 8481 17085 8493 17119
rect 8527 17085 8539 17119
rect 8481 17079 8539 17085
rect 7098 17057 7104 17060
rect 2976 17020 4752 17048
rect 6288 17020 7052 17048
rect 3510 16940 3516 16992
rect 3568 16980 3574 16992
rect 4724 16989 4752 17020
rect 7092 17011 7104 17057
rect 7156 17048 7162 17060
rect 7156 17020 7192 17048
rect 7098 17008 7104 17011
rect 7156 17008 7162 17020
rect 7282 17008 7288 17060
rect 7340 17048 7346 17060
rect 8496 17048 8524 17079
rect 7340 17020 8524 17048
rect 8748 17051 8806 17057
rect 7340 17008 7346 17020
rect 8748 17017 8760 17051
rect 8794 17048 8806 17051
rect 9766 17048 9772 17060
rect 8794 17020 9772 17048
rect 8794 17017 8806 17020
rect 8748 17011 8806 17017
rect 9766 17008 9772 17020
rect 9824 17008 9830 17060
rect 9876 17048 9904 17215
rect 12434 17212 12440 17224
rect 12492 17212 12498 17264
rect 10134 17184 10140 17196
rect 10095 17156 10140 17184
rect 10134 17144 10140 17156
rect 10192 17144 10198 17196
rect 11146 17144 11152 17196
rect 11204 17184 11210 17196
rect 11793 17187 11851 17193
rect 11793 17184 11805 17187
rect 11204 17156 11805 17184
rect 11204 17144 11210 17156
rect 11793 17153 11805 17156
rect 11839 17153 11851 17187
rect 14458 17184 14464 17196
rect 11793 17147 11851 17153
rect 13096 17156 14464 17184
rect 10226 17076 10232 17128
rect 10284 17116 10290 17128
rect 13096 17116 13124 17156
rect 14458 17144 14464 17156
rect 14516 17144 14522 17196
rect 10284 17088 13124 17116
rect 10284 17076 10290 17088
rect 13170 17076 13176 17128
rect 13228 17116 13234 17128
rect 13449 17119 13507 17125
rect 13449 17116 13461 17119
rect 13228 17088 13461 17116
rect 13228 17076 13234 17088
rect 13449 17085 13461 17088
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 10382 17051 10440 17057
rect 10382 17048 10394 17051
rect 9876 17020 10394 17048
rect 10382 17017 10394 17020
rect 10428 17017 10440 17051
rect 10382 17011 10440 17017
rect 11054 17008 11060 17060
rect 11112 17048 11118 17060
rect 11112 17020 11560 17048
rect 11112 17008 11118 17020
rect 4065 16983 4123 16989
rect 4065 16980 4077 16983
rect 3568 16952 4077 16980
rect 3568 16940 3574 16952
rect 4065 16949 4077 16952
rect 4111 16949 4123 16983
rect 4065 16943 4123 16949
rect 4709 16983 4767 16989
rect 4709 16949 4721 16983
rect 4755 16949 4767 16983
rect 5074 16980 5080 16992
rect 5035 16952 5080 16980
rect 4709 16943 4767 16949
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 5169 16983 5227 16989
rect 5169 16949 5181 16983
rect 5215 16980 5227 16983
rect 5626 16980 5632 16992
rect 5215 16952 5632 16980
rect 5215 16949 5227 16952
rect 5169 16943 5227 16949
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 6086 16980 6092 16992
rect 6047 16952 6092 16980
rect 6086 16940 6092 16952
rect 6144 16940 6150 16992
rect 6181 16983 6239 16989
rect 6181 16949 6193 16983
rect 6227 16980 6239 16983
rect 7374 16980 7380 16992
rect 6227 16952 7380 16980
rect 6227 16949 6239 16952
rect 6181 16943 6239 16949
rect 7374 16940 7380 16952
rect 7432 16940 7438 16992
rect 7650 16940 7656 16992
rect 7708 16980 7714 16992
rect 11422 16980 11428 16992
rect 7708 16952 11428 16980
rect 7708 16940 7714 16952
rect 11422 16940 11428 16952
rect 11480 16940 11486 16992
rect 11532 16989 11560 17020
rect 11517 16983 11575 16989
rect 11517 16949 11529 16983
rect 11563 16949 11575 16983
rect 11517 16943 11575 16949
rect 11606 16940 11612 16992
rect 11664 16980 11670 16992
rect 12437 16983 12495 16989
rect 12437 16980 12449 16983
rect 11664 16952 12449 16980
rect 11664 16940 11670 16952
rect 12437 16949 12449 16952
rect 12483 16949 12495 16983
rect 12437 16943 12495 16949
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 2222 16736 2228 16788
rect 2280 16776 2286 16788
rect 2961 16779 3019 16785
rect 2961 16776 2973 16779
rect 2280 16748 2973 16776
rect 2280 16736 2286 16748
rect 2961 16745 2973 16748
rect 3007 16745 3019 16779
rect 2961 16739 3019 16745
rect 3421 16779 3479 16785
rect 3421 16745 3433 16779
rect 3467 16776 3479 16779
rect 7098 16776 7104 16788
rect 3467 16748 6101 16776
rect 7059 16748 7104 16776
rect 3467 16745 3479 16748
rect 3421 16739 3479 16745
rect 2774 16708 2780 16720
rect 1504 16680 2780 16708
rect 1504 16649 1532 16680
rect 2774 16668 2780 16680
rect 2832 16668 2838 16720
rect 3050 16668 3056 16720
rect 3108 16708 3114 16720
rect 3108 16680 5856 16708
rect 3108 16668 3114 16680
rect 1489 16643 1547 16649
rect 1489 16609 1501 16643
rect 1535 16609 1547 16643
rect 1489 16603 1547 16609
rect 2041 16643 2099 16649
rect 2041 16609 2053 16643
rect 2087 16640 2099 16643
rect 2314 16640 2320 16652
rect 2087 16612 2320 16640
rect 2087 16609 2099 16612
rect 2041 16603 2099 16609
rect 2314 16600 2320 16612
rect 2372 16600 2378 16652
rect 2958 16600 2964 16652
rect 3016 16640 3022 16652
rect 3329 16643 3387 16649
rect 3329 16640 3341 16643
rect 3016 16612 3341 16640
rect 3016 16600 3022 16612
rect 3329 16609 3341 16612
rect 3375 16609 3387 16643
rect 4154 16640 4160 16652
rect 3329 16603 3387 16609
rect 3988 16612 4160 16640
rect 2222 16572 2228 16584
rect 2183 16544 2228 16572
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 3605 16575 3663 16581
rect 3605 16541 3617 16575
rect 3651 16572 3663 16575
rect 3988 16572 4016 16612
rect 4154 16600 4160 16612
rect 4212 16640 4218 16652
rect 4321 16643 4379 16649
rect 4321 16640 4333 16643
rect 4212 16612 4333 16640
rect 4212 16600 4218 16612
rect 4321 16609 4333 16612
rect 4367 16609 4379 16643
rect 5828 16640 5856 16680
rect 5902 16668 5908 16720
rect 5960 16717 5966 16720
rect 5960 16711 6024 16717
rect 5960 16677 5978 16711
rect 6012 16677 6024 16711
rect 6073 16708 6101 16748
rect 7098 16736 7104 16748
rect 7156 16736 7162 16788
rect 7374 16776 7380 16788
rect 7335 16748 7380 16776
rect 7374 16736 7380 16748
rect 7432 16736 7438 16788
rect 8389 16779 8447 16785
rect 8389 16745 8401 16779
rect 8435 16745 8447 16779
rect 8846 16776 8852 16788
rect 8759 16748 8852 16776
rect 8389 16739 8447 16745
rect 7285 16711 7343 16717
rect 7285 16708 7297 16711
rect 6073 16680 7297 16708
rect 5960 16671 6024 16677
rect 7285 16677 7297 16680
rect 7331 16677 7343 16711
rect 8404 16708 8432 16739
rect 8846 16736 8852 16748
rect 8904 16776 8910 16788
rect 9950 16776 9956 16788
rect 8904 16748 9956 16776
rect 8904 16736 8910 16748
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 10042 16736 10048 16788
rect 10100 16776 10106 16788
rect 10870 16776 10876 16788
rect 10100 16748 10145 16776
rect 10831 16748 10876 16776
rect 10100 16736 10106 16748
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 11241 16779 11299 16785
rect 11241 16745 11253 16779
rect 11287 16776 11299 16779
rect 11606 16776 11612 16788
rect 11287 16748 11612 16776
rect 11287 16745 11299 16748
rect 11241 16739 11299 16745
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 11882 16776 11888 16788
rect 11843 16748 11888 16776
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12250 16736 12256 16788
rect 12308 16776 12314 16788
rect 12345 16779 12403 16785
rect 12345 16776 12357 16779
rect 12308 16748 12357 16776
rect 12308 16736 12314 16748
rect 12345 16745 12357 16748
rect 12391 16745 12403 16779
rect 12345 16739 12403 16745
rect 10226 16708 10232 16720
rect 7285 16671 7343 16677
rect 7659 16680 8432 16708
rect 8680 16680 10232 16708
rect 5960 16668 5966 16671
rect 7374 16640 7380 16652
rect 5828 16612 7380 16640
rect 4321 16603 4379 16609
rect 7374 16600 7380 16612
rect 7432 16600 7438 16652
rect 3651 16544 4016 16572
rect 4065 16575 4123 16581
rect 3651 16541 3663 16544
rect 3605 16535 3663 16541
rect 4065 16541 4077 16575
rect 4111 16541 4123 16575
rect 4065 16535 4123 16541
rect 3970 16464 3976 16516
rect 4028 16504 4034 16516
rect 4080 16504 4108 16535
rect 5534 16532 5540 16584
rect 5592 16572 5598 16584
rect 5721 16575 5779 16581
rect 5721 16572 5733 16575
rect 5592 16544 5733 16572
rect 5592 16532 5598 16544
rect 5721 16541 5733 16544
rect 5767 16541 5779 16575
rect 5721 16535 5779 16541
rect 7285 16575 7343 16581
rect 7285 16541 7297 16575
rect 7331 16572 7343 16575
rect 7659 16572 7687 16680
rect 7745 16643 7803 16649
rect 7745 16609 7757 16643
rect 7791 16640 7803 16643
rect 8680 16640 8708 16680
rect 10226 16668 10232 16680
rect 10284 16668 10290 16720
rect 11514 16708 11520 16720
rect 11072 16680 11520 16708
rect 7791 16612 8708 16640
rect 7791 16609 7803 16612
rect 7745 16603 7803 16609
rect 8754 16600 8760 16652
rect 8812 16640 8818 16652
rect 8812 16612 8857 16640
rect 8812 16600 8818 16612
rect 9030 16600 9036 16652
rect 9088 16640 9094 16652
rect 11072 16640 11100 16680
rect 11514 16668 11520 16680
rect 11572 16668 11578 16720
rect 13170 16708 13176 16720
rect 13131 16680 13176 16708
rect 13170 16668 13176 16680
rect 13228 16668 13234 16720
rect 9088 16612 11100 16640
rect 9088 16600 9094 16612
rect 11146 16600 11152 16652
rect 11204 16640 11210 16652
rect 11333 16643 11391 16649
rect 11333 16640 11345 16643
rect 11204 16612 11345 16640
rect 11204 16600 11210 16612
rect 11333 16609 11345 16612
rect 11379 16609 11391 16643
rect 11333 16603 11391 16609
rect 11790 16600 11796 16652
rect 11848 16640 11854 16652
rect 12253 16643 12311 16649
rect 12253 16640 12265 16643
rect 11848 16612 12265 16640
rect 11848 16600 11854 16612
rect 12253 16609 12265 16612
rect 12299 16640 12311 16643
rect 12342 16640 12348 16652
rect 12299 16612 12348 16640
rect 12299 16609 12311 16612
rect 12253 16603 12311 16609
rect 12342 16600 12348 16612
rect 12400 16600 12406 16652
rect 12618 16600 12624 16652
rect 12676 16640 12682 16652
rect 12897 16643 12955 16649
rect 12897 16640 12909 16643
rect 12676 16612 12909 16640
rect 12676 16600 12682 16612
rect 12897 16609 12909 16612
rect 12943 16609 12955 16643
rect 12897 16603 12955 16609
rect 7834 16572 7840 16584
rect 7331 16544 7687 16572
rect 7795 16544 7840 16572
rect 7331 16541 7343 16544
rect 7285 16535 7343 16541
rect 7834 16532 7840 16544
rect 7892 16532 7898 16584
rect 8021 16575 8079 16581
rect 8021 16541 8033 16575
rect 8067 16541 8079 16575
rect 8021 16535 8079 16541
rect 8941 16575 8999 16581
rect 8941 16541 8953 16575
rect 8987 16541 8999 16575
rect 10137 16575 10195 16581
rect 10137 16572 10149 16575
rect 8941 16535 8999 16541
rect 9508 16544 10149 16572
rect 4028 16476 4108 16504
rect 4028 16464 4034 16476
rect 7098 16464 7104 16516
rect 7156 16504 7162 16516
rect 8036 16504 8064 16535
rect 7156 16476 8064 16504
rect 7156 16464 7162 16476
rect 8754 16464 8760 16516
rect 8812 16504 8818 16516
rect 8956 16504 8984 16535
rect 9508 16504 9536 16544
rect 10137 16541 10149 16544
rect 10183 16541 10195 16575
rect 10318 16572 10324 16584
rect 10279 16544 10324 16572
rect 10137 16535 10195 16541
rect 10318 16532 10324 16544
rect 10376 16532 10382 16584
rect 11054 16532 11060 16584
rect 11112 16572 11118 16584
rect 11425 16575 11483 16581
rect 11425 16572 11437 16575
rect 11112 16544 11437 16572
rect 11112 16532 11118 16544
rect 11425 16541 11437 16544
rect 11471 16572 11483 16575
rect 12437 16575 12495 16581
rect 12437 16572 12449 16575
rect 11471 16544 12449 16572
rect 11471 16541 11483 16544
rect 11425 16535 11483 16541
rect 12437 16541 12449 16544
rect 12483 16541 12495 16575
rect 12437 16535 12495 16541
rect 8812 16476 8984 16504
rect 9048 16476 9536 16504
rect 8812 16464 8818 16476
rect 1670 16436 1676 16448
rect 1631 16408 1676 16436
rect 1670 16396 1676 16408
rect 1728 16396 1734 16448
rect 5442 16436 5448 16448
rect 5403 16408 5448 16436
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 6362 16396 6368 16448
rect 6420 16436 6426 16448
rect 9048 16436 9076 16476
rect 9766 16464 9772 16516
rect 9824 16504 9830 16516
rect 10336 16504 10364 16532
rect 9824 16476 10364 16504
rect 9824 16464 9830 16476
rect 9674 16436 9680 16448
rect 6420 16408 9076 16436
rect 9635 16408 9680 16436
rect 6420 16396 6426 16408
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 3973 16235 4031 16241
rect 3973 16201 3985 16235
rect 4019 16232 4031 16235
rect 4154 16232 4160 16244
rect 4019 16204 4160 16232
rect 4019 16201 4031 16204
rect 3973 16195 4031 16201
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 5629 16235 5687 16241
rect 5629 16201 5641 16235
rect 5675 16232 5687 16235
rect 5902 16232 5908 16244
rect 5675 16204 5908 16232
rect 5675 16201 5687 16204
rect 5629 16195 5687 16201
rect 5902 16192 5908 16204
rect 5960 16192 5966 16244
rect 6086 16192 6092 16244
rect 6144 16232 6150 16244
rect 6825 16235 6883 16241
rect 6825 16232 6837 16235
rect 6144 16204 6837 16232
rect 6144 16192 6150 16204
rect 6825 16201 6837 16204
rect 6871 16201 6883 16235
rect 6825 16195 6883 16201
rect 7374 16192 7380 16244
rect 7432 16232 7438 16244
rect 8757 16235 8815 16241
rect 8757 16232 8769 16235
rect 7432 16204 8769 16232
rect 7432 16192 7438 16204
rect 8757 16201 8769 16204
rect 8803 16201 8815 16235
rect 8757 16195 8815 16201
rect 9214 16192 9220 16244
rect 9272 16232 9278 16244
rect 13817 16235 13875 16241
rect 13817 16232 13829 16235
rect 9272 16204 13829 16232
rect 9272 16192 9278 16204
rect 13817 16201 13829 16204
rect 13863 16201 13875 16235
rect 13817 16195 13875 16201
rect 8386 16164 8392 16176
rect 5920 16136 8392 16164
rect 1854 16028 1860 16040
rect 1815 16000 1860 16028
rect 1854 15988 1860 16000
rect 1912 15988 1918 16040
rect 2593 16031 2651 16037
rect 2593 15997 2605 16031
rect 2639 16028 2651 16031
rect 2682 16028 2688 16040
rect 2639 16000 2688 16028
rect 2639 15997 2651 16000
rect 2593 15991 2651 15997
rect 2682 15988 2688 16000
rect 2740 16028 2746 16040
rect 3970 16028 3976 16040
rect 2740 16000 3976 16028
rect 2740 15988 2746 16000
rect 3970 15988 3976 16000
rect 4028 16028 4034 16040
rect 4154 16028 4160 16040
rect 4028 16000 4160 16028
rect 4028 15988 4034 16000
rect 4154 15988 4160 16000
rect 4212 16028 4218 16040
rect 4249 16031 4307 16037
rect 4249 16028 4261 16031
rect 4212 16000 4261 16028
rect 4212 15988 4218 16000
rect 4249 15997 4261 16000
rect 4295 16028 4307 16031
rect 5534 16028 5540 16040
rect 4295 16000 5540 16028
rect 4295 15997 4307 16000
rect 4249 15991 4307 15997
rect 5534 15988 5540 16000
rect 5592 15988 5598 16040
rect 5920 16037 5948 16136
rect 8386 16124 8392 16136
rect 8444 16124 8450 16176
rect 8573 16167 8631 16173
rect 8573 16133 8585 16167
rect 8619 16164 8631 16167
rect 8619 16136 9720 16164
rect 8619 16133 8631 16136
rect 8573 16127 8631 16133
rect 6086 16056 6092 16108
rect 6144 16096 6150 16108
rect 6144 16068 6776 16096
rect 6144 16056 6150 16068
rect 5905 16031 5963 16037
rect 5905 15997 5917 16031
rect 5951 15997 5963 16031
rect 5905 15991 5963 15997
rect 6178 15988 6184 16040
rect 6236 16028 6242 16040
rect 6641 16031 6699 16037
rect 6641 16028 6653 16031
rect 6236 16000 6653 16028
rect 6236 15988 6242 16000
rect 6641 15997 6653 16000
rect 6687 15997 6699 16031
rect 6748 16028 6776 16068
rect 7098 16056 7104 16108
rect 7156 16096 7162 16108
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 7156 16068 7389 16096
rect 7156 16056 7162 16068
rect 7377 16065 7389 16068
rect 7423 16065 7435 16099
rect 7377 16059 7435 16065
rect 8754 16056 8760 16108
rect 8812 16096 8818 16108
rect 9214 16096 9220 16108
rect 8812 16068 9220 16096
rect 8812 16056 8818 16068
rect 9214 16056 9220 16068
rect 9272 16056 9278 16108
rect 9401 16099 9459 16105
rect 9401 16065 9413 16099
rect 9447 16096 9459 16099
rect 9490 16096 9496 16108
rect 9447 16068 9496 16096
rect 9447 16065 9459 16068
rect 9401 16059 9459 16065
rect 9490 16056 9496 16068
rect 9548 16056 9554 16108
rect 8573 16031 8631 16037
rect 8573 16028 8585 16031
rect 6748 16000 8585 16028
rect 6641 15991 6699 15997
rect 8573 15997 8585 16000
rect 8619 15997 8631 16031
rect 8573 15991 8631 15997
rect 9125 16031 9183 16037
rect 9125 15997 9137 16031
rect 9171 16028 9183 16031
rect 9582 16028 9588 16040
rect 9171 16000 9588 16028
rect 9171 15997 9183 16000
rect 9125 15991 9183 15997
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 9692 16028 9720 16136
rect 9766 16124 9772 16176
rect 9824 16164 9830 16176
rect 10686 16164 10692 16176
rect 9824 16136 10692 16164
rect 9824 16124 9830 16136
rect 10686 16124 10692 16136
rect 10744 16164 10750 16176
rect 10744 16136 12480 16164
rect 10744 16124 10750 16136
rect 10318 16056 10324 16108
rect 10376 16096 10382 16108
rect 11149 16099 11207 16105
rect 11149 16096 11161 16099
rect 10376 16068 11161 16096
rect 10376 16056 10382 16068
rect 11149 16065 11161 16068
rect 11195 16065 11207 16099
rect 11149 16059 11207 16065
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 11793 16099 11851 16105
rect 11793 16096 11805 16099
rect 11756 16068 11805 16096
rect 11756 16056 11762 16068
rect 11793 16065 11805 16068
rect 11839 16065 11851 16099
rect 12452 16096 12480 16136
rect 12452 16068 12572 16096
rect 11793 16059 11851 16065
rect 10226 16028 10232 16040
rect 9692 16000 10232 16028
rect 10226 15988 10232 16000
rect 10284 16028 10290 16040
rect 10502 16028 10508 16040
rect 10284 16000 10508 16028
rect 10284 15988 10290 16000
rect 10502 15988 10508 16000
rect 10560 15988 10566 16040
rect 11330 15988 11336 16040
rect 11388 16028 11394 16040
rect 11609 16031 11667 16037
rect 11609 16028 11621 16031
rect 11388 16000 11621 16028
rect 11388 15988 11394 16000
rect 11609 15997 11621 16000
rect 11655 15997 11667 16031
rect 12434 16028 12440 16040
rect 12395 16000 12440 16028
rect 11609 15991 11667 15997
rect 12434 15988 12440 16000
rect 12492 15988 12498 16040
rect 12544 16028 12572 16068
rect 13998 16028 14004 16040
rect 12544 16000 14004 16028
rect 13998 15988 14004 16000
rect 14056 15988 14062 16040
rect 1486 15920 1492 15972
rect 1544 15960 1550 15972
rect 2133 15963 2191 15969
rect 2133 15960 2145 15963
rect 1544 15932 2145 15960
rect 1544 15920 1550 15932
rect 2133 15929 2145 15932
rect 2179 15929 2191 15963
rect 2133 15923 2191 15929
rect 2860 15963 2918 15969
rect 2860 15929 2872 15963
rect 2906 15960 2918 15963
rect 3602 15960 3608 15972
rect 2906 15932 3608 15960
rect 2906 15929 2918 15932
rect 2860 15923 2918 15929
rect 3602 15920 3608 15932
rect 3660 15920 3666 15972
rect 4516 15963 4574 15969
rect 4516 15929 4528 15963
rect 4562 15960 4574 15963
rect 5442 15960 5448 15972
rect 4562 15932 5448 15960
rect 4562 15929 4574 15932
rect 4516 15923 4574 15929
rect 5442 15920 5448 15932
rect 5500 15920 5506 15972
rect 6914 15960 6920 15972
rect 6472 15932 6920 15960
rect 1397 15895 1455 15901
rect 1397 15861 1409 15895
rect 1443 15892 1455 15895
rect 3326 15892 3332 15904
rect 1443 15864 3332 15892
rect 1443 15861 1455 15864
rect 1397 15855 1455 15861
rect 3326 15852 3332 15864
rect 3384 15852 3390 15904
rect 4982 15852 4988 15904
rect 5040 15892 5046 15904
rect 6472 15901 6500 15932
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 7193 15963 7251 15969
rect 7193 15929 7205 15963
rect 7239 15960 7251 15963
rect 7837 15963 7895 15969
rect 7837 15960 7849 15963
rect 7239 15932 7849 15960
rect 7239 15929 7251 15932
rect 7193 15923 7251 15929
rect 7837 15929 7849 15932
rect 7883 15929 7895 15963
rect 7837 15923 7895 15929
rect 8297 15963 8355 15969
rect 8297 15929 8309 15963
rect 8343 15960 8355 15963
rect 10042 15960 10048 15972
rect 8343 15932 10048 15960
rect 8343 15929 8355 15932
rect 8297 15923 8355 15929
rect 10042 15920 10048 15932
rect 10100 15920 10106 15972
rect 10965 15963 11023 15969
rect 10965 15929 10977 15963
rect 11011 15960 11023 15963
rect 11698 15960 11704 15972
rect 11011 15932 11704 15960
rect 11011 15929 11023 15932
rect 10965 15923 11023 15929
rect 11698 15920 11704 15932
rect 11756 15960 11762 15972
rect 12158 15960 12164 15972
rect 11756 15932 12164 15960
rect 11756 15920 11762 15932
rect 12158 15920 12164 15932
rect 12216 15920 12222 15972
rect 12710 15969 12716 15972
rect 12704 15960 12716 15969
rect 12671 15932 12716 15960
rect 12704 15923 12716 15932
rect 12710 15920 12716 15923
rect 12768 15920 12774 15972
rect 6089 15895 6147 15901
rect 6089 15892 6101 15895
rect 5040 15864 6101 15892
rect 5040 15852 5046 15864
rect 6089 15861 6101 15864
rect 6135 15861 6147 15895
rect 6089 15855 6147 15861
rect 6457 15895 6515 15901
rect 6457 15861 6469 15895
rect 6503 15861 6515 15895
rect 6457 15855 6515 15861
rect 6546 15852 6552 15904
rect 6604 15892 6610 15904
rect 6730 15892 6736 15904
rect 6604 15864 6736 15892
rect 6604 15852 6610 15864
rect 6730 15852 6736 15864
rect 6788 15892 6794 15904
rect 7285 15895 7343 15901
rect 7285 15892 7297 15895
rect 6788 15864 7297 15892
rect 6788 15852 6794 15864
rect 7285 15861 7297 15864
rect 7331 15861 7343 15895
rect 7285 15855 7343 15861
rect 9217 15895 9275 15901
rect 9217 15861 9229 15895
rect 9263 15892 9275 15895
rect 10597 15895 10655 15901
rect 10597 15892 10609 15895
rect 9263 15864 10609 15892
rect 9263 15861 9275 15864
rect 9217 15855 9275 15861
rect 10597 15861 10609 15864
rect 10643 15861 10655 15895
rect 10597 15855 10655 15861
rect 11057 15895 11115 15901
rect 11057 15861 11069 15895
rect 11103 15892 11115 15895
rect 11974 15892 11980 15904
rect 11103 15864 11980 15892
rect 11103 15861 11115 15864
rect 11057 15855 11115 15861
rect 11974 15852 11980 15864
rect 12032 15892 12038 15904
rect 13354 15892 13360 15904
rect 12032 15864 13360 15892
rect 12032 15852 12038 15864
rect 13354 15852 13360 15864
rect 13412 15852 13418 15904
rect 14093 15895 14151 15901
rect 14093 15861 14105 15895
rect 14139 15892 14151 15895
rect 14366 15892 14372 15904
rect 14139 15864 14372 15892
rect 14139 15861 14151 15864
rect 14093 15855 14151 15861
rect 14366 15852 14372 15864
rect 14424 15852 14430 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1578 15688 1584 15700
rect 1539 15660 1584 15688
rect 1578 15648 1584 15660
rect 1636 15648 1642 15700
rect 2038 15648 2044 15700
rect 2096 15688 2102 15700
rect 2409 15691 2467 15697
rect 2409 15688 2421 15691
rect 2096 15660 2421 15688
rect 2096 15648 2102 15660
rect 2409 15657 2421 15660
rect 2455 15657 2467 15691
rect 2958 15688 2964 15700
rect 2919 15660 2964 15688
rect 2409 15651 2467 15657
rect 2958 15648 2964 15660
rect 3016 15648 3022 15700
rect 3326 15688 3332 15700
rect 3287 15660 3332 15688
rect 3326 15648 3332 15660
rect 3384 15648 3390 15700
rect 4801 15691 4859 15697
rect 4801 15657 4813 15691
rect 4847 15688 4859 15691
rect 5074 15688 5080 15700
rect 4847 15660 5080 15688
rect 4847 15657 4859 15660
rect 4801 15651 4859 15657
rect 5074 15648 5080 15660
rect 5132 15648 5138 15700
rect 5626 15648 5632 15700
rect 5684 15688 5690 15700
rect 5813 15691 5871 15697
rect 5813 15688 5825 15691
rect 5684 15660 5825 15688
rect 5684 15648 5690 15660
rect 5813 15657 5825 15660
rect 5859 15657 5871 15691
rect 5813 15651 5871 15657
rect 6086 15648 6092 15700
rect 6144 15688 6150 15700
rect 6273 15691 6331 15697
rect 6273 15688 6285 15691
rect 6144 15660 6285 15688
rect 6144 15648 6150 15660
rect 6273 15657 6285 15660
rect 6319 15657 6331 15691
rect 6273 15651 6331 15657
rect 6917 15691 6975 15697
rect 6917 15657 6929 15691
rect 6963 15688 6975 15691
rect 9398 15688 9404 15700
rect 6963 15660 9404 15688
rect 6963 15657 6975 15660
rect 6917 15651 6975 15657
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 11330 15688 11336 15700
rect 11291 15660 11336 15688
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 11793 15691 11851 15697
rect 11793 15657 11805 15691
rect 11839 15688 11851 15691
rect 12526 15688 12532 15700
rect 11839 15660 12532 15688
rect 11839 15657 11851 15660
rect 11793 15651 11851 15657
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 13725 15691 13783 15697
rect 13725 15657 13737 15691
rect 13771 15657 13783 15691
rect 14366 15688 14372 15700
rect 14327 15660 14372 15688
rect 13725 15651 13783 15657
rect 4341 15623 4399 15629
rect 4341 15620 4353 15623
rect 1412 15592 4353 15620
rect 1412 15561 1440 15592
rect 4341 15589 4353 15592
rect 4387 15589 4399 15623
rect 4341 15583 4399 15589
rect 6181 15623 6239 15629
rect 6181 15589 6193 15623
rect 6227 15620 6239 15623
rect 10686 15620 10692 15632
rect 6227 15592 10692 15620
rect 6227 15589 6239 15592
rect 6181 15583 6239 15589
rect 10686 15580 10692 15592
rect 10744 15620 10750 15632
rect 11882 15620 11888 15632
rect 10744 15592 11888 15620
rect 10744 15580 10750 15592
rect 11882 15580 11888 15592
rect 11940 15580 11946 15632
rect 12710 15620 12716 15632
rect 11992 15592 12716 15620
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15521 1455 15555
rect 1397 15515 1455 15521
rect 2317 15555 2375 15561
rect 2317 15521 2329 15555
rect 2363 15552 2375 15555
rect 2866 15552 2872 15564
rect 2363 15524 2872 15552
rect 2363 15521 2375 15524
rect 2317 15515 2375 15521
rect 2866 15512 2872 15524
rect 2924 15512 2930 15564
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15552 4123 15555
rect 4982 15552 4988 15564
rect 4111 15524 4988 15552
rect 4111 15521 4123 15524
rect 4065 15515 4123 15521
rect 4982 15512 4988 15524
rect 5040 15512 5046 15564
rect 5169 15555 5227 15561
rect 5169 15521 5181 15555
rect 5215 15552 5227 15555
rect 6086 15552 6092 15564
rect 5215 15524 6092 15552
rect 5215 15521 5227 15524
rect 5169 15515 5227 15521
rect 6086 15512 6092 15524
rect 6144 15512 6150 15564
rect 7282 15552 7288 15564
rect 7243 15524 7288 15552
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 8202 15561 8208 15564
rect 8196 15515 8208 15561
rect 8260 15552 8266 15564
rect 8260 15524 8296 15552
rect 8202 15512 8208 15515
rect 8260 15512 8266 15524
rect 9030 15512 9036 15564
rect 9088 15552 9094 15564
rect 9677 15555 9735 15561
rect 9677 15552 9689 15555
rect 9088 15524 9689 15552
rect 9088 15512 9094 15524
rect 9677 15521 9689 15524
rect 9723 15521 9735 15555
rect 9933 15555 9991 15561
rect 9933 15552 9945 15555
rect 9677 15515 9735 15521
rect 9784 15524 9945 15552
rect 2038 15444 2044 15496
rect 2096 15484 2102 15496
rect 2501 15487 2559 15493
rect 2501 15484 2513 15487
rect 2096 15456 2513 15484
rect 2096 15444 2102 15456
rect 2501 15453 2513 15456
rect 2547 15453 2559 15487
rect 3418 15484 3424 15496
rect 3331 15456 3424 15484
rect 2501 15447 2559 15453
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 3602 15484 3608 15496
rect 3563 15456 3608 15484
rect 3602 15444 3608 15456
rect 3660 15444 3666 15496
rect 5261 15487 5319 15493
rect 5261 15453 5273 15487
rect 5307 15453 5319 15487
rect 5442 15484 5448 15496
rect 5355 15456 5448 15484
rect 5261 15447 5319 15453
rect 3436 15416 3464 15444
rect 4890 15416 4896 15428
rect 3436 15388 4896 15416
rect 4890 15376 4896 15388
rect 4948 15376 4954 15428
rect 5166 15376 5172 15428
rect 5224 15416 5230 15428
rect 5276 15416 5304 15447
rect 5442 15444 5448 15456
rect 5500 15484 5506 15496
rect 6365 15487 6423 15493
rect 6365 15484 6377 15487
rect 5500 15456 6377 15484
rect 5500 15444 5506 15456
rect 6365 15453 6377 15456
rect 6411 15453 6423 15487
rect 6365 15447 6423 15453
rect 7006 15444 7012 15496
rect 7064 15484 7070 15496
rect 7377 15487 7435 15493
rect 7377 15484 7389 15487
rect 7064 15456 7389 15484
rect 7064 15444 7070 15456
rect 7377 15453 7389 15456
rect 7423 15453 7435 15487
rect 7377 15447 7435 15453
rect 7561 15487 7619 15493
rect 7561 15453 7573 15487
rect 7607 15453 7619 15487
rect 7561 15447 7619 15453
rect 5224 15388 5304 15416
rect 5224 15376 5230 15388
rect 1949 15351 2007 15357
rect 1949 15317 1961 15351
rect 1995 15348 2007 15351
rect 3050 15348 3056 15360
rect 1995 15320 3056 15348
rect 1995 15317 2007 15320
rect 1949 15311 2007 15317
rect 3050 15308 3056 15320
rect 3108 15308 3114 15360
rect 3694 15308 3700 15360
rect 3752 15348 3758 15360
rect 5074 15348 5080 15360
rect 3752 15320 5080 15348
rect 3752 15308 3758 15320
rect 5074 15308 5080 15320
rect 5132 15308 5138 15360
rect 5276 15348 5304 15388
rect 5442 15348 5448 15360
rect 5276 15320 5448 15348
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 7576 15348 7604 15447
rect 7834 15444 7840 15496
rect 7892 15484 7898 15496
rect 7929 15487 7987 15493
rect 7929 15484 7941 15487
rect 7892 15456 7941 15484
rect 7892 15444 7898 15456
rect 7929 15453 7941 15456
rect 7975 15453 7987 15487
rect 9784 15484 9812 15524
rect 9933 15521 9945 15524
rect 9979 15521 9991 15555
rect 9933 15515 9991 15521
rect 11701 15555 11759 15561
rect 11701 15521 11713 15555
rect 11747 15521 11759 15555
rect 11701 15515 11759 15521
rect 7929 15447 7987 15453
rect 9324 15456 9812 15484
rect 9122 15348 9128 15360
rect 7576 15320 9128 15348
rect 9122 15308 9128 15320
rect 9180 15348 9186 15360
rect 9324 15357 9352 15456
rect 9309 15351 9367 15357
rect 9309 15348 9321 15351
rect 9180 15320 9321 15348
rect 9180 15308 9186 15320
rect 9309 15317 9321 15320
rect 9355 15317 9367 15351
rect 11054 15348 11060 15360
rect 11015 15320 11060 15348
rect 9309 15311 9367 15317
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 11716 15348 11744 15515
rect 11992 15493 12020 15592
rect 12710 15580 12716 15592
rect 12768 15620 12774 15632
rect 13740 15620 13768 15651
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 12768 15592 13768 15620
rect 12768 15580 12774 15592
rect 13998 15580 14004 15632
rect 14056 15620 14062 15632
rect 14461 15623 14519 15629
rect 14461 15620 14473 15623
rect 14056 15592 14473 15620
rect 14056 15580 14062 15592
rect 14461 15589 14473 15592
rect 14507 15589 14519 15623
rect 14461 15583 14519 15589
rect 12345 15555 12403 15561
rect 12345 15521 12357 15555
rect 12391 15552 12403 15555
rect 12434 15552 12440 15564
rect 12391 15524 12440 15552
rect 12391 15521 12403 15524
rect 12345 15515 12403 15521
rect 12434 15512 12440 15524
rect 12492 15512 12498 15564
rect 12612 15555 12670 15561
rect 12612 15521 12624 15555
rect 12658 15552 12670 15555
rect 14274 15552 14280 15564
rect 12658 15524 14280 15552
rect 12658 15521 12670 15524
rect 12612 15515 12670 15521
rect 14274 15512 14280 15524
rect 14332 15552 14338 15564
rect 14332 15524 14596 15552
rect 14332 15512 14338 15524
rect 14568 15493 14596 15524
rect 11977 15487 12035 15493
rect 11977 15453 11989 15487
rect 12023 15453 12035 15487
rect 11977 15447 12035 15453
rect 14553 15487 14611 15493
rect 14553 15453 14565 15487
rect 14599 15453 14611 15487
rect 14553 15447 14611 15453
rect 14001 15419 14059 15425
rect 14001 15416 14013 15419
rect 13280 15388 14013 15416
rect 13280 15348 13308 15388
rect 14001 15385 14013 15388
rect 14047 15385 14059 15419
rect 14001 15379 14059 15385
rect 11716 15320 13308 15348
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 1578 15144 1584 15156
rect 1539 15116 1584 15144
rect 1578 15104 1584 15116
rect 1636 15104 1642 15156
rect 2866 15104 2872 15156
rect 2924 15144 2930 15156
rect 2924 15116 4108 15144
rect 2924 15104 2930 15116
rect 1949 15079 2007 15085
rect 1949 15045 1961 15079
rect 1995 15076 2007 15079
rect 1995 15048 3004 15076
rect 1995 15045 2007 15048
rect 1949 15039 2007 15045
rect 198 14968 204 15020
rect 256 15008 262 15020
rect 1670 15008 1676 15020
rect 256 14980 1676 15008
rect 256 14968 262 14980
rect 1670 14968 1676 14980
rect 1728 15008 1734 15020
rect 2409 15011 2467 15017
rect 2409 15008 2421 15011
rect 1728 14980 2421 15008
rect 1728 14968 1734 14980
rect 2409 14977 2421 14980
rect 2455 14977 2467 15011
rect 2590 15008 2596 15020
rect 2551 14980 2596 15008
rect 2409 14971 2467 14977
rect 2590 14968 2596 14980
rect 2648 14968 2654 15020
rect 2976 15008 3004 15048
rect 4080 15008 4108 15116
rect 4246 15104 4252 15156
rect 4304 15144 4310 15156
rect 4341 15147 4399 15153
rect 4341 15144 4353 15147
rect 4304 15116 4353 15144
rect 4304 15104 4310 15116
rect 4341 15113 4353 15116
rect 4387 15113 4399 15147
rect 4341 15107 4399 15113
rect 5721 15147 5779 15153
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 7006 15144 7012 15156
rect 5767 15116 7012 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 7742 15104 7748 15156
rect 7800 15104 7806 15156
rect 8202 15144 8208 15156
rect 8115 15116 8208 15144
rect 8202 15104 8208 15116
rect 8260 15144 8266 15156
rect 9490 15144 9496 15156
rect 8260 15116 9496 15144
rect 8260 15104 8266 15116
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 9585 15147 9643 15153
rect 9585 15113 9597 15147
rect 9631 15144 9643 15147
rect 12618 15144 12624 15156
rect 9631 15116 12624 15144
rect 9631 15113 9643 15116
rect 9585 15107 9643 15113
rect 12618 15104 12624 15116
rect 12676 15104 12682 15156
rect 5534 15076 5540 15088
rect 5184 15048 5540 15076
rect 5184 15017 5212 15048
rect 5534 15036 5540 15048
rect 5592 15036 5598 15088
rect 7760 15076 7788 15104
rect 10502 15076 10508 15088
rect 7760 15048 10508 15076
rect 10502 15036 10508 15048
rect 10560 15036 10566 15088
rect 5169 15011 5227 15017
rect 5169 15008 5181 15011
rect 2976 14980 3096 15008
rect 4080 14980 5181 15008
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 1486 14940 1492 14952
rect 1443 14912 1492 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 1486 14900 1492 14912
rect 1544 14900 1550 14952
rect 2130 14900 2136 14952
rect 2188 14940 2194 14952
rect 2958 14940 2964 14952
rect 2188 14912 2964 14940
rect 2188 14900 2194 14912
rect 2958 14900 2964 14912
rect 3016 14900 3022 14952
rect 3068 14940 3096 14980
rect 5169 14977 5181 14980
rect 5215 14977 5227 15011
rect 5350 15008 5356 15020
rect 5263 14980 5356 15008
rect 5169 14971 5227 14977
rect 5350 14968 5356 14980
rect 5408 15008 5414 15020
rect 6365 15011 6423 15017
rect 5408 14980 6316 15008
rect 5408 14968 5414 14980
rect 6181 14943 6239 14949
rect 6181 14940 6193 14943
rect 3068 14912 6193 14940
rect 6181 14909 6193 14912
rect 6227 14909 6239 14943
rect 6288 14940 6316 14980
rect 6365 14977 6377 15011
rect 6411 15008 6423 15011
rect 9122 15008 9128 15020
rect 6411 14980 6960 15008
rect 9083 14980 9128 15008
rect 6411 14977 6423 14980
rect 6365 14971 6423 14977
rect 6932 14952 6960 14980
rect 9122 14968 9128 14980
rect 9180 14968 9186 15020
rect 9398 14968 9404 15020
rect 9456 15008 9462 15020
rect 10045 15011 10103 15017
rect 10045 15008 10057 15011
rect 9456 14980 10057 15008
rect 9456 14968 9462 14980
rect 10045 14977 10057 14980
rect 10091 14977 10103 15011
rect 10045 14971 10103 14977
rect 10229 15011 10287 15017
rect 10229 14977 10241 15011
rect 10275 15008 10287 15011
rect 10275 14980 10732 15008
rect 10275 14977 10287 14980
rect 10229 14971 10287 14977
rect 6641 14943 6699 14949
rect 6641 14940 6653 14943
rect 6288 14912 6653 14940
rect 6181 14903 6239 14909
rect 6641 14909 6653 14912
rect 6687 14909 6699 14943
rect 6822 14940 6828 14952
rect 6783 14912 6828 14940
rect 6641 14903 6699 14909
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 6914 14900 6920 14952
rect 6972 14900 6978 14952
rect 7650 14940 7656 14952
rect 7024 14912 7656 14940
rect 658 14832 664 14884
rect 716 14872 722 14884
rect 2317 14875 2375 14881
rect 2317 14872 2329 14875
rect 716 14844 2329 14872
rect 716 14832 722 14844
rect 2317 14841 2329 14844
rect 2363 14841 2375 14875
rect 2317 14835 2375 14841
rect 3228 14875 3286 14881
rect 3228 14841 3240 14875
rect 3274 14841 3286 14875
rect 3228 14835 3286 14841
rect 2332 14804 2360 14835
rect 2958 14804 2964 14816
rect 2332 14776 2964 14804
rect 2958 14764 2964 14776
rect 3016 14764 3022 14816
rect 3243 14804 3271 14835
rect 3326 14832 3332 14884
rect 3384 14872 3390 14884
rect 6089 14875 6147 14881
rect 6089 14872 6101 14875
rect 3384 14844 6101 14872
rect 3384 14832 3390 14844
rect 6089 14841 6101 14844
rect 6135 14841 6147 14875
rect 7024 14872 7052 14912
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 9490 14940 9496 14952
rect 8496 14912 9496 14940
rect 8496 14884 8524 14912
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 10134 14900 10140 14952
rect 10192 14940 10198 14952
rect 10594 14940 10600 14952
rect 10192 14912 10600 14940
rect 10192 14900 10198 14912
rect 10594 14900 10600 14912
rect 10652 14900 10658 14952
rect 6089 14835 6147 14841
rect 6564 14844 7052 14872
rect 7092 14875 7150 14881
rect 3786 14804 3792 14816
rect 3243 14776 3792 14804
rect 3786 14764 3792 14776
rect 3844 14764 3850 14816
rect 4154 14764 4160 14816
rect 4212 14804 4218 14816
rect 4338 14804 4344 14816
rect 4212 14776 4344 14804
rect 4212 14764 4218 14776
rect 4338 14764 4344 14776
rect 4396 14764 4402 14816
rect 4706 14804 4712 14816
rect 4667 14776 4712 14804
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 5074 14804 5080 14816
rect 5035 14776 5080 14804
rect 5074 14764 5080 14776
rect 5132 14804 5138 14816
rect 6564 14804 6592 14844
rect 7092 14841 7104 14875
rect 7138 14872 7150 14875
rect 8478 14872 8484 14884
rect 7138 14844 8484 14872
rect 7138 14841 7150 14844
rect 7092 14835 7150 14841
rect 5132 14776 6592 14804
rect 6641 14807 6699 14813
rect 5132 14764 5138 14776
rect 6641 14773 6653 14807
rect 6687 14804 6699 14807
rect 7107 14804 7135 14835
rect 8478 14832 8484 14844
rect 8536 14832 8542 14884
rect 9953 14875 10011 14881
rect 9953 14872 9965 14875
rect 8588 14844 9965 14872
rect 8588 14813 8616 14844
rect 9953 14841 9965 14844
rect 9999 14841 10011 14875
rect 10704 14872 10732 14980
rect 12066 14968 12072 15020
rect 12124 15008 12130 15020
rect 12124 14980 12572 15008
rect 12124 14968 12130 14980
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 11164 14912 12449 14940
rect 10864 14875 10922 14881
rect 10864 14872 10876 14875
rect 10704 14844 10876 14872
rect 9953 14835 10011 14841
rect 10864 14841 10876 14844
rect 10910 14872 10922 14875
rect 11054 14872 11060 14884
rect 10910 14844 11060 14872
rect 10910 14841 10922 14844
rect 10864 14835 10922 14841
rect 11054 14832 11060 14844
rect 11112 14832 11118 14884
rect 6687 14776 7135 14804
rect 8573 14807 8631 14813
rect 6687 14773 6699 14776
rect 6641 14767 6699 14773
rect 8573 14773 8585 14807
rect 8619 14773 8631 14807
rect 8938 14804 8944 14816
rect 8899 14776 8944 14804
rect 8573 14767 8631 14773
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 9030 14764 9036 14816
rect 9088 14804 9094 14816
rect 9088 14776 9133 14804
rect 9088 14764 9094 14776
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 11164 14804 11192 14912
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12544 14940 12572 14980
rect 13998 14968 14004 15020
rect 14056 15008 14062 15020
rect 14645 15011 14703 15017
rect 14645 15008 14657 15011
rect 14056 14980 14657 15008
rect 14056 14968 14062 14980
rect 14645 14977 14657 14980
rect 14691 14977 14703 15011
rect 14645 14971 14703 14977
rect 15010 14940 15016 14952
rect 12544 14912 15016 14940
rect 12437 14903 12495 14909
rect 15010 14900 15016 14912
rect 15068 14900 15074 14952
rect 12682 14875 12740 14881
rect 12682 14872 12694 14875
rect 11992 14844 12694 14872
rect 11992 14816 12020 14844
rect 12682 14841 12694 14844
rect 12728 14841 12740 14875
rect 12682 14835 12740 14841
rect 13170 14832 13176 14884
rect 13228 14872 13234 14884
rect 14461 14875 14519 14881
rect 14461 14872 14473 14875
rect 13228 14844 14473 14872
rect 13228 14832 13234 14844
rect 14461 14841 14473 14844
rect 14507 14872 14519 14875
rect 15286 14872 15292 14884
rect 14507 14844 15292 14872
rect 14507 14841 14519 14844
rect 14461 14835 14519 14841
rect 15286 14832 15292 14844
rect 15344 14832 15350 14884
rect 11974 14804 11980 14816
rect 10652 14776 11192 14804
rect 11887 14776 11980 14804
rect 10652 14764 10658 14776
rect 11974 14764 11980 14776
rect 12032 14764 12038 14816
rect 13817 14807 13875 14813
rect 13817 14773 13829 14807
rect 13863 14804 13875 14807
rect 13906 14804 13912 14816
rect 13863 14776 13912 14804
rect 13863 14773 13875 14776
rect 13817 14767 13875 14773
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 14090 14804 14096 14816
rect 14051 14776 14096 14804
rect 14090 14764 14096 14776
rect 14148 14764 14154 14816
rect 14550 14804 14556 14816
rect 14511 14776 14556 14804
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 2961 14603 3019 14609
rect 2961 14569 2973 14603
rect 3007 14600 3019 14603
rect 3142 14600 3148 14612
rect 3007 14572 3148 14600
rect 3007 14569 3019 14572
rect 2961 14563 3019 14569
rect 3142 14560 3148 14572
rect 3200 14560 3206 14612
rect 3970 14600 3976 14612
rect 3344 14572 3976 14600
rect 1762 14492 1768 14544
rect 1820 14532 1826 14544
rect 3344 14541 3372 14572
rect 3970 14560 3976 14572
rect 4028 14560 4034 14612
rect 4706 14560 4712 14612
rect 4764 14600 4770 14612
rect 7009 14603 7067 14609
rect 7009 14600 7021 14603
rect 4764 14572 7021 14600
rect 4764 14560 4770 14572
rect 7009 14569 7021 14572
rect 7055 14569 7067 14603
rect 7009 14563 7067 14569
rect 7101 14603 7159 14609
rect 7101 14569 7113 14603
rect 7147 14600 7159 14603
rect 7466 14600 7472 14612
rect 7147 14572 7472 14600
rect 7147 14569 7159 14572
rect 7101 14563 7159 14569
rect 7466 14560 7472 14572
rect 7524 14560 7530 14612
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 8113 14603 8171 14609
rect 8113 14600 8125 14603
rect 7708 14572 8125 14600
rect 7708 14560 7714 14572
rect 8113 14569 8125 14572
rect 8159 14569 8171 14603
rect 8113 14563 8171 14569
rect 8938 14560 8944 14612
rect 8996 14600 9002 14612
rect 9953 14603 10011 14609
rect 9953 14600 9965 14603
rect 8996 14572 9965 14600
rect 8996 14560 9002 14572
rect 9953 14569 9965 14572
rect 9999 14569 10011 14603
rect 9953 14563 10011 14569
rect 10594 14560 10600 14612
rect 10652 14600 10658 14612
rect 10870 14600 10876 14612
rect 10652 14572 10876 14600
rect 10652 14560 10658 14572
rect 10870 14560 10876 14572
rect 10928 14600 10934 14612
rect 10965 14603 11023 14609
rect 10965 14600 10977 14603
rect 10928 14572 10977 14600
rect 10928 14560 10934 14572
rect 10965 14569 10977 14572
rect 11011 14569 11023 14603
rect 10965 14563 11023 14569
rect 11333 14603 11391 14609
rect 11333 14569 11345 14603
rect 11379 14600 11391 14603
rect 14550 14600 14556 14612
rect 11379 14572 14556 14600
rect 11379 14569 11391 14572
rect 11333 14563 11391 14569
rect 14550 14560 14556 14572
rect 14608 14560 14614 14612
rect 3329 14535 3387 14541
rect 3329 14532 3341 14535
rect 1820 14504 3341 14532
rect 1820 14492 1826 14504
rect 3329 14501 3341 14504
rect 3375 14501 3387 14535
rect 5626 14532 5632 14544
rect 3329 14495 3387 14501
rect 3436 14504 5632 14532
rect 1857 14467 1915 14473
rect 1857 14433 1869 14467
rect 1903 14464 1915 14467
rect 2317 14467 2375 14473
rect 2317 14464 2329 14467
rect 1903 14436 2329 14464
rect 1903 14433 1915 14436
rect 1857 14427 1915 14433
rect 2317 14433 2329 14436
rect 2363 14464 2375 14467
rect 2498 14464 2504 14476
rect 2363 14436 2504 14464
rect 2363 14433 2375 14436
rect 2317 14427 2375 14433
rect 2498 14424 2504 14436
rect 2556 14424 2562 14476
rect 2406 14396 2412 14408
rect 2367 14368 2412 14396
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14396 2651 14399
rect 2682 14396 2688 14408
rect 2639 14368 2688 14396
rect 2639 14365 2651 14368
rect 2593 14359 2651 14365
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 3436 14405 3464 14504
rect 5626 14492 5632 14504
rect 5684 14492 5690 14544
rect 6086 14492 6092 14544
rect 6144 14532 6150 14544
rect 6181 14535 6239 14541
rect 6181 14532 6193 14535
rect 6144 14504 6193 14532
rect 6144 14492 6150 14504
rect 6181 14501 6193 14504
rect 6227 14501 6239 14535
rect 6181 14495 6239 14501
rect 9490 14492 9496 14544
rect 9548 14532 9554 14544
rect 11054 14532 11060 14544
rect 9548 14504 11060 14532
rect 9548 14492 9554 14504
rect 11054 14492 11060 14504
rect 11112 14492 11118 14544
rect 12618 14532 12624 14544
rect 11164 14504 12624 14532
rect 3694 14424 3700 14476
rect 3752 14464 3758 14476
rect 4792 14467 4850 14473
rect 4792 14464 4804 14467
rect 3752 14436 4804 14464
rect 3752 14424 3758 14436
rect 4792 14433 4804 14436
rect 4838 14464 4850 14467
rect 6546 14464 6552 14476
rect 4838 14436 6552 14464
rect 4838 14433 4850 14436
rect 4792 14427 4850 14433
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 8018 14464 8024 14476
rect 7979 14436 8024 14464
rect 8018 14424 8024 14436
rect 8076 14424 8082 14476
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14464 9183 14467
rect 10321 14467 10379 14473
rect 10321 14464 10333 14467
rect 9171 14436 10333 14464
rect 9171 14433 9183 14436
rect 9125 14427 9183 14433
rect 10321 14433 10333 14436
rect 10367 14433 10379 14467
rect 10321 14427 10379 14433
rect 10413 14467 10471 14473
rect 10413 14433 10425 14467
rect 10459 14464 10471 14467
rect 10778 14464 10784 14476
rect 10459 14436 10784 14464
rect 10459 14433 10471 14436
rect 10413 14427 10471 14433
rect 10778 14424 10784 14436
rect 10836 14424 10842 14476
rect 11164 14473 11192 14504
rect 12618 14492 12624 14504
rect 12676 14532 12682 14544
rect 15657 14535 15715 14541
rect 12676 14504 12848 14532
rect 12676 14492 12682 14504
rect 12820 14473 12848 14504
rect 15657 14501 15669 14535
rect 15703 14532 15715 14535
rect 15746 14532 15752 14544
rect 15703 14504 15752 14532
rect 15703 14501 15715 14504
rect 15657 14495 15715 14501
rect 15746 14492 15752 14504
rect 15804 14532 15810 14544
rect 16206 14532 16212 14544
rect 15804 14504 16212 14532
rect 15804 14492 15810 14504
rect 16206 14492 16212 14504
rect 16264 14492 16270 14544
rect 11149 14467 11207 14473
rect 11149 14433 11161 14467
rect 11195 14433 11207 14467
rect 11149 14427 11207 14433
rect 11701 14467 11759 14473
rect 11701 14433 11713 14467
rect 11747 14433 11759 14467
rect 11701 14427 11759 14433
rect 12805 14467 12863 14473
rect 12805 14433 12817 14467
rect 12851 14433 12863 14467
rect 12805 14427 12863 14433
rect 12897 14467 12955 14473
rect 12897 14433 12909 14467
rect 12943 14464 12955 14467
rect 12986 14464 12992 14476
rect 12943 14436 12992 14464
rect 12943 14433 12955 14436
rect 12897 14427 12955 14433
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14396 2927 14399
rect 3421 14399 3479 14405
rect 3421 14396 3433 14399
rect 2915 14368 3433 14396
rect 2915 14365 2927 14368
rect 2869 14359 2927 14365
rect 3421 14365 3433 14368
rect 3467 14365 3479 14399
rect 3602 14396 3608 14408
rect 3563 14368 3608 14396
rect 3421 14359 3479 14365
rect 3602 14356 3608 14368
rect 3660 14356 3666 14408
rect 4338 14356 4344 14408
rect 4396 14396 4402 14408
rect 4525 14399 4583 14405
rect 4525 14396 4537 14399
rect 4396 14368 4537 14396
rect 4396 14356 4402 14368
rect 4525 14365 4537 14368
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 6914 14356 6920 14408
rect 6972 14396 6978 14408
rect 7193 14399 7251 14405
rect 7193 14396 7205 14399
rect 6972 14368 7205 14396
rect 6972 14356 6978 14368
rect 7193 14365 7205 14368
rect 7239 14396 7251 14399
rect 8110 14396 8116 14408
rect 7239 14368 8116 14396
rect 7239 14365 7251 14368
rect 7193 14359 7251 14365
rect 8110 14356 8116 14368
rect 8168 14356 8174 14408
rect 8202 14356 8208 14408
rect 8260 14396 8266 14408
rect 8297 14399 8355 14405
rect 8297 14396 8309 14399
rect 8260 14368 8309 14396
rect 8260 14356 8266 14368
rect 8297 14365 8309 14368
rect 8343 14396 8355 14399
rect 9306 14396 9312 14408
rect 8343 14368 9312 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 9306 14356 9312 14368
rect 9364 14356 9370 14408
rect 9582 14356 9588 14408
rect 9640 14396 9646 14408
rect 10502 14396 10508 14408
rect 9640 14368 10508 14396
rect 9640 14356 9646 14368
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 10594 14356 10600 14408
rect 10652 14396 10658 14408
rect 11716 14396 11744 14427
rect 10652 14368 11744 14396
rect 11793 14399 11851 14405
rect 10652 14356 10658 14368
rect 11793 14365 11805 14399
rect 11839 14365 11851 14399
rect 11974 14396 11980 14408
rect 11935 14368 11980 14396
rect 11793 14359 11851 14365
rect 1949 14331 2007 14337
rect 1949 14297 1961 14331
rect 1995 14328 2007 14331
rect 4154 14328 4160 14340
rect 1995 14300 4160 14328
rect 1995 14297 2007 14300
rect 1949 14291 2007 14297
rect 4154 14288 4160 14300
rect 4212 14288 4218 14340
rect 6641 14331 6699 14337
rect 6641 14297 6653 14331
rect 6687 14328 6699 14331
rect 7282 14328 7288 14340
rect 6687 14300 7288 14328
rect 6687 14297 6699 14300
rect 6641 14291 6699 14297
rect 7282 14288 7288 14300
rect 7340 14288 7346 14340
rect 11808 14328 11836 14359
rect 11974 14356 11980 14368
rect 12032 14356 12038 14408
rect 7383 14300 11836 14328
rect 1118 14220 1124 14272
rect 1176 14260 1182 14272
rect 2869 14263 2927 14269
rect 2869 14260 2881 14263
rect 1176 14232 2881 14260
rect 1176 14220 1182 14232
rect 2869 14229 2881 14232
rect 2915 14229 2927 14263
rect 2869 14223 2927 14229
rect 3602 14220 3608 14272
rect 3660 14260 3666 14272
rect 5905 14263 5963 14269
rect 5905 14260 5917 14263
rect 3660 14232 5917 14260
rect 3660 14220 3666 14232
rect 5905 14229 5917 14232
rect 5951 14229 5963 14263
rect 5905 14223 5963 14229
rect 5994 14220 6000 14272
rect 6052 14260 6058 14272
rect 7383 14260 7411 14300
rect 12434 14288 12440 14340
rect 12492 14328 12498 14340
rect 12621 14331 12679 14337
rect 12621 14328 12633 14331
rect 12492 14300 12633 14328
rect 12492 14288 12498 14300
rect 12621 14297 12633 14300
rect 12667 14328 12679 14331
rect 12912 14328 12940 14427
rect 12986 14424 12992 14436
rect 13044 14424 13050 14476
rect 13164 14467 13222 14473
rect 13164 14433 13176 14467
rect 13210 14464 13222 14467
rect 13446 14464 13452 14476
rect 13210 14436 13452 14464
rect 13210 14433 13222 14436
rect 13164 14427 13222 14433
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 19150 14464 19156 14476
rect 14660 14436 19156 14464
rect 13906 14356 13912 14408
rect 13964 14396 13970 14408
rect 14660 14396 14688 14436
rect 19150 14424 19156 14436
rect 19208 14424 19214 14476
rect 13964 14368 14688 14396
rect 13964 14356 13970 14368
rect 15286 14356 15292 14408
rect 15344 14396 15350 14408
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 15344 14368 15761 14396
rect 15344 14356 15350 14368
rect 15749 14365 15761 14368
rect 15795 14365 15807 14399
rect 15749 14359 15807 14365
rect 14274 14328 14280 14340
rect 12667 14300 12940 14328
rect 14235 14300 14280 14328
rect 12667 14297 12679 14300
rect 12621 14291 12679 14297
rect 14274 14288 14280 14300
rect 14332 14288 14338 14340
rect 15194 14328 15200 14340
rect 14384 14300 15200 14328
rect 7650 14260 7656 14272
rect 6052 14232 7411 14260
rect 7611 14232 7656 14260
rect 6052 14220 6058 14232
rect 7650 14220 7656 14232
rect 7708 14220 7714 14272
rect 9490 14220 9496 14272
rect 9548 14260 9554 14272
rect 12802 14260 12808 14272
rect 9548 14232 12808 14260
rect 9548 14220 9554 14232
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 12894 14220 12900 14272
rect 12952 14260 12958 14272
rect 14384 14260 14412 14300
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 15764 14328 15792 14359
rect 15838 14356 15844 14408
rect 15896 14396 15902 14408
rect 15896 14368 15941 14396
rect 15896 14356 15902 14368
rect 22462 14328 22468 14340
rect 15764 14300 22468 14328
rect 22462 14288 22468 14300
rect 22520 14288 22526 14340
rect 15286 14260 15292 14272
rect 12952 14232 14412 14260
rect 15247 14232 15292 14260
rect 12952 14220 12958 14232
rect 15286 14220 15292 14232
rect 15344 14220 15350 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 1397 14059 1455 14065
rect 1397 14025 1409 14059
rect 1443 14056 1455 14059
rect 3418 14056 3424 14068
rect 1443 14028 3424 14056
rect 1443 14025 1455 14028
rect 1397 14019 1455 14025
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 5994 14056 6000 14068
rect 4172 14028 6000 14056
rect 1670 13880 1676 13932
rect 1728 13920 1734 13932
rect 1857 13923 1915 13929
rect 1857 13920 1869 13923
rect 1728 13892 1869 13920
rect 1728 13880 1734 13892
rect 1857 13889 1869 13892
rect 1903 13889 1915 13923
rect 2038 13920 2044 13932
rect 1999 13892 2044 13920
rect 1857 13883 1915 13889
rect 1118 13812 1124 13864
rect 1176 13852 1182 13864
rect 1765 13855 1823 13861
rect 1765 13852 1777 13855
rect 1176 13824 1777 13852
rect 1176 13812 1182 13824
rect 1765 13821 1777 13824
rect 1811 13821 1823 13855
rect 1872 13852 1900 13883
rect 2038 13880 2044 13892
rect 2096 13880 2102 13932
rect 2130 13880 2136 13932
rect 2188 13920 2194 13932
rect 2409 13923 2467 13929
rect 2409 13920 2421 13923
rect 2188 13892 2421 13920
rect 2188 13880 2194 13892
rect 2409 13889 2421 13892
rect 2455 13889 2467 13923
rect 2409 13883 2467 13889
rect 4172 13852 4200 14028
rect 5994 14016 6000 14028
rect 6052 14016 6058 14068
rect 7101 14059 7159 14065
rect 7101 14056 7113 14059
rect 6840 14028 7113 14056
rect 6840 13988 6868 14028
rect 7101 14025 7113 14028
rect 7147 14025 7159 14059
rect 7101 14019 7159 14025
rect 7745 14059 7803 14065
rect 7745 14025 7757 14059
rect 7791 14056 7803 14059
rect 8938 14056 8944 14068
rect 7791 14028 8944 14056
rect 7791 14025 7803 14028
rect 7745 14019 7803 14025
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 9030 14016 9036 14068
rect 9088 14056 9094 14068
rect 9861 14059 9919 14065
rect 9861 14056 9873 14059
rect 9088 14028 9873 14056
rect 9088 14016 9094 14028
rect 9861 14025 9873 14028
rect 9907 14025 9919 14059
rect 9861 14019 9919 14025
rect 10778 14016 10784 14068
rect 10836 14056 10842 14068
rect 10873 14059 10931 14065
rect 10873 14056 10885 14059
rect 10836 14028 10885 14056
rect 10836 14016 10842 14028
rect 10873 14025 10885 14028
rect 10919 14025 10931 14059
rect 12526 14056 12532 14068
rect 12487 14028 12532 14056
rect 10873 14019 10931 14025
rect 12526 14016 12532 14028
rect 12584 14016 12590 14068
rect 13357 14059 13415 14065
rect 13357 14025 13369 14059
rect 13403 14056 13415 14059
rect 14274 14056 14280 14068
rect 13403 14028 14280 14056
rect 13403 14025 13415 14028
rect 13357 14019 13415 14025
rect 14274 14016 14280 14028
rect 14332 14016 14338 14068
rect 6288 13960 6868 13988
rect 4246 13880 4252 13932
rect 4304 13920 4310 13932
rect 4304 13892 4568 13920
rect 4304 13880 4310 13892
rect 1872 13824 4200 13852
rect 4433 13855 4491 13861
rect 1765 13815 1823 13821
rect 4433 13821 4445 13855
rect 4479 13821 4491 13855
rect 4540 13852 4568 13892
rect 4689 13855 4747 13861
rect 4689 13852 4701 13855
rect 4540 13824 4701 13852
rect 4433 13815 4491 13821
rect 4689 13821 4701 13824
rect 4735 13821 4747 13855
rect 4689 13815 4747 13821
rect 2682 13793 2688 13796
rect 2665 13787 2688 13793
rect 2665 13753 2677 13787
rect 2740 13784 2746 13796
rect 3602 13784 3608 13796
rect 2740 13756 3608 13784
rect 2665 13747 2688 13753
rect 2682 13744 2688 13747
rect 2740 13744 2746 13756
rect 3602 13744 3608 13756
rect 3660 13744 3666 13796
rect 4246 13744 4252 13796
rect 4304 13784 4310 13796
rect 4448 13784 4476 13815
rect 6178 13812 6184 13864
rect 6236 13852 6242 13864
rect 6288 13861 6316 13960
rect 6914 13948 6920 14000
rect 6972 13988 6978 14000
rect 8018 13988 8024 14000
rect 6972 13960 8024 13988
rect 6972 13948 6978 13960
rect 8018 13948 8024 13960
rect 8076 13948 8082 14000
rect 8294 13948 8300 14000
rect 8352 13988 8358 14000
rect 8757 13991 8815 13997
rect 8757 13988 8769 13991
rect 8352 13960 8769 13988
rect 8352 13948 8358 13960
rect 8757 13957 8769 13960
rect 8803 13957 8815 13991
rect 15286 13988 15292 14000
rect 8757 13951 8815 13957
rect 10336 13960 15292 13988
rect 8036 13920 8064 13948
rect 8389 13923 8447 13929
rect 8036 13892 8340 13920
rect 6273 13855 6331 13861
rect 6273 13852 6285 13855
rect 6236 13824 6285 13852
rect 6236 13812 6242 13824
rect 6273 13821 6285 13824
rect 6319 13821 6331 13855
rect 7282 13852 7288 13864
rect 7243 13824 7288 13852
rect 6273 13815 6331 13821
rect 7282 13812 7288 13824
rect 7340 13812 7346 13864
rect 7650 13812 7656 13864
rect 7708 13852 7714 13864
rect 8113 13855 8171 13861
rect 8113 13852 8125 13855
rect 7708 13824 8125 13852
rect 7708 13812 7714 13824
rect 8113 13821 8125 13824
rect 8159 13821 8171 13855
rect 8312 13852 8340 13892
rect 8389 13889 8401 13923
rect 8435 13920 8447 13923
rect 8478 13920 8484 13932
rect 8435 13892 8484 13920
rect 8435 13889 8447 13892
rect 8389 13883 8447 13889
rect 8478 13880 8484 13892
rect 8536 13880 8542 13932
rect 9306 13920 9312 13932
rect 9267 13892 9312 13920
rect 9306 13880 9312 13892
rect 9364 13880 9370 13932
rect 10336 13929 10364 13960
rect 15286 13948 15292 13960
rect 15344 13948 15350 14000
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13889 10379 13923
rect 10502 13920 10508 13932
rect 10463 13892 10508 13920
rect 10321 13883 10379 13889
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 10888 13892 11468 13920
rect 10888 13852 10916 13892
rect 8312 13824 10916 13852
rect 8113 13815 8171 13821
rect 10962 13812 10968 13864
rect 11020 13852 11026 13864
rect 11333 13855 11391 13861
rect 11333 13852 11345 13855
rect 11020 13824 11345 13852
rect 11020 13812 11026 13824
rect 11333 13821 11345 13824
rect 11379 13821 11391 13855
rect 11440 13852 11468 13892
rect 11514 13880 11520 13932
rect 11572 13920 11578 13932
rect 11572 13892 11617 13920
rect 11572 13880 11578 13892
rect 12802 13880 12808 13932
rect 12860 13920 12866 13932
rect 13173 13923 13231 13929
rect 12860 13892 13032 13920
rect 12860 13880 12866 13892
rect 12894 13852 12900 13864
rect 11440 13824 12900 13852
rect 11333 13815 11391 13821
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 13004 13852 13032 13892
rect 13173 13889 13185 13923
rect 13219 13920 13231 13923
rect 13357 13923 13415 13929
rect 13357 13920 13369 13923
rect 13219 13892 13369 13920
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 13357 13889 13369 13892
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 13446 13880 13452 13932
rect 13504 13920 13510 13932
rect 14093 13923 14151 13929
rect 14093 13920 14105 13923
rect 13504 13892 14105 13920
rect 13504 13880 13510 13892
rect 14093 13889 14105 13892
rect 14139 13889 14151 13923
rect 15010 13920 15016 13932
rect 14971 13892 15016 13920
rect 14093 13883 14151 13889
rect 15010 13880 15016 13892
rect 15068 13880 15074 13932
rect 15194 13920 15200 13932
rect 15107 13892 15200 13920
rect 15194 13880 15200 13892
rect 15252 13920 15258 13932
rect 15838 13920 15844 13932
rect 15252 13892 15844 13920
rect 15252 13880 15258 13892
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 13906 13852 13912 13864
rect 13004 13824 13912 13852
rect 13906 13812 13912 13824
rect 13964 13812 13970 13864
rect 4304 13756 4476 13784
rect 8205 13787 8263 13793
rect 4304 13744 4310 13756
rect 8205 13753 8217 13787
rect 8251 13784 8263 13787
rect 8294 13784 8300 13796
rect 8251 13756 8300 13784
rect 8251 13753 8263 13756
rect 8205 13747 8263 13753
rect 8294 13744 8300 13756
rect 8352 13744 8358 13796
rect 10134 13784 10140 13796
rect 8404 13756 10140 13784
rect 2958 13676 2964 13728
rect 3016 13716 3022 13728
rect 3694 13716 3700 13728
rect 3016 13688 3700 13716
rect 3016 13676 3022 13688
rect 3694 13676 3700 13688
rect 3752 13676 3758 13728
rect 3786 13676 3792 13728
rect 3844 13716 3850 13728
rect 5810 13716 5816 13728
rect 3844 13688 3889 13716
rect 5771 13688 5816 13716
rect 3844 13676 3850 13688
rect 5810 13676 5816 13688
rect 5868 13676 5874 13728
rect 5994 13676 6000 13728
rect 6052 13716 6058 13728
rect 6089 13719 6147 13725
rect 6089 13716 6101 13719
rect 6052 13688 6101 13716
rect 6052 13676 6058 13688
rect 6089 13685 6101 13688
rect 6135 13685 6147 13719
rect 6089 13679 6147 13685
rect 6546 13676 6552 13728
rect 6604 13716 6610 13728
rect 8404 13716 8432 13756
rect 10134 13744 10140 13756
rect 10192 13744 10198 13796
rect 10229 13787 10287 13793
rect 10229 13753 10241 13787
rect 10275 13784 10287 13787
rect 10275 13756 14596 13784
rect 10275 13753 10287 13756
rect 10229 13747 10287 13753
rect 6604 13688 8432 13716
rect 6604 13676 6610 13688
rect 8754 13676 8760 13728
rect 8812 13716 8818 13728
rect 9122 13716 9128 13728
rect 8812 13688 9128 13716
rect 8812 13676 8818 13688
rect 9122 13676 9128 13688
rect 9180 13676 9186 13728
rect 9214 13676 9220 13728
rect 9272 13716 9278 13728
rect 9272 13688 9317 13716
rect 9272 13676 9278 13688
rect 9674 13676 9680 13728
rect 9732 13716 9738 13728
rect 10870 13716 10876 13728
rect 9732 13688 10876 13716
rect 9732 13676 9738 13688
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 11238 13716 11244 13728
rect 11199 13688 11244 13716
rect 11238 13676 11244 13688
rect 11296 13676 11302 13728
rect 12894 13716 12900 13728
rect 12855 13688 12900 13716
rect 12894 13676 12900 13688
rect 12952 13676 12958 13728
rect 12989 13719 13047 13725
rect 12989 13685 13001 13719
rect 13035 13716 13047 13719
rect 13541 13719 13599 13725
rect 13541 13716 13553 13719
rect 13035 13688 13553 13716
rect 13035 13685 13047 13688
rect 12989 13679 13047 13685
rect 13541 13685 13553 13688
rect 13587 13685 13599 13719
rect 13541 13679 13599 13685
rect 13722 13676 13728 13728
rect 13780 13716 13786 13728
rect 14001 13719 14059 13725
rect 14001 13716 14013 13719
rect 13780 13688 14013 13716
rect 13780 13676 13786 13688
rect 14001 13685 14013 13688
rect 14047 13716 14059 13719
rect 14366 13716 14372 13728
rect 14047 13688 14372 13716
rect 14047 13685 14059 13688
rect 14001 13679 14059 13685
rect 14366 13676 14372 13688
rect 14424 13676 14430 13728
rect 14568 13725 14596 13756
rect 14642 13744 14648 13796
rect 14700 13784 14706 13796
rect 14921 13787 14979 13793
rect 14921 13784 14933 13787
rect 14700 13756 14933 13784
rect 14700 13744 14706 13756
rect 14921 13753 14933 13756
rect 14967 13753 14979 13787
rect 14921 13747 14979 13753
rect 14553 13719 14611 13725
rect 14553 13685 14565 13719
rect 14599 13685 14611 13719
rect 14553 13679 14611 13685
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 2961 13515 3019 13521
rect 2961 13481 2973 13515
rect 3007 13512 3019 13515
rect 4525 13515 4583 13521
rect 4525 13512 4537 13515
rect 3007 13484 4537 13512
rect 3007 13481 3019 13484
rect 2961 13475 3019 13481
rect 4525 13481 4537 13484
rect 4571 13481 4583 13515
rect 4525 13475 4583 13481
rect 4706 13472 4712 13524
rect 4764 13512 4770 13524
rect 9214 13512 9220 13524
rect 4764 13484 9220 13512
rect 4764 13472 4770 13484
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 9309 13515 9367 13521
rect 9309 13481 9321 13515
rect 9355 13481 9367 13515
rect 13170 13512 13176 13524
rect 9309 13475 9367 13481
rect 10060 13484 13176 13512
rect 2222 13444 2228 13456
rect 1412 13416 2228 13444
rect 1412 13385 1440 13416
rect 2222 13404 2228 13416
rect 2280 13404 2286 13456
rect 3418 13444 3424 13456
rect 3379 13416 3424 13444
rect 3418 13404 3424 13416
rect 3476 13404 3482 13456
rect 4154 13404 4160 13456
rect 4212 13444 4218 13456
rect 4433 13447 4491 13453
rect 4433 13444 4445 13447
rect 4212 13416 4445 13444
rect 4212 13404 4218 13416
rect 4433 13413 4445 13416
rect 4479 13413 4491 13447
rect 5626 13444 5632 13456
rect 5587 13416 5632 13444
rect 4433 13407 4491 13413
rect 5626 13404 5632 13416
rect 5684 13404 5690 13456
rect 5810 13404 5816 13456
rect 5868 13444 5874 13456
rect 6426 13447 6484 13453
rect 6426 13444 6438 13447
rect 5868 13416 6438 13444
rect 5868 13404 5874 13416
rect 6426 13413 6438 13416
rect 6472 13413 6484 13447
rect 9324 13444 9352 13475
rect 9582 13444 9588 13456
rect 6426 13407 6484 13413
rect 6564 13416 8892 13444
rect 9324 13416 9588 13444
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13345 1455 13379
rect 1397 13339 1455 13345
rect 1578 13336 1584 13388
rect 1636 13376 1642 13388
rect 2317 13379 2375 13385
rect 2317 13376 2329 13379
rect 1636 13348 2329 13376
rect 1636 13336 1642 13348
rect 2317 13345 2329 13348
rect 2363 13345 2375 13379
rect 2317 13339 2375 13345
rect 3050 13336 3056 13388
rect 3108 13376 3114 13388
rect 3329 13379 3387 13385
rect 3329 13376 3341 13379
rect 3108 13348 3341 13376
rect 3108 13336 3114 13348
rect 3329 13345 3341 13348
rect 3375 13345 3387 13379
rect 5534 13376 5540 13388
rect 3329 13339 3387 13345
rect 3436 13348 4732 13376
rect 5495 13348 5540 13376
rect 3436 13320 3464 13348
rect 2409 13311 2467 13317
rect 2409 13277 2421 13311
rect 2455 13308 2467 13311
rect 2498 13308 2504 13320
rect 2455 13280 2504 13308
rect 2455 13277 2467 13280
rect 2409 13271 2467 13277
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 2593 13311 2651 13317
rect 2593 13277 2605 13311
rect 2639 13277 2651 13311
rect 2593 13271 2651 13277
rect 2608 13240 2636 13271
rect 3418 13268 3424 13320
rect 3476 13268 3482 13320
rect 3602 13308 3608 13320
rect 3563 13280 3608 13308
rect 3602 13268 3608 13280
rect 3660 13268 3666 13320
rect 3786 13268 3792 13320
rect 3844 13308 3850 13320
rect 4617 13311 4675 13317
rect 4617 13308 4629 13311
rect 3844 13280 4629 13308
rect 3844 13268 3850 13280
rect 4617 13277 4629 13280
rect 4663 13277 4675 13311
rect 4704 13308 4732 13348
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 6564 13376 6592 13416
rect 5644 13348 6592 13376
rect 8196 13379 8254 13385
rect 5644 13308 5672 13348
rect 8196 13345 8208 13379
rect 8242 13376 8254 13379
rect 8478 13376 8484 13388
rect 8242 13348 8484 13376
rect 8242 13345 8254 13348
rect 8196 13339 8254 13345
rect 8478 13336 8484 13348
rect 8536 13376 8542 13388
rect 8754 13376 8760 13388
rect 8536 13348 8760 13376
rect 8536 13336 8542 13348
rect 8754 13336 8760 13348
rect 8812 13336 8818 13388
rect 8864 13376 8892 13416
rect 9582 13404 9588 13416
rect 9640 13444 9646 13456
rect 9922 13447 9980 13453
rect 9922 13444 9934 13447
rect 9640 13416 9934 13444
rect 9640 13404 9646 13416
rect 9922 13413 9934 13416
rect 9968 13413 9980 13447
rect 9922 13407 9980 13413
rect 10060 13376 10088 13484
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 13446 13512 13452 13524
rect 13407 13484 13452 13512
rect 13446 13472 13452 13484
rect 13504 13472 13510 13524
rect 14090 13472 14096 13524
rect 14148 13512 14154 13524
rect 14185 13515 14243 13521
rect 14185 13512 14197 13515
rect 14148 13484 14197 13512
rect 14148 13472 14154 13484
rect 14185 13481 14197 13484
rect 14231 13481 14243 13515
rect 14185 13475 14243 13481
rect 14366 13472 14372 13524
rect 14424 13512 14430 13524
rect 15654 13512 15660 13524
rect 14424 13484 15660 13512
rect 14424 13472 14430 13484
rect 15654 13472 15660 13484
rect 15712 13472 15718 13524
rect 20533 13515 20591 13521
rect 20533 13481 20545 13515
rect 20579 13481 20591 13515
rect 20533 13475 20591 13481
rect 10134 13404 10140 13456
rect 10192 13444 10198 13456
rect 20548 13444 20576 13475
rect 10192 13416 20576 13444
rect 10192 13404 10198 13416
rect 8864 13348 10088 13376
rect 11054 13336 11060 13388
rect 11112 13376 11118 13388
rect 11333 13379 11391 13385
rect 11333 13376 11345 13379
rect 11112 13348 11345 13376
rect 11112 13336 11118 13348
rect 11333 13345 11345 13348
rect 11379 13345 11391 13379
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 11333 13339 11391 13345
rect 11440 13348 12081 13376
rect 4704 13280 5672 13308
rect 5813 13311 5871 13317
rect 4617 13271 4675 13277
rect 5813 13277 5825 13311
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 3804 13240 3832 13268
rect 4062 13240 4068 13252
rect 2608 13212 3832 13240
rect 4023 13212 4068 13240
rect 4062 13200 4068 13212
rect 4120 13200 4126 13252
rect 5258 13200 5264 13252
rect 5316 13240 5322 13252
rect 5828 13240 5856 13271
rect 5994 13268 6000 13320
rect 6052 13308 6058 13320
rect 6181 13311 6239 13317
rect 6181 13308 6193 13311
rect 6052 13280 6193 13308
rect 6052 13268 6058 13280
rect 6181 13277 6193 13280
rect 6227 13277 6239 13311
rect 6181 13271 6239 13277
rect 7374 13268 7380 13320
rect 7432 13308 7438 13320
rect 7742 13308 7748 13320
rect 7432 13280 7748 13308
rect 7432 13268 7438 13280
rect 7742 13268 7748 13280
rect 7800 13308 7806 13320
rect 7929 13311 7987 13317
rect 7929 13308 7941 13311
rect 7800 13280 7941 13308
rect 7800 13268 7806 13280
rect 7929 13277 7941 13280
rect 7975 13277 7987 13311
rect 9674 13308 9680 13320
rect 9635 13280 9680 13308
rect 7929 13271 7987 13277
rect 9674 13268 9680 13280
rect 9732 13268 9738 13320
rect 10870 13268 10876 13320
rect 10928 13308 10934 13320
rect 11440 13308 11468 13348
rect 12069 13345 12081 13348
rect 12115 13345 12127 13379
rect 12069 13339 12127 13345
rect 12158 13336 12164 13388
rect 12216 13376 12222 13388
rect 12325 13379 12383 13385
rect 12325 13376 12337 13379
rect 12216 13348 12337 13376
rect 12216 13336 12222 13348
rect 12325 13345 12337 13348
rect 12371 13345 12383 13379
rect 12325 13339 12383 13345
rect 14093 13379 14151 13385
rect 14093 13345 14105 13379
rect 14139 13376 14151 13379
rect 15286 13376 15292 13388
rect 14139 13348 15292 13376
rect 14139 13345 14151 13348
rect 14093 13339 14151 13345
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 19426 13385 19432 13388
rect 19420 13339 19432 13385
rect 19484 13376 19490 13388
rect 19484 13348 19520 13376
rect 19426 13336 19432 13339
rect 19484 13336 19490 13348
rect 11606 13308 11612 13320
rect 10928 13280 11468 13308
rect 11567 13280 11612 13308
rect 10928 13268 10934 13280
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 14366 13308 14372 13320
rect 14327 13280 14372 13308
rect 14366 13268 14372 13280
rect 14424 13268 14430 13320
rect 19150 13308 19156 13320
rect 19111 13280 19156 13308
rect 19150 13268 19156 13280
rect 19208 13268 19214 13320
rect 11238 13240 11244 13252
rect 5316 13212 6224 13240
rect 5316 13200 5322 13212
rect 1949 13175 2007 13181
rect 1949 13141 1961 13175
rect 1995 13172 2007 13175
rect 3510 13172 3516 13184
rect 1995 13144 3516 13172
rect 1995 13141 2007 13144
rect 1949 13135 2007 13141
rect 3510 13132 3516 13144
rect 3568 13132 3574 13184
rect 3970 13132 3976 13184
rect 4028 13172 4034 13184
rect 5074 13172 5080 13184
rect 4028 13144 5080 13172
rect 4028 13132 4034 13144
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 5169 13175 5227 13181
rect 5169 13141 5181 13175
rect 5215 13172 5227 13175
rect 6086 13172 6092 13184
rect 5215 13144 6092 13172
rect 5215 13141 5227 13144
rect 5169 13135 5227 13141
rect 6086 13132 6092 13144
rect 6144 13132 6150 13184
rect 6196 13172 6224 13212
rect 10980 13212 11244 13240
rect 7098 13172 7104 13184
rect 6196 13144 7104 13172
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 7561 13175 7619 13181
rect 7561 13141 7573 13175
rect 7607 13172 7619 13175
rect 7650 13172 7656 13184
rect 7607 13144 7656 13172
rect 7607 13141 7619 13144
rect 7561 13135 7619 13141
rect 7650 13132 7656 13144
rect 7708 13172 7714 13184
rect 8202 13172 8208 13184
rect 7708 13144 8208 13172
rect 7708 13132 7714 13144
rect 8202 13132 8208 13144
rect 8260 13132 8266 13184
rect 8294 13132 8300 13184
rect 8352 13172 8358 13184
rect 10980 13172 11008 13212
rect 11238 13200 11244 13212
rect 11296 13240 11302 13252
rect 12066 13240 12072 13252
rect 11296 13212 12072 13240
rect 11296 13200 11302 13212
rect 12066 13200 12072 13212
rect 12124 13200 12130 13252
rect 14090 13200 14096 13252
rect 14148 13240 14154 13252
rect 14458 13240 14464 13252
rect 14148 13212 14464 13240
rect 14148 13200 14154 13212
rect 14458 13200 14464 13212
rect 14516 13200 14522 13252
rect 8352 13144 11008 13172
rect 11057 13175 11115 13181
rect 8352 13132 8358 13144
rect 11057 13141 11069 13175
rect 11103 13172 11115 13175
rect 11606 13172 11612 13184
rect 11103 13144 11612 13172
rect 11103 13141 11115 13144
rect 11057 13135 11115 13141
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 13725 13175 13783 13181
rect 13725 13141 13737 13175
rect 13771 13172 13783 13175
rect 14274 13172 14280 13184
rect 13771 13144 14280 13172
rect 13771 13141 13783 13144
rect 13725 13135 13783 13141
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 2406 12968 2412 12980
rect 2367 12940 2412 12968
rect 2406 12928 2412 12940
rect 2464 12928 2470 12980
rect 3605 12971 3663 12977
rect 3605 12937 3617 12971
rect 3651 12968 3663 12971
rect 3694 12968 3700 12980
rect 3651 12940 3700 12968
rect 3651 12937 3663 12940
rect 3605 12931 3663 12937
rect 3694 12928 3700 12940
rect 3752 12928 3758 12980
rect 3970 12928 3976 12980
rect 4028 12968 4034 12980
rect 10870 12968 10876 12980
rect 4028 12940 10876 12968
rect 4028 12928 4034 12940
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 12069 12971 12127 12977
rect 12069 12937 12081 12971
rect 12115 12968 12127 12971
rect 12158 12968 12164 12980
rect 12115 12940 12164 12968
rect 12115 12937 12127 12940
rect 12069 12931 12127 12937
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 12618 12928 12624 12980
rect 12676 12968 12682 12980
rect 12897 12971 12955 12977
rect 12897 12968 12909 12971
rect 12676 12940 12909 12968
rect 12676 12928 12682 12940
rect 12897 12937 12909 12940
rect 12943 12937 12955 12971
rect 12897 12931 12955 12937
rect 12986 12928 12992 12980
rect 13044 12968 13050 12980
rect 13538 12968 13544 12980
rect 13044 12940 13544 12968
rect 13044 12928 13050 12940
rect 2682 12900 2688 12912
rect 2240 12872 2688 12900
rect 2240 12841 2268 12872
rect 2682 12860 2688 12872
rect 2740 12860 2746 12912
rect 3510 12860 3516 12912
rect 3568 12900 3574 12912
rect 8754 12900 8760 12912
rect 3568 12872 6868 12900
rect 8667 12872 8760 12900
rect 3568 12860 3574 12872
rect 2225 12835 2283 12841
rect 2225 12801 2237 12835
rect 2271 12801 2283 12835
rect 2958 12832 2964 12844
rect 2919 12804 2964 12832
rect 2225 12795 2283 12801
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 3234 12792 3240 12844
rect 3292 12832 3298 12844
rect 3292 12804 3464 12832
rect 3292 12792 3298 12804
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12764 2007 12767
rect 2682 12764 2688 12776
rect 1995 12736 2688 12764
rect 1995 12733 2007 12736
rect 1949 12727 2007 12733
rect 2682 12724 2688 12736
rect 2740 12724 2746 12776
rect 3436 12764 3464 12804
rect 4062 12792 4068 12844
rect 4120 12832 4126 12844
rect 4157 12835 4215 12841
rect 4157 12832 4169 12835
rect 4120 12804 4169 12832
rect 4120 12792 4126 12804
rect 4157 12801 4169 12804
rect 4203 12801 4215 12835
rect 4157 12795 4215 12801
rect 5077 12835 5135 12841
rect 5077 12801 5089 12835
rect 5123 12832 5135 12835
rect 5166 12832 5172 12844
rect 5123 12804 5172 12832
rect 5123 12801 5135 12804
rect 5077 12795 5135 12801
rect 5166 12792 5172 12804
rect 5224 12792 5230 12844
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12832 5319 12835
rect 5810 12832 5816 12844
rect 5307 12804 5816 12832
rect 5307 12801 5319 12804
rect 5261 12795 5319 12801
rect 5810 12792 5816 12804
rect 5868 12792 5874 12844
rect 6178 12832 6184 12844
rect 6139 12804 6184 12832
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 6086 12764 6092 12776
rect 3436 12736 5764 12764
rect 6047 12736 6092 12764
rect 2777 12699 2835 12705
rect 2777 12665 2789 12699
rect 2823 12696 2835 12699
rect 3234 12696 3240 12708
rect 2823 12668 3240 12696
rect 2823 12665 2835 12668
rect 2777 12659 2835 12665
rect 3234 12656 3240 12668
rect 3292 12656 3298 12708
rect 3878 12656 3884 12708
rect 3936 12696 3942 12708
rect 4065 12699 4123 12705
rect 4065 12696 4077 12699
rect 3936 12668 4077 12696
rect 3936 12656 3942 12668
rect 4065 12665 4077 12668
rect 4111 12665 4123 12699
rect 4798 12696 4804 12708
rect 4065 12659 4123 12665
rect 4325 12668 4804 12696
rect 2038 12628 2044 12640
rect 1999 12600 2044 12628
rect 2038 12588 2044 12600
rect 2096 12588 2102 12640
rect 2869 12631 2927 12637
rect 2869 12597 2881 12631
rect 2915 12628 2927 12631
rect 3418 12628 3424 12640
rect 2915 12600 3424 12628
rect 2915 12597 2927 12600
rect 2869 12591 2927 12597
rect 3418 12588 3424 12600
rect 3476 12588 3482 12640
rect 3513 12631 3571 12637
rect 3513 12597 3525 12631
rect 3559 12628 3571 12631
rect 3973 12631 4031 12637
rect 3973 12628 3985 12631
rect 3559 12600 3985 12628
rect 3559 12597 3571 12600
rect 3513 12591 3571 12597
rect 3973 12597 3985 12600
rect 4019 12628 4031 12631
rect 4325 12628 4353 12668
rect 4798 12656 4804 12668
rect 4856 12656 4862 12708
rect 4985 12699 5043 12705
rect 4985 12665 4997 12699
rect 5031 12696 5043 12699
rect 5074 12696 5080 12708
rect 5031 12668 5080 12696
rect 5031 12665 5043 12668
rect 4985 12659 5043 12665
rect 5074 12656 5080 12668
rect 5132 12656 5138 12708
rect 4019 12600 4353 12628
rect 4617 12631 4675 12637
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 4617 12597 4629 12631
rect 4663 12628 4675 12631
rect 4706 12628 4712 12640
rect 4663 12600 4712 12628
rect 4663 12597 4675 12600
rect 4617 12591 4675 12597
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 5626 12628 5632 12640
rect 5587 12600 5632 12628
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 5736 12628 5764 12736
rect 6086 12724 6092 12736
rect 6144 12724 6150 12776
rect 6840 12773 6868 12872
rect 8754 12860 8760 12872
rect 8812 12900 8818 12912
rect 9122 12900 9128 12912
rect 8812 12872 9128 12900
rect 8812 12860 8818 12872
rect 9122 12860 9128 12872
rect 9180 12860 9186 12912
rect 10410 12900 10416 12912
rect 9416 12872 10416 12900
rect 7374 12832 7380 12844
rect 7335 12804 7380 12832
rect 7374 12792 7380 12804
rect 7432 12792 7438 12844
rect 8849 12835 8907 12841
rect 8849 12801 8861 12835
rect 8895 12832 8907 12835
rect 9416 12832 9444 12872
rect 10410 12860 10416 12872
rect 10468 12860 10474 12912
rect 9582 12832 9588 12844
rect 8895 12804 9444 12832
rect 9543 12804 9588 12832
rect 8895 12801 8907 12804
rect 8849 12795 8907 12801
rect 9582 12792 9588 12804
rect 9640 12792 9646 12844
rect 13280 12841 13308 12940
rect 13538 12928 13544 12940
rect 13596 12968 13602 12980
rect 19150 12968 19156 12980
rect 13596 12940 19156 12968
rect 13596 12928 13602 12940
rect 19150 12928 19156 12940
rect 19208 12928 19214 12980
rect 13265 12835 13323 12841
rect 13265 12801 13277 12835
rect 13311 12801 13323 12835
rect 17310 12832 17316 12844
rect 17271 12804 17316 12832
rect 13265 12795 13323 12801
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 7650 12773 7656 12776
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12733 6883 12767
rect 7644 12764 7656 12773
rect 7611 12736 7656 12764
rect 6825 12727 6883 12733
rect 7644 12727 7656 12736
rect 7650 12724 7656 12727
rect 7708 12724 7714 12776
rect 8938 12724 8944 12776
rect 8996 12764 9002 12776
rect 9493 12767 9551 12773
rect 9493 12764 9505 12767
rect 8996 12736 9505 12764
rect 8996 12724 9002 12736
rect 9493 12733 9505 12736
rect 9539 12733 9551 12767
rect 9493 12727 9551 12733
rect 10410 12724 10416 12776
rect 10468 12764 10474 12776
rect 10689 12767 10747 12773
rect 10689 12764 10701 12767
rect 10468 12736 10701 12764
rect 10468 12724 10474 12736
rect 10689 12733 10701 12736
rect 10735 12764 10747 12767
rect 10778 12764 10784 12776
rect 10735 12736 10784 12764
rect 10735 12733 10747 12736
rect 10689 12727 10747 12733
rect 10778 12724 10784 12736
rect 10836 12724 10842 12776
rect 12986 12724 12992 12776
rect 13044 12764 13050 12776
rect 13081 12767 13139 12773
rect 13081 12764 13093 12767
rect 13044 12736 13093 12764
rect 13044 12724 13050 12736
rect 13081 12733 13093 12736
rect 13127 12733 13139 12767
rect 13081 12727 13139 12733
rect 13532 12767 13590 12773
rect 13532 12733 13544 12767
rect 13578 12764 13590 12767
rect 14366 12764 14372 12776
rect 13578 12736 14372 12764
rect 13578 12733 13590 12736
rect 13532 12727 13590 12733
rect 14366 12724 14372 12736
rect 14424 12724 14430 12776
rect 17034 12764 17040 12776
rect 16995 12736 17040 12764
rect 17034 12724 17040 12736
rect 17092 12724 17098 12776
rect 5997 12699 6055 12705
rect 5997 12665 6009 12699
rect 6043 12696 6055 12699
rect 10956 12699 11014 12705
rect 6043 12668 7604 12696
rect 6043 12665 6055 12668
rect 5997 12659 6055 12665
rect 7009 12631 7067 12637
rect 7009 12628 7021 12631
rect 5736 12600 7021 12628
rect 7009 12597 7021 12600
rect 7055 12597 7067 12631
rect 7576 12628 7604 12668
rect 10956 12665 10968 12699
rect 11002 12696 11014 12699
rect 11882 12696 11888 12708
rect 11002 12668 11888 12696
rect 11002 12665 11014 12668
rect 10956 12659 11014 12665
rect 11882 12656 11888 12668
rect 11940 12656 11946 12708
rect 14182 12696 14188 12708
rect 11992 12668 12756 12696
rect 8386 12628 8392 12640
rect 7576 12600 8392 12628
rect 7009 12591 7067 12597
rect 8386 12588 8392 12600
rect 8444 12588 8450 12640
rect 8849 12631 8907 12637
rect 8849 12597 8861 12631
rect 8895 12628 8907 12631
rect 9033 12631 9091 12637
rect 9033 12628 9045 12631
rect 8895 12600 9045 12628
rect 8895 12597 8907 12600
rect 8849 12591 8907 12597
rect 9033 12597 9045 12600
rect 9079 12597 9091 12631
rect 9398 12628 9404 12640
rect 9359 12600 9404 12628
rect 9033 12591 9091 12597
rect 9398 12588 9404 12600
rect 9456 12588 9462 12640
rect 9582 12588 9588 12640
rect 9640 12628 9646 12640
rect 11992 12628 12020 12668
rect 9640 12600 12020 12628
rect 12437 12631 12495 12637
rect 9640 12588 9646 12600
rect 12437 12597 12449 12631
rect 12483 12628 12495 12631
rect 12526 12628 12532 12640
rect 12483 12600 12532 12628
rect 12483 12597 12495 12600
rect 12437 12591 12495 12597
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 12728 12628 12756 12668
rect 13280 12668 14188 12696
rect 13280 12628 13308 12668
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 12728 12600 13308 12628
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 14645 12631 14703 12637
rect 14645 12628 14657 12631
rect 13964 12600 14657 12628
rect 13964 12588 13970 12600
rect 14645 12597 14657 12600
rect 14691 12597 14703 12631
rect 14645 12591 14703 12597
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 1489 12427 1547 12433
rect 1489 12393 1501 12427
rect 1535 12424 1547 12427
rect 1854 12424 1860 12436
rect 1535 12396 1860 12424
rect 1535 12393 1547 12396
rect 1489 12387 1547 12393
rect 1854 12384 1860 12396
rect 1912 12384 1918 12436
rect 2498 12424 2504 12436
rect 2459 12396 2504 12424
rect 2498 12384 2504 12396
rect 2556 12384 2562 12436
rect 2682 12384 2688 12436
rect 2740 12424 2746 12436
rect 3513 12427 3571 12433
rect 3513 12424 3525 12427
rect 2740 12396 3525 12424
rect 2740 12384 2746 12396
rect 3513 12393 3525 12396
rect 3559 12393 3571 12427
rect 3513 12387 3571 12393
rect 5626 12384 5632 12436
rect 5684 12424 5690 12436
rect 6549 12427 6607 12433
rect 6549 12424 6561 12427
rect 5684 12396 6561 12424
rect 5684 12384 5690 12396
rect 6549 12393 6561 12396
rect 6595 12393 6607 12427
rect 7558 12424 7564 12436
rect 7519 12396 7564 12424
rect 6549 12387 6607 12393
rect 7558 12384 7564 12396
rect 7616 12384 7622 12436
rect 7650 12384 7656 12436
rect 7708 12424 7714 12436
rect 8573 12427 8631 12433
rect 7708 12396 7753 12424
rect 7708 12384 7714 12396
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 9398 12424 9404 12436
rect 8619 12396 9404 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 9398 12384 9404 12396
rect 9456 12384 9462 12436
rect 9953 12427 10011 12433
rect 9953 12393 9965 12427
rect 9999 12393 10011 12427
rect 9953 12387 10011 12393
rect 10965 12427 11023 12433
rect 10965 12393 10977 12427
rect 11011 12424 11023 12427
rect 11054 12424 11060 12436
rect 11011 12396 11060 12424
rect 11011 12393 11023 12396
rect 10965 12387 11023 12393
rect 2869 12359 2927 12365
rect 2869 12325 2881 12359
rect 2915 12356 2927 12359
rect 2958 12356 2964 12368
rect 2915 12328 2964 12356
rect 2915 12325 2927 12328
rect 2869 12319 2927 12325
rect 2958 12316 2964 12328
rect 3016 12316 3022 12368
rect 4246 12316 4252 12368
rect 4304 12356 4310 12368
rect 5994 12356 6000 12368
rect 4304 12328 6000 12356
rect 4304 12316 4310 12328
rect 1854 12288 1860 12300
rect 1815 12260 1860 12288
rect 1854 12248 1860 12260
rect 1912 12248 1918 12300
rect 4448 12297 4476 12328
rect 5994 12316 6000 12328
rect 6052 12316 6058 12368
rect 6638 12316 6644 12368
rect 6696 12356 6702 12368
rect 7374 12356 7380 12368
rect 6696 12328 7380 12356
rect 6696 12316 6702 12328
rect 7374 12316 7380 12328
rect 7432 12316 7438 12368
rect 8386 12316 8392 12368
rect 8444 12356 8450 12368
rect 9968 12356 9996 12387
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 11333 12427 11391 12433
rect 11333 12393 11345 12427
rect 11379 12424 11391 12427
rect 11977 12427 12035 12433
rect 11977 12424 11989 12427
rect 11379 12396 11989 12424
rect 11379 12393 11391 12396
rect 11333 12387 11391 12393
rect 11977 12393 11989 12396
rect 12023 12393 12035 12427
rect 11977 12387 12035 12393
rect 12345 12427 12403 12433
rect 12345 12393 12357 12427
rect 12391 12424 12403 12427
rect 12526 12424 12532 12436
rect 12391 12396 12532 12424
rect 12391 12393 12403 12396
rect 12345 12387 12403 12393
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 12618 12384 12624 12436
rect 12676 12424 12682 12436
rect 12986 12424 12992 12436
rect 12676 12396 12992 12424
rect 12676 12384 12682 12396
rect 12986 12384 12992 12396
rect 13044 12384 13050 12436
rect 14921 12427 14979 12433
rect 14921 12424 14933 12427
rect 14016 12396 14933 12424
rect 14016 12368 14044 12396
rect 14921 12393 14933 12396
rect 14967 12393 14979 12427
rect 15286 12424 15292 12436
rect 15247 12396 15292 12424
rect 14921 12387 14979 12393
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 15470 12384 15476 12436
rect 15528 12424 15534 12436
rect 15749 12427 15807 12433
rect 15749 12424 15761 12427
rect 15528 12396 15761 12424
rect 15528 12384 15534 12396
rect 15749 12393 15761 12396
rect 15795 12424 15807 12427
rect 16298 12424 16304 12436
rect 15795 12396 16304 12424
rect 15795 12393 15807 12396
rect 15749 12387 15807 12393
rect 16298 12384 16304 12396
rect 16356 12384 16362 12436
rect 8444 12328 9996 12356
rect 10321 12359 10379 12365
rect 8444 12316 8450 12328
rect 10321 12325 10333 12359
rect 10367 12356 10379 12359
rect 11790 12356 11796 12368
rect 10367 12328 11796 12356
rect 10367 12325 10379 12328
rect 10321 12319 10379 12325
rect 11790 12316 11796 12328
rect 11848 12316 11854 12368
rect 12434 12316 12440 12368
rect 12492 12356 12498 12368
rect 13262 12356 13268 12368
rect 12492 12328 13268 12356
rect 12492 12316 12498 12328
rect 13262 12316 13268 12328
rect 13320 12316 13326 12368
rect 13808 12359 13866 12365
rect 13808 12325 13820 12359
rect 13854 12356 13866 12359
rect 13906 12356 13912 12368
rect 13854 12328 13912 12356
rect 13854 12325 13866 12328
rect 13808 12319 13866 12325
rect 13906 12316 13912 12328
rect 13964 12316 13970 12368
rect 13998 12316 14004 12368
rect 14056 12316 14062 12368
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12257 4491 12291
rect 4433 12251 4491 12257
rect 4700 12291 4758 12297
rect 4700 12257 4712 12291
rect 4746 12288 4758 12291
rect 5258 12288 5264 12300
rect 4746 12260 5264 12288
rect 4746 12257 4758 12260
rect 4700 12251 4758 12257
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 5626 12248 5632 12300
rect 5684 12288 5690 12300
rect 6457 12291 6515 12297
rect 6457 12288 6469 12291
rect 5684 12260 6469 12288
rect 5684 12248 5690 12260
rect 6457 12257 6469 12260
rect 6503 12257 6515 12291
rect 8938 12288 8944 12300
rect 8899 12260 8944 12288
rect 6457 12251 6515 12257
rect 8938 12248 8944 12260
rect 8996 12248 9002 12300
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12288 11483 12291
rect 11698 12288 11704 12300
rect 11471 12260 11704 12288
rect 11471 12257 11483 12260
rect 11425 12251 11483 12257
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 11882 12248 11888 12300
rect 11940 12288 11946 12300
rect 13538 12288 13544 12300
rect 11940 12260 12572 12288
rect 13499 12260 13544 12288
rect 11940 12248 11946 12260
rect 1946 12220 1952 12232
rect 1907 12192 1952 12220
rect 1946 12180 1952 12192
rect 2004 12180 2010 12232
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12189 2191 12223
rect 2133 12183 2191 12189
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12220 3019 12223
rect 3050 12220 3056 12232
rect 3007 12192 3056 12220
rect 3007 12189 3019 12192
rect 2961 12183 3019 12189
rect 2148 12084 2176 12183
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 3145 12223 3203 12229
rect 3145 12189 3157 12223
rect 3191 12220 3203 12223
rect 3602 12220 3608 12232
rect 3191 12192 3608 12220
rect 3191 12189 3203 12192
rect 3145 12183 3203 12189
rect 3602 12180 3608 12192
rect 3660 12180 3666 12232
rect 6638 12220 6644 12232
rect 6599 12192 6644 12220
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 7745 12223 7803 12229
rect 7745 12220 7757 12223
rect 7524 12192 7757 12220
rect 7524 12180 7530 12192
rect 7745 12189 7757 12192
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 8570 12180 8576 12232
rect 8628 12220 8634 12232
rect 9033 12223 9091 12229
rect 9033 12220 9045 12223
rect 8628 12192 9045 12220
rect 8628 12180 8634 12192
rect 9033 12189 9045 12192
rect 9079 12189 9091 12223
rect 9033 12183 9091 12189
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 10413 12223 10471 12229
rect 9180 12192 9225 12220
rect 9180 12180 9186 12192
rect 10413 12189 10425 12223
rect 10459 12189 10471 12223
rect 10594 12220 10600 12232
rect 10555 12192 10600 12220
rect 10413 12183 10471 12189
rect 6089 12155 6147 12161
rect 6089 12121 6101 12155
rect 6135 12152 6147 12155
rect 9858 12152 9864 12164
rect 6135 12124 9864 12152
rect 6135 12121 6147 12124
rect 6089 12115 6147 12121
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 9950 12112 9956 12164
rect 10008 12152 10014 12164
rect 10428 12152 10456 12183
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 11609 12223 11667 12229
rect 11609 12189 11621 12223
rect 11655 12220 11667 12223
rect 12158 12220 12164 12232
rect 11655 12192 12164 12220
rect 11655 12189 11667 12192
rect 11609 12183 11667 12189
rect 12158 12180 12164 12192
rect 12216 12180 12222 12232
rect 12544 12229 12572 12260
rect 13538 12248 13544 12260
rect 13596 12248 13602 12300
rect 15657 12291 15715 12297
rect 15657 12257 15669 12291
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 12529 12223 12587 12229
rect 12529 12189 12541 12223
rect 12575 12189 12587 12223
rect 12529 12183 12587 12189
rect 12986 12180 12992 12232
rect 13044 12220 13050 12232
rect 13556 12220 13584 12248
rect 13044 12192 13584 12220
rect 13044 12180 13050 12192
rect 14918 12180 14924 12232
rect 14976 12220 14982 12232
rect 15672 12220 15700 12251
rect 15838 12220 15844 12232
rect 14976 12192 15700 12220
rect 15799 12192 15844 12220
rect 14976 12180 14982 12192
rect 15838 12180 15844 12192
rect 15896 12180 15902 12232
rect 13538 12152 13544 12164
rect 10008 12124 13544 12152
rect 10008 12112 10014 12124
rect 13538 12112 13544 12124
rect 13596 12112 13602 12164
rect 5718 12084 5724 12096
rect 2148 12056 5724 12084
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 5813 12087 5871 12093
rect 5813 12053 5825 12087
rect 5859 12084 5871 12087
rect 6178 12084 6184 12096
rect 5859 12056 6184 12084
rect 5859 12053 5871 12056
rect 5813 12047 5871 12053
rect 6178 12044 6184 12056
rect 6236 12044 6242 12096
rect 7193 12087 7251 12093
rect 7193 12053 7205 12087
rect 7239 12084 7251 12087
rect 7742 12084 7748 12096
rect 7239 12056 7748 12084
rect 7239 12053 7251 12056
rect 7193 12047 7251 12053
rect 7742 12044 7748 12056
rect 7800 12044 7806 12096
rect 12894 12044 12900 12096
rect 12952 12084 12958 12096
rect 13170 12084 13176 12096
rect 12952 12056 13176 12084
rect 12952 12044 12958 12056
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 2774 11880 2780 11892
rect 1627 11852 2780 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 2774 11840 2780 11852
rect 2832 11840 2838 11892
rect 3970 11840 3976 11892
rect 4028 11880 4034 11892
rect 6181 11883 6239 11889
rect 4028 11852 6132 11880
rect 4028 11840 4034 11852
rect 6104 11812 6132 11852
rect 6181 11849 6193 11883
rect 6227 11880 6239 11883
rect 6638 11880 6644 11892
rect 6227 11852 6644 11880
rect 6227 11849 6239 11852
rect 6181 11843 6239 11849
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 8754 11880 8760 11892
rect 6840 11852 8760 11880
rect 6840 11812 6868 11852
rect 8754 11840 8760 11852
rect 8812 11840 8818 11892
rect 8938 11880 8944 11892
rect 8899 11852 8944 11880
rect 8938 11840 8944 11852
rect 8996 11840 9002 11892
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 9272 11852 11560 11880
rect 9272 11840 9278 11852
rect 10594 11812 10600 11824
rect 6104 11784 6868 11812
rect 7852 11784 10600 11812
rect 2406 11704 2412 11756
rect 2464 11744 2470 11756
rect 2501 11747 2559 11753
rect 2501 11744 2513 11747
rect 2464 11716 2513 11744
rect 2464 11704 2470 11716
rect 2501 11713 2513 11716
rect 2547 11713 2559 11747
rect 3602 11744 3608 11756
rect 3563 11716 3608 11744
rect 2501 11707 2559 11713
rect 3602 11704 3608 11716
rect 3660 11704 3666 11756
rect 5994 11704 6000 11756
rect 6052 11744 6058 11756
rect 6052 11716 6316 11744
rect 6052 11704 6058 11716
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11676 3479 11679
rect 3694 11676 3700 11688
rect 3467 11648 3700 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 3694 11636 3700 11648
rect 3752 11636 3758 11688
rect 3786 11636 3792 11688
rect 3844 11676 3850 11688
rect 3973 11679 4031 11685
rect 3973 11676 3985 11679
rect 3844 11648 3985 11676
rect 3844 11636 3850 11648
rect 3973 11645 3985 11648
rect 4019 11645 4031 11679
rect 4798 11676 4804 11688
rect 3973 11639 4031 11645
rect 4080 11648 4660 11676
rect 4759 11648 4804 11676
rect 2317 11611 2375 11617
rect 2317 11577 2329 11611
rect 2363 11608 2375 11611
rect 3050 11608 3056 11620
rect 2363 11580 3056 11608
rect 2363 11577 2375 11580
rect 2317 11571 2375 11577
rect 3050 11568 3056 11580
rect 3108 11568 3114 11620
rect 3878 11568 3884 11620
rect 3936 11608 3942 11620
rect 4080 11608 4108 11648
rect 4246 11608 4252 11620
rect 3936 11580 4108 11608
rect 4207 11580 4252 11608
rect 3936 11568 3942 11580
rect 4246 11568 4252 11580
rect 4304 11568 4310 11620
rect 4632 11608 4660 11648
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 5068 11679 5126 11685
rect 5068 11645 5080 11679
rect 5114 11676 5126 11679
rect 5534 11676 5540 11688
rect 5114 11648 5540 11676
rect 5114 11645 5126 11648
rect 5068 11639 5126 11645
rect 5534 11636 5540 11648
rect 5592 11676 5598 11688
rect 6178 11676 6184 11688
rect 5592 11648 6184 11676
rect 5592 11636 5598 11648
rect 6178 11636 6184 11648
rect 6236 11636 6242 11688
rect 6288 11676 6316 11716
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 6696 11716 6960 11744
rect 6696 11704 6702 11716
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6288 11648 6837 11676
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 6932 11676 6960 11716
rect 7081 11679 7139 11685
rect 7081 11676 7093 11679
rect 6932 11648 7093 11676
rect 6825 11639 6883 11645
rect 7081 11645 7093 11648
rect 7127 11645 7139 11679
rect 7852 11676 7880 11784
rect 10594 11772 10600 11784
rect 10652 11772 10658 11824
rect 11532 11812 11560 11852
rect 11882 11840 11888 11892
rect 11940 11880 11946 11892
rect 11977 11883 12035 11889
rect 11977 11880 11989 11883
rect 11940 11852 11989 11880
rect 11940 11840 11946 11852
rect 11977 11849 11989 11852
rect 12023 11849 12035 11883
rect 14366 11880 14372 11892
rect 14327 11852 14372 11880
rect 11977 11843 12035 11849
rect 14366 11840 14372 11852
rect 14424 11840 14430 11892
rect 12894 11812 12900 11824
rect 11532 11784 12900 11812
rect 12894 11772 12900 11784
rect 12952 11772 12958 11824
rect 7926 11704 7932 11756
rect 7984 11744 7990 11756
rect 7984 11716 9260 11744
rect 7984 11704 7990 11716
rect 8662 11676 8668 11688
rect 7081 11639 7139 11645
rect 7208 11648 7880 11676
rect 8623 11648 8668 11676
rect 7208 11620 7236 11648
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 9232 11676 9260 11716
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 9493 11747 9551 11753
rect 9493 11744 9505 11747
rect 9364 11716 9505 11744
rect 9364 11704 9370 11716
rect 9493 11713 9505 11716
rect 9539 11713 9551 11747
rect 12986 11744 12992 11756
rect 9493 11707 9551 11713
rect 9600 11716 10732 11744
rect 12947 11716 12992 11744
rect 9600 11676 9628 11716
rect 9232 11648 9628 11676
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 10410 11676 10416 11688
rect 9732 11648 10416 11676
rect 9732 11636 9738 11648
rect 10410 11636 10416 11648
rect 10468 11676 10474 11688
rect 10597 11679 10655 11685
rect 10597 11676 10609 11679
rect 10468 11648 10609 11676
rect 10468 11636 10474 11648
rect 10597 11645 10609 11648
rect 10643 11645 10655 11679
rect 10704 11676 10732 11716
rect 12986 11704 12992 11716
rect 13044 11704 13050 11756
rect 14384 11744 14412 11840
rect 15197 11747 15255 11753
rect 15197 11744 15209 11747
rect 14384 11716 15209 11744
rect 15197 11713 15209 11716
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 12158 11676 12164 11688
rect 10704 11648 12164 11676
rect 10597 11639 10655 11645
rect 11532 11620 11560 11648
rect 12158 11636 12164 11648
rect 12216 11636 12222 11688
rect 13256 11679 13314 11685
rect 13256 11645 13268 11679
rect 13302 11676 13314 11679
rect 13722 11676 13728 11688
rect 13302 11648 13728 11676
rect 13302 11645 13314 11648
rect 13256 11639 13314 11645
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 14182 11636 14188 11688
rect 14240 11676 14246 11688
rect 14918 11676 14924 11688
rect 14240 11648 14924 11676
rect 14240 11636 14246 11648
rect 14918 11636 14924 11648
rect 14976 11636 14982 11688
rect 6914 11608 6920 11620
rect 4632 11580 6920 11608
rect 6914 11568 6920 11580
rect 6972 11568 6978 11620
rect 7190 11568 7196 11620
rect 7248 11568 7254 11620
rect 7282 11568 7288 11620
rect 7340 11608 7346 11620
rect 9309 11611 9367 11617
rect 7340 11580 8524 11608
rect 7340 11568 7346 11580
rect 1486 11500 1492 11552
rect 1544 11540 1550 11552
rect 1949 11543 2007 11549
rect 1949 11540 1961 11543
rect 1544 11512 1961 11540
rect 1544 11500 1550 11512
rect 1949 11509 1961 11512
rect 1995 11509 2007 11543
rect 1949 11503 2007 11509
rect 2409 11543 2467 11549
rect 2409 11509 2421 11543
rect 2455 11540 2467 11543
rect 2961 11543 3019 11549
rect 2961 11540 2973 11543
rect 2455 11512 2973 11540
rect 2455 11509 2467 11512
rect 2409 11503 2467 11509
rect 2961 11509 2973 11512
rect 3007 11509 3019 11543
rect 3326 11540 3332 11552
rect 3287 11512 3332 11540
rect 2961 11503 3019 11509
rect 3326 11500 3332 11512
rect 3384 11500 3390 11552
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 8496 11549 8524 11580
rect 9309 11577 9321 11611
rect 9355 11608 9367 11611
rect 9953 11611 10011 11617
rect 9953 11608 9965 11611
rect 9355 11580 9965 11608
rect 9355 11577 9367 11580
rect 9309 11571 9367 11577
rect 9953 11577 9965 11580
rect 9999 11577 10011 11611
rect 9953 11571 10011 11577
rect 10864 11611 10922 11617
rect 10864 11577 10876 11611
rect 10910 11608 10922 11611
rect 11054 11608 11060 11620
rect 10910 11580 11060 11608
rect 10910 11577 10922 11580
rect 10864 11571 10922 11577
rect 11054 11568 11060 11580
rect 11112 11568 11118 11620
rect 11514 11568 11520 11620
rect 11572 11568 11578 11620
rect 12526 11568 12532 11620
rect 12584 11608 12590 11620
rect 13354 11608 13360 11620
rect 12584 11580 13360 11608
rect 12584 11568 12590 11580
rect 13354 11568 13360 11580
rect 13412 11568 13418 11620
rect 13740 11608 13768 11636
rect 14090 11608 14096 11620
rect 13740 11580 14096 11608
rect 14090 11568 14096 11580
rect 14148 11608 14154 11620
rect 15838 11608 15844 11620
rect 14148 11580 15844 11608
rect 14148 11568 14154 11580
rect 15838 11568 15844 11580
rect 15896 11568 15902 11620
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 7524 11512 8217 11540
rect 7524 11500 7530 11512
rect 8205 11509 8217 11512
rect 8251 11509 8263 11543
rect 8205 11503 8263 11509
rect 8481 11543 8539 11549
rect 8481 11509 8493 11543
rect 8527 11509 8539 11543
rect 8481 11503 8539 11509
rect 9214 11500 9220 11552
rect 9272 11540 9278 11552
rect 9401 11543 9459 11549
rect 9401 11540 9413 11543
rect 9272 11512 9413 11540
rect 9272 11500 9278 11512
rect 9401 11509 9413 11512
rect 9447 11509 9459 11543
rect 9401 11503 9459 11509
rect 10594 11500 10600 11552
rect 10652 11540 10658 11552
rect 14366 11540 14372 11552
rect 10652 11512 14372 11540
rect 10652 11500 10658 11512
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 14550 11500 14556 11552
rect 14608 11540 14614 11552
rect 14645 11543 14703 11549
rect 14645 11540 14657 11543
rect 14608 11512 14657 11540
rect 14608 11500 14614 11512
rect 14645 11509 14657 11512
rect 14691 11509 14703 11543
rect 15010 11540 15016 11552
rect 14971 11512 15016 11540
rect 14645 11503 14703 11509
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 15160 11512 15205 11540
rect 15160 11500 15166 11512
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 3326 11296 3332 11348
rect 3384 11336 3390 11348
rect 5077 11339 5135 11345
rect 5077 11336 5089 11339
rect 3384 11308 5089 11336
rect 3384 11296 3390 11308
rect 5077 11305 5089 11308
rect 5123 11305 5135 11339
rect 5077 11299 5135 11305
rect 5445 11339 5503 11345
rect 5445 11305 5457 11339
rect 5491 11336 5503 11339
rect 7650 11336 7656 11348
rect 5491 11308 7656 11336
rect 5491 11305 5503 11308
rect 5445 11299 5503 11305
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 8570 11336 8576 11348
rect 8531 11308 8576 11336
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 11609 11339 11667 11345
rect 11609 11336 11621 11339
rect 8720 11308 11621 11336
rect 8720 11296 8726 11308
rect 11609 11305 11621 11308
rect 11655 11305 11667 11339
rect 11609 11299 11667 11305
rect 1394 11228 1400 11280
rect 1452 11268 1458 11280
rect 1857 11271 1915 11277
rect 1857 11268 1869 11271
rect 1452 11240 1869 11268
rect 1452 11228 1458 11240
rect 1857 11237 1869 11240
rect 1903 11237 1915 11271
rect 1857 11231 1915 11237
rect 4525 11271 4583 11277
rect 4525 11237 4537 11271
rect 4571 11268 4583 11271
rect 4614 11268 4620 11280
rect 4571 11240 4620 11268
rect 4571 11237 4583 11240
rect 4525 11231 4583 11237
rect 4614 11228 4620 11240
rect 4672 11228 4678 11280
rect 5258 11228 5264 11280
rect 5316 11268 5322 11280
rect 5537 11271 5595 11277
rect 5537 11268 5549 11271
rect 5316 11240 5549 11268
rect 5316 11228 5322 11240
rect 5537 11237 5549 11240
rect 5583 11237 5595 11271
rect 5537 11231 5595 11237
rect 5902 11228 5908 11280
rect 5960 11268 5966 11280
rect 11422 11268 11428 11280
rect 5960 11240 11428 11268
rect 5960 11228 5966 11240
rect 11422 11228 11428 11240
rect 11480 11228 11486 11280
rect 11624 11268 11652 11299
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 12161 11339 12219 11345
rect 12161 11336 12173 11339
rect 11756 11308 12173 11336
rect 11756 11296 11762 11308
rect 12161 11305 12173 11308
rect 12207 11305 12219 11339
rect 12161 11299 12219 11305
rect 12250 11296 12256 11348
rect 12308 11336 12314 11348
rect 13449 11339 13507 11345
rect 13449 11336 13461 11339
rect 12308 11308 13461 11336
rect 12308 11296 12314 11308
rect 13449 11305 13461 11308
rect 13495 11305 13507 11339
rect 13814 11336 13820 11348
rect 13775 11308 13820 11336
rect 13449 11299 13507 11305
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 14274 11336 14280 11348
rect 14235 11308 14280 11336
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 12710 11268 12716 11280
rect 11624 11240 12716 11268
rect 12710 11228 12716 11240
rect 12768 11228 12774 11280
rect 12802 11228 12808 11280
rect 12860 11228 12866 11280
rect 12894 11228 12900 11280
rect 12952 11268 12958 11280
rect 13357 11271 13415 11277
rect 13357 11268 13369 11271
rect 12952 11240 13369 11268
rect 12952 11228 12958 11240
rect 13357 11237 13369 11240
rect 13403 11237 13415 11271
rect 13357 11231 13415 11237
rect 14185 11271 14243 11277
rect 14185 11237 14197 11271
rect 14231 11268 14243 11271
rect 14550 11268 14556 11280
rect 14231 11240 14556 11268
rect 14231 11237 14243 11240
rect 14185 11231 14243 11237
rect 14550 11228 14556 11240
rect 14608 11228 14614 11280
rect 1578 11200 1584 11212
rect 1539 11172 1584 11200
rect 1578 11160 1584 11172
rect 1636 11160 1642 11212
rect 2584 11203 2642 11209
rect 2584 11169 2596 11203
rect 2630 11200 2642 11203
rect 4433 11203 4491 11209
rect 2630 11172 4108 11200
rect 2630 11169 2642 11172
rect 2584 11163 2642 11169
rect 4080 11144 4108 11172
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 4890 11200 4896 11212
rect 4479 11172 4896 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 4890 11160 4896 11172
rect 4948 11160 4954 11212
rect 6454 11200 6460 11212
rect 6415 11172 6460 11200
rect 6454 11160 6460 11172
rect 6512 11160 6518 11212
rect 6549 11203 6607 11209
rect 6549 11169 6561 11203
rect 6595 11200 6607 11203
rect 6914 11200 6920 11212
rect 6595 11172 6920 11200
rect 6595 11169 6607 11172
rect 6549 11163 6607 11169
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7282 11200 7288 11212
rect 7243 11172 7288 11200
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 7745 11203 7803 11209
rect 7745 11169 7757 11203
rect 7791 11200 7803 11203
rect 8570 11200 8576 11212
rect 7791 11172 8576 11200
rect 7791 11169 7803 11172
rect 7745 11163 7803 11169
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 8938 11200 8944 11212
rect 8899 11172 8944 11200
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 9030 11160 9036 11212
rect 9088 11200 9094 11212
rect 9490 11200 9496 11212
rect 9088 11172 9496 11200
rect 9088 11160 9094 11172
rect 9490 11160 9496 11172
rect 9548 11160 9554 11212
rect 10318 11200 10324 11212
rect 10279 11172 10324 11200
rect 10318 11160 10324 11172
rect 10376 11160 10382 11212
rect 12529 11203 12587 11209
rect 12529 11169 12541 11203
rect 12575 11169 12587 11203
rect 12529 11163 12587 11169
rect 12621 11203 12679 11209
rect 12621 11169 12633 11203
rect 12667 11200 12679 11203
rect 12820 11200 12848 11228
rect 13998 11200 14004 11212
rect 12667 11172 12848 11200
rect 13832 11172 14004 11200
rect 12667 11169 12679 11172
rect 12621 11163 12679 11169
rect 1670 11092 1676 11144
rect 1728 11132 1734 11144
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 1728 11104 2329 11132
rect 1728 11092 1734 11104
rect 2317 11101 2329 11104
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 4062 11092 4068 11144
rect 4120 11092 4126 11144
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 5629 11135 5687 11141
rect 5629 11101 5641 11135
rect 5675 11101 5687 11135
rect 5629 11095 5687 11101
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11132 6791 11135
rect 7190 11132 7196 11144
rect 6779 11104 7196 11132
rect 6779 11101 6791 11104
rect 6733 11095 6791 11101
rect 4080 11064 4108 11092
rect 4632 11064 4660 11095
rect 4706 11064 4712 11076
rect 4080 11036 4712 11064
rect 4706 11024 4712 11036
rect 4764 11064 4770 11076
rect 5644 11064 5672 11095
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 7374 11092 7380 11144
rect 7432 11132 7438 11144
rect 7837 11135 7895 11141
rect 7837 11132 7849 11135
rect 7432 11104 7849 11132
rect 7432 11092 7438 11104
rect 7837 11101 7849 11104
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11132 8079 11135
rect 8110 11132 8116 11144
rect 8067 11104 8116 11132
rect 8067 11101 8079 11104
rect 8021 11095 8079 11101
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11132 9275 11135
rect 9306 11132 9312 11144
rect 9263 11104 9312 11132
rect 9263 11101 9275 11104
rect 9217 11095 9275 11101
rect 9306 11092 9312 11104
rect 9364 11092 9370 11144
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 11330 11132 11336 11144
rect 9640 11104 11336 11132
rect 9640 11092 9646 11104
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 12250 11092 12256 11144
rect 12308 11132 12314 11144
rect 12544 11132 12572 11163
rect 13832 11144 13860 11172
rect 13998 11160 14004 11172
rect 14056 11160 14062 11212
rect 12308 11104 12572 11132
rect 12713 11135 12771 11141
rect 12308 11092 12314 11104
rect 12713 11101 12725 11135
rect 12759 11101 12771 11135
rect 12713 11095 12771 11101
rect 4764 11036 5672 11064
rect 4764 11024 4770 11036
rect 5718 11024 5724 11076
rect 5776 11064 5782 11076
rect 7101 11067 7159 11073
rect 7101 11064 7113 11067
rect 5776 11036 7113 11064
rect 5776 11024 5782 11036
rect 7101 11033 7113 11036
rect 7147 11033 7159 11067
rect 7392 11064 7420 11092
rect 7101 11027 7159 11033
rect 7208 11036 7420 11064
rect 3694 10996 3700 11008
rect 3655 10968 3700 10996
rect 3694 10956 3700 10968
rect 3752 10956 3758 11008
rect 4062 10996 4068 11008
rect 4023 10968 4068 10996
rect 4062 10956 4068 10968
rect 4120 10956 4126 11008
rect 5902 10956 5908 11008
rect 5960 10996 5966 11008
rect 6089 10999 6147 11005
rect 6089 10996 6101 10999
rect 5960 10968 6101 10996
rect 5960 10956 5966 10968
rect 6089 10965 6101 10968
rect 6135 10965 6147 10999
rect 6089 10959 6147 10965
rect 6638 10956 6644 11008
rect 6696 10996 6702 11008
rect 7208 10996 7236 11036
rect 7650 11024 7656 11076
rect 7708 11064 7714 11076
rect 11146 11064 11152 11076
rect 7708 11036 11152 11064
rect 7708 11024 7714 11036
rect 11146 11024 11152 11036
rect 11204 11064 11210 11076
rect 11204 11036 11836 11064
rect 11204 11024 11210 11036
rect 7374 10996 7380 11008
rect 6696 10968 7236 10996
rect 7335 10968 7380 10996
rect 6696 10956 6702 10968
rect 7374 10956 7380 10968
rect 7432 10956 7438 11008
rect 11808 10996 11836 11036
rect 11882 11024 11888 11076
rect 11940 11064 11946 11076
rect 12719 11064 12747 11095
rect 12894 11092 12900 11144
rect 12952 11132 12958 11144
rect 13170 11132 13176 11144
rect 12952 11104 13176 11132
rect 12952 11092 12958 11104
rect 13170 11092 13176 11104
rect 13228 11092 13234 11144
rect 13262 11092 13268 11144
rect 13320 11132 13326 11144
rect 13541 11135 13599 11141
rect 13541 11132 13553 11135
rect 13320 11104 13553 11132
rect 13320 11092 13326 11104
rect 13541 11101 13553 11104
rect 13587 11132 13599 11135
rect 13814 11132 13820 11144
rect 13587 11104 13820 11132
rect 13587 11101 13599 11104
rect 13541 11095 13599 11101
rect 13814 11092 13820 11104
rect 13872 11092 13878 11144
rect 13906 11092 13912 11144
rect 13964 11132 13970 11144
rect 14369 11135 14427 11141
rect 14369 11132 14381 11135
rect 13964 11104 14381 11132
rect 13964 11092 13970 11104
rect 14369 11101 14381 11104
rect 14415 11101 14427 11135
rect 14642 11132 14648 11144
rect 14603 11104 14648 11132
rect 14369 11095 14427 11101
rect 14642 11092 14648 11104
rect 14700 11092 14706 11144
rect 11940 11036 12747 11064
rect 12989 11067 13047 11073
rect 11940 11024 11946 11036
rect 12989 11033 13001 11067
rect 13035 11064 13047 11067
rect 13354 11064 13360 11076
rect 13035 11036 13360 11064
rect 13035 11033 13047 11036
rect 12989 11027 13047 11033
rect 13354 11024 13360 11036
rect 13412 11024 13418 11076
rect 14550 11064 14556 11076
rect 13464 11036 14556 11064
rect 13464 10996 13492 11036
rect 14550 11024 14556 11036
rect 14608 11024 14614 11076
rect 11808 10968 13492 10996
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 2406 10752 2412 10804
rect 2464 10792 2470 10804
rect 2777 10795 2835 10801
rect 2777 10792 2789 10795
rect 2464 10764 2789 10792
rect 2464 10752 2470 10764
rect 2777 10761 2789 10764
rect 2823 10761 2835 10795
rect 3050 10792 3056 10804
rect 3011 10764 3056 10792
rect 2777 10755 2835 10761
rect 3050 10752 3056 10764
rect 3108 10752 3114 10804
rect 5077 10795 5135 10801
rect 5077 10761 5089 10795
rect 5123 10792 5135 10795
rect 5626 10792 5632 10804
rect 5123 10764 5632 10792
rect 5123 10761 5135 10764
rect 5077 10755 5135 10761
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 9217 10795 9275 10801
rect 9217 10792 9229 10795
rect 7484 10764 9229 10792
rect 4982 10684 4988 10736
rect 5040 10724 5046 10736
rect 6825 10727 6883 10733
rect 6825 10724 6837 10727
rect 5040 10696 6837 10724
rect 5040 10684 5046 10696
rect 6825 10693 6837 10696
rect 6871 10693 6883 10727
rect 6825 10687 6883 10693
rect 3605 10659 3663 10665
rect 3605 10656 3617 10659
rect 3160 10628 3617 10656
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10557 1455 10591
rect 1397 10551 1455 10557
rect 1664 10591 1722 10597
rect 1664 10557 1676 10591
rect 1710 10588 1722 10591
rect 3160 10588 3188 10628
rect 3605 10625 3617 10628
rect 3651 10656 3663 10659
rect 3694 10656 3700 10668
rect 3651 10628 3700 10656
rect 3651 10625 3663 10628
rect 3605 10619 3663 10625
rect 3694 10616 3700 10628
rect 3752 10616 3758 10668
rect 4706 10656 4712 10668
rect 4667 10628 4712 10656
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 5074 10616 5080 10668
rect 5132 10656 5138 10668
rect 5537 10659 5595 10665
rect 5537 10656 5549 10659
rect 5132 10628 5549 10656
rect 5132 10616 5138 10628
rect 5537 10625 5549 10628
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 6089 10659 6147 10665
rect 5684 10628 5729 10656
rect 5684 10616 5690 10628
rect 6089 10625 6101 10659
rect 6135 10656 6147 10659
rect 6454 10656 6460 10668
rect 6135 10628 6460 10656
rect 6135 10625 6147 10628
rect 6089 10619 6147 10625
rect 6454 10616 6460 10628
rect 6512 10616 6518 10668
rect 7484 10665 7512 10764
rect 9217 10761 9229 10764
rect 9263 10761 9275 10795
rect 11054 10792 11060 10804
rect 11015 10764 11060 10792
rect 9217 10755 9275 10761
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10625 7527 10659
rect 9232 10656 9260 10755
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11149 10795 11207 10801
rect 11149 10761 11161 10795
rect 11195 10792 11207 10795
rect 12802 10792 12808 10804
rect 11195 10764 12808 10792
rect 11195 10761 11207 10764
rect 11149 10755 11207 10761
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 13173 10795 13231 10801
rect 13173 10761 13185 10795
rect 13219 10792 13231 10795
rect 15010 10792 15016 10804
rect 13219 10764 15016 10792
rect 13219 10761 13231 10764
rect 13173 10755 13231 10761
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 11072 10656 11100 10752
rect 17494 10724 17500 10736
rect 12636 10696 17500 10724
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 9232 10628 9812 10656
rect 11072 10628 11713 10656
rect 7469 10619 7527 10625
rect 1710 10560 3188 10588
rect 3513 10591 3571 10597
rect 1710 10557 1722 10560
rect 1664 10551 1722 10557
rect 3513 10557 3525 10591
rect 3559 10588 3571 10591
rect 4062 10588 4068 10600
rect 3559 10560 4068 10588
rect 3559 10557 3571 10560
rect 3513 10551 3571 10557
rect 1412 10520 1440 10551
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4338 10548 4344 10600
rect 4396 10588 4402 10600
rect 4525 10591 4583 10597
rect 4525 10588 4537 10591
rect 4396 10560 4537 10588
rect 4396 10548 4402 10560
rect 4525 10557 4537 10560
rect 4571 10588 4583 10591
rect 6546 10588 6552 10600
rect 4571 10560 6552 10588
rect 4571 10557 4583 10560
rect 4525 10551 4583 10557
rect 6546 10548 6552 10560
rect 6604 10548 6610 10600
rect 7193 10591 7251 10597
rect 7193 10557 7205 10591
rect 7239 10588 7251 10591
rect 7374 10588 7380 10600
rect 7239 10560 7380 10588
rect 7239 10557 7251 10560
rect 7193 10551 7251 10557
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 7650 10548 7656 10600
rect 7708 10588 7714 10600
rect 8110 10597 8116 10600
rect 7837 10591 7895 10597
rect 7837 10588 7849 10591
rect 7708 10560 7849 10588
rect 7708 10548 7714 10560
rect 7837 10557 7849 10560
rect 7883 10557 7895 10591
rect 8104 10588 8116 10597
rect 8071 10560 8116 10588
rect 7837 10551 7895 10557
rect 8104 10551 8116 10560
rect 8110 10548 8116 10551
rect 8168 10548 8174 10600
rect 8570 10548 8576 10600
rect 8628 10588 8634 10600
rect 9401 10591 9459 10597
rect 9401 10588 9413 10591
rect 8628 10560 9413 10588
rect 8628 10548 8634 10560
rect 9401 10557 9413 10560
rect 9447 10557 9459 10591
rect 9674 10588 9680 10600
rect 9635 10560 9680 10588
rect 9401 10551 9459 10557
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 9784 10588 9812 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 9933 10591 9991 10597
rect 9933 10588 9945 10591
rect 9784 10560 9945 10588
rect 9933 10557 9945 10560
rect 9979 10557 9991 10591
rect 9933 10551 9991 10557
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 11112 10560 11529 10588
rect 11112 10548 11118 10560
rect 11517 10557 11529 10560
rect 11563 10588 11575 10591
rect 12636 10588 12664 10696
rect 17494 10684 17500 10696
rect 17552 10684 17558 10736
rect 13722 10656 13728 10668
rect 13683 10628 13728 10656
rect 13722 10616 13728 10628
rect 13780 10616 13786 10668
rect 13814 10616 13820 10668
rect 13872 10656 13878 10668
rect 14737 10659 14795 10665
rect 14737 10656 14749 10659
rect 13872 10628 14749 10656
rect 13872 10616 13878 10628
rect 14737 10625 14749 10628
rect 14783 10625 14795 10659
rect 14737 10619 14795 10625
rect 11563 10560 12664 10588
rect 11563 10557 11575 10560
rect 11517 10551 11575 10557
rect 12710 10548 12716 10600
rect 12768 10588 12774 10600
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12768 10560 12817 10588
rect 12768 10548 12774 10560
rect 12805 10557 12817 10560
rect 12851 10557 12863 10591
rect 12805 10551 12863 10557
rect 13541 10591 13599 10597
rect 13541 10557 13553 10591
rect 13587 10588 13599 10591
rect 14642 10588 14648 10600
rect 13587 10560 14648 10588
rect 13587 10557 13599 10560
rect 13541 10551 13599 10557
rect 14642 10548 14648 10560
rect 14700 10548 14706 10600
rect 3421 10523 3479 10529
rect 1412 10492 1716 10520
rect 1688 10464 1716 10492
rect 3421 10489 3433 10523
rect 3467 10520 3479 10523
rect 3467 10492 4108 10520
rect 3467 10489 3479 10492
rect 3421 10483 3479 10489
rect 1670 10412 1676 10464
rect 1728 10412 1734 10464
rect 4080 10461 4108 10492
rect 11698 10480 11704 10532
rect 11756 10520 11762 10532
rect 14553 10523 14611 10529
rect 14553 10520 14565 10523
rect 11756 10492 14565 10520
rect 11756 10480 11762 10492
rect 14553 10489 14565 10492
rect 14599 10489 14611 10523
rect 14553 10483 14611 10489
rect 4065 10455 4123 10461
rect 4065 10421 4077 10455
rect 4111 10421 4123 10455
rect 4430 10452 4436 10464
rect 4391 10424 4436 10452
rect 4065 10415 4123 10421
rect 4430 10412 4436 10424
rect 4488 10412 4494 10464
rect 5445 10455 5503 10461
rect 5445 10421 5457 10455
rect 5491 10452 5503 10455
rect 5902 10452 5908 10464
rect 5491 10424 5908 10452
rect 5491 10421 5503 10424
rect 5445 10415 5503 10421
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 7282 10452 7288 10464
rect 7243 10424 7288 10452
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 8478 10412 8484 10464
rect 8536 10452 8542 10464
rect 9582 10452 9588 10464
rect 8536 10424 9588 10452
rect 8536 10412 8542 10424
rect 9582 10412 9588 10424
rect 9640 10452 9646 10464
rect 11609 10455 11667 10461
rect 11609 10452 11621 10455
rect 9640 10424 11621 10452
rect 9640 10412 9646 10424
rect 11609 10421 11621 10424
rect 11655 10421 11667 10455
rect 12618 10452 12624 10464
rect 12579 10424 12624 10452
rect 11609 10415 11667 10421
rect 12618 10412 12624 10424
rect 12676 10412 12682 10464
rect 13630 10452 13636 10464
rect 13591 10424 13636 10452
rect 13630 10412 13636 10424
rect 13688 10452 13694 10464
rect 13906 10452 13912 10464
rect 13688 10424 13912 10452
rect 13688 10412 13694 10424
rect 13906 10412 13912 10424
rect 13964 10412 13970 10464
rect 14182 10452 14188 10464
rect 14143 10424 14188 10452
rect 14182 10412 14188 10424
rect 14240 10412 14246 10464
rect 14274 10412 14280 10464
rect 14332 10452 14338 10464
rect 14645 10455 14703 10461
rect 14645 10452 14657 10455
rect 14332 10424 14657 10452
rect 14332 10412 14338 10424
rect 14645 10421 14657 10424
rect 14691 10452 14703 10455
rect 16390 10452 16396 10464
rect 14691 10424 16396 10452
rect 14691 10421 14703 10424
rect 14645 10415 14703 10421
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 2866 10248 2872 10260
rect 1627 10220 2872 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 3421 10251 3479 10257
rect 3421 10217 3433 10251
rect 3467 10248 3479 10251
rect 4430 10248 4436 10260
rect 3467 10220 4436 10248
rect 3467 10217 3479 10220
rect 3421 10211 3479 10217
rect 4430 10208 4436 10220
rect 4488 10208 4494 10260
rect 4617 10251 4675 10257
rect 4617 10217 4629 10251
rect 4663 10248 4675 10251
rect 4982 10248 4988 10260
rect 4663 10220 4988 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 4982 10208 4988 10220
rect 5040 10208 5046 10260
rect 8202 10208 8208 10260
rect 8260 10248 8266 10260
rect 8849 10251 8907 10257
rect 8849 10248 8861 10251
rect 8260 10220 8861 10248
rect 8260 10208 8266 10220
rect 8849 10217 8861 10220
rect 8895 10217 8907 10251
rect 10962 10248 10968 10260
rect 8849 10211 8907 10217
rect 9876 10220 10968 10248
rect 4246 10180 4252 10192
rect 1412 10152 4252 10180
rect 1412 10121 1440 10152
rect 4246 10140 4252 10152
rect 4304 10140 4310 10192
rect 5077 10183 5135 10189
rect 5077 10149 5089 10183
rect 5123 10180 5135 10183
rect 5166 10180 5172 10192
rect 5123 10152 5172 10180
rect 5123 10149 5135 10152
rect 5077 10143 5135 10149
rect 5166 10140 5172 10152
rect 5224 10140 5230 10192
rect 5810 10140 5816 10192
rect 5868 10180 5874 10192
rect 6058 10183 6116 10189
rect 6058 10180 6070 10183
rect 5868 10152 6070 10180
rect 5868 10140 5874 10152
rect 6058 10149 6070 10152
rect 6104 10149 6116 10183
rect 9876 10180 9904 10220
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11057 10251 11115 10257
rect 11057 10217 11069 10251
rect 11103 10248 11115 10251
rect 11146 10248 11152 10260
rect 11103 10220 11152 10248
rect 11103 10217 11115 10220
rect 11057 10211 11115 10217
rect 11146 10208 11152 10220
rect 11204 10248 11210 10260
rect 11882 10248 11888 10260
rect 11204 10220 11888 10248
rect 11204 10208 11210 10220
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 14366 10248 14372 10260
rect 14327 10220 14372 10248
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 6058 10143 6116 10149
rect 7116 10152 9904 10180
rect 9944 10183 10002 10189
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10081 1455 10115
rect 1397 10075 1455 10081
rect 2032 10115 2090 10121
rect 2032 10081 2044 10115
rect 2078 10112 2090 10115
rect 2406 10112 2412 10124
rect 2078 10084 2412 10112
rect 2078 10081 2090 10084
rect 2032 10075 2090 10081
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 4982 10112 4988 10124
rect 4943 10084 4988 10112
rect 4982 10072 4988 10084
rect 5040 10072 5046 10124
rect 7116 10112 7144 10152
rect 9944 10149 9956 10183
rect 9990 10180 10002 10183
rect 12434 10180 12440 10192
rect 9990 10152 12440 10180
rect 9990 10149 10002 10152
rect 9944 10143 10002 10149
rect 12434 10140 12440 10152
rect 12492 10140 12498 10192
rect 13234 10183 13292 10189
rect 13234 10180 13246 10183
rect 12728 10152 13246 10180
rect 7736 10115 7794 10121
rect 7736 10112 7748 10115
rect 5184 10084 7144 10112
rect 7208 10084 7748 10112
rect 1670 10004 1676 10056
rect 1728 10044 1734 10056
rect 1765 10047 1823 10053
rect 1765 10044 1777 10047
rect 1728 10016 1777 10044
rect 1728 10004 1734 10016
rect 1765 10013 1777 10016
rect 1811 10013 1823 10047
rect 1765 10007 1823 10013
rect 4062 10004 4068 10056
rect 4120 10044 4126 10056
rect 5184 10044 5212 10084
rect 4120 10016 5212 10044
rect 5261 10047 5319 10053
rect 4120 10004 4126 10016
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 5350 10044 5356 10056
rect 5307 10016 5356 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10013 5871 10047
rect 5813 10007 5871 10013
rect 4798 9936 4804 9988
rect 4856 9976 4862 9988
rect 5828 9976 5856 10007
rect 7208 9985 7236 10084
rect 7736 10081 7748 10084
rect 7782 10112 7794 10115
rect 8478 10112 8484 10124
rect 7782 10084 8484 10112
rect 7782 10081 7794 10084
rect 7736 10075 7794 10081
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 11333 10115 11391 10121
rect 11333 10112 11345 10115
rect 9692 10084 11345 10112
rect 9692 10056 9720 10084
rect 11333 10081 11345 10084
rect 11379 10081 11391 10115
rect 11333 10075 11391 10081
rect 11589 10115 11647 10121
rect 11589 10081 11601 10115
rect 11635 10112 11647 10115
rect 11882 10112 11888 10124
rect 11635 10084 11888 10112
rect 11635 10081 11647 10084
rect 11589 10075 11647 10081
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10013 7527 10047
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 7469 10007 7527 10013
rect 4856 9948 5856 9976
rect 7193 9979 7251 9985
rect 4856 9936 4862 9948
rect 7193 9945 7205 9979
rect 7239 9945 7251 9979
rect 7193 9939 7251 9945
rect 3142 9908 3148 9920
rect 3103 9880 3148 9908
rect 3142 9868 3148 9880
rect 3200 9868 3206 9920
rect 3234 9868 3240 9920
rect 3292 9908 3298 9920
rect 5074 9908 5080 9920
rect 3292 9880 5080 9908
rect 3292 9868 3298 9880
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 7484 9908 7512 10007
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 7650 9908 7656 9920
rect 7484 9880 7656 9908
rect 7650 9868 7656 9880
rect 7708 9908 7714 9920
rect 9674 9908 9680 9920
rect 7708 9880 9680 9908
rect 7708 9868 7714 9880
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 11974 9868 11980 9920
rect 12032 9908 12038 9920
rect 12728 9917 12756 10152
rect 13234 10149 13246 10152
rect 13280 10149 13292 10183
rect 13234 10143 13292 10149
rect 12989 10115 13047 10121
rect 12989 10081 13001 10115
rect 13035 10112 13047 10115
rect 13538 10112 13544 10124
rect 13035 10084 13544 10112
rect 13035 10081 13047 10084
rect 12989 10075 13047 10081
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 12713 9911 12771 9917
rect 12713 9908 12725 9911
rect 12032 9880 12725 9908
rect 12032 9868 12038 9880
rect 12713 9877 12725 9880
rect 12759 9877 12771 9911
rect 12713 9871 12771 9877
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 4157 9707 4215 9713
rect 4157 9673 4169 9707
rect 4203 9704 4215 9707
rect 4706 9704 4712 9716
rect 4203 9676 4712 9704
rect 4203 9673 4215 9676
rect 4157 9667 4215 9673
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 6273 9707 6331 9713
rect 6273 9704 6285 9707
rect 5868 9676 6285 9704
rect 5868 9664 5874 9676
rect 6273 9673 6285 9676
rect 6319 9673 6331 9707
rect 6273 9667 6331 9673
rect 7282 9664 7288 9716
rect 7340 9704 7346 9716
rect 7837 9707 7895 9713
rect 7837 9704 7849 9707
rect 7340 9676 7849 9704
rect 7340 9664 7346 9676
rect 7837 9673 7849 9676
rect 7883 9673 7895 9707
rect 7837 9667 7895 9673
rect 8294 9664 8300 9716
rect 8352 9704 8358 9716
rect 11146 9704 11152 9716
rect 8352 9676 10272 9704
rect 8352 9664 8358 9676
rect 1765 9639 1823 9645
rect 1765 9605 1777 9639
rect 1811 9636 1823 9639
rect 2774 9636 2780 9648
rect 1811 9608 2780 9636
rect 1811 9605 1823 9608
rect 1765 9599 1823 9605
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 4617 9639 4675 9645
rect 4617 9605 4629 9639
rect 4663 9636 4675 9639
rect 4798 9636 4804 9648
rect 4663 9608 4804 9636
rect 4663 9605 4675 9608
rect 4617 9599 4675 9605
rect 2314 9568 2320 9580
rect 2275 9540 2320 9568
rect 2314 9528 2320 9540
rect 2372 9528 2378 9580
rect 1670 9460 1676 9512
rect 1728 9500 1734 9512
rect 2777 9503 2835 9509
rect 2777 9500 2789 9503
rect 1728 9472 2789 9500
rect 1728 9460 1734 9472
rect 2777 9469 2789 9472
rect 2823 9500 2835 9503
rect 4724 9500 4752 9608
rect 4798 9596 4804 9608
rect 4856 9596 4862 9648
rect 6638 9596 6644 9648
rect 6696 9596 6702 9648
rect 6822 9636 6828 9648
rect 6783 9608 6828 9636
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 7098 9596 7104 9648
rect 7156 9636 7162 9648
rect 9766 9636 9772 9648
rect 7156 9608 9772 9636
rect 7156 9596 7162 9608
rect 9766 9596 9772 9608
rect 9824 9596 9830 9648
rect 4816 9540 5028 9568
rect 4816 9509 4844 9540
rect 2823 9472 4752 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 2133 9435 2191 9441
rect 2133 9401 2145 9435
rect 2179 9432 2191 9435
rect 2498 9432 2504 9444
rect 2179 9404 2504 9432
rect 2179 9401 2191 9404
rect 2133 9395 2191 9401
rect 2498 9392 2504 9404
rect 2556 9392 2562 9444
rect 3044 9435 3102 9441
rect 3044 9401 3056 9435
rect 3090 9432 3102 9435
rect 3234 9432 3240 9444
rect 3090 9404 3240 9432
rect 3090 9401 3102 9404
rect 3044 9395 3102 9401
rect 3234 9392 3240 9404
rect 3292 9392 3298 9444
rect 4724 9432 4752 9472
rect 4801 9503 4859 9509
rect 4801 9469 4813 9503
rect 4847 9469 4859 9503
rect 4801 9463 4859 9469
rect 4893 9503 4951 9509
rect 4893 9469 4905 9503
rect 4939 9469 4951 9503
rect 5000 9500 5028 9540
rect 5718 9500 5724 9512
rect 5000 9472 5724 9500
rect 4893 9463 4951 9469
rect 4908 9432 4936 9463
rect 5718 9460 5724 9472
rect 5776 9460 5782 9512
rect 4724 9404 4936 9432
rect 5160 9435 5218 9441
rect 5160 9401 5172 9435
rect 5206 9432 5218 9435
rect 6454 9432 6460 9444
rect 5206 9404 6460 9432
rect 5206 9401 5218 9404
rect 5160 9395 5218 9401
rect 6454 9392 6460 9404
rect 6512 9392 6518 9444
rect 1854 9324 1860 9376
rect 1912 9364 1918 9376
rect 2225 9367 2283 9373
rect 2225 9364 2237 9367
rect 1912 9336 2237 9364
rect 1912 9324 1918 9336
rect 2225 9333 2237 9336
rect 2271 9333 2283 9367
rect 2225 9327 2283 9333
rect 5350 9324 5356 9376
rect 5408 9364 5414 9376
rect 6656 9364 6684 9596
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 7469 9571 7527 9577
rect 6788 9540 7144 9568
rect 6788 9528 6794 9540
rect 7116 9432 7144 9540
rect 7469 9537 7481 9571
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 7484 9500 7512 9531
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 8389 9571 8447 9577
rect 8389 9568 8401 9571
rect 8260 9540 8401 9568
rect 8260 9528 8266 9540
rect 8389 9537 8401 9540
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 8754 9528 8760 9580
rect 8812 9568 8818 9580
rect 9950 9568 9956 9580
rect 8812 9540 9956 9568
rect 8812 9528 8818 9540
rect 9950 9528 9956 9540
rect 10008 9528 10014 9580
rect 10244 9577 10272 9676
rect 11072 9676 11152 9704
rect 11072 9577 11100 9676
rect 11146 9664 11152 9676
rect 11204 9664 11210 9716
rect 12176 9676 12664 9704
rect 11882 9596 11888 9648
rect 11940 9636 11946 9648
rect 12176 9636 12204 9676
rect 11940 9608 12204 9636
rect 12253 9639 12311 9645
rect 11940 9596 11946 9608
rect 12253 9605 12265 9639
rect 12299 9636 12311 9639
rect 12437 9639 12495 9645
rect 12437 9636 12449 9639
rect 12299 9608 12449 9636
rect 12299 9605 12311 9608
rect 12253 9599 12311 9605
rect 12437 9605 12449 9608
rect 12483 9605 12495 9639
rect 12437 9599 12495 9605
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9537 10287 9571
rect 10229 9531 10287 9537
rect 10965 9571 11023 9577
rect 10965 9537 10977 9571
rect 11011 9537 11023 9571
rect 10965 9531 11023 9537
rect 11057 9571 11115 9577
rect 11057 9537 11069 9571
rect 11103 9537 11115 9571
rect 11057 9531 11115 9537
rect 10042 9500 10048 9512
rect 7484 9472 10048 9500
rect 10042 9460 10048 9472
rect 10100 9460 10106 9512
rect 10980 9500 11008 9531
rect 11514 9528 11520 9580
rect 11572 9568 11578 9580
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11572 9540 11805 9568
rect 11572 9528 11578 9540
rect 11793 9537 11805 9540
rect 11839 9537 11851 9571
rect 11974 9568 11980 9580
rect 11935 9540 11980 9568
rect 11793 9531 11851 9537
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 12526 9568 12532 9580
rect 12084 9540 12532 9568
rect 12084 9500 12112 9540
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12636 9568 12664 9676
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 12636 9540 12909 9568
rect 12897 9537 12909 9540
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 10980 9472 12112 9500
rect 12158 9460 12164 9512
rect 12216 9500 12222 9512
rect 13004 9500 13032 9531
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 14001 9571 14059 9577
rect 14001 9568 14013 9571
rect 13780 9540 14013 9568
rect 13780 9528 13786 9540
rect 14001 9537 14013 9540
rect 14047 9537 14059 9571
rect 14001 9531 14059 9537
rect 14090 9528 14096 9580
rect 14148 9568 14154 9580
rect 14550 9568 14556 9580
rect 14148 9540 14556 9568
rect 14148 9528 14154 9540
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 15010 9568 15016 9580
rect 14971 9540 15016 9568
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 12216 9472 13032 9500
rect 13357 9503 13415 9509
rect 12216 9460 12222 9472
rect 13357 9469 13369 9503
rect 13403 9500 13415 9503
rect 15102 9500 15108 9512
rect 13403 9472 15108 9500
rect 13403 9469 13415 9472
rect 13357 9463 13415 9469
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 7558 9432 7564 9444
rect 7116 9404 7564 9432
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 8205 9435 8263 9441
rect 8205 9401 8217 9435
rect 8251 9432 8263 9435
rect 8846 9432 8852 9444
rect 8251 9404 8852 9432
rect 8251 9401 8263 9404
rect 8205 9395 8263 9401
rect 8846 9392 8852 9404
rect 8904 9392 8910 9444
rect 8938 9392 8944 9444
rect 8996 9432 9002 9444
rect 10873 9435 10931 9441
rect 8996 9404 9996 9432
rect 8996 9392 9002 9404
rect 9968 9376 9996 9404
rect 10873 9401 10885 9435
rect 10919 9432 10931 9435
rect 11701 9435 11759 9441
rect 10919 9404 11652 9432
rect 10919 9401 10931 9404
rect 10873 9395 10931 9401
rect 7190 9364 7196 9376
rect 5408 9336 6684 9364
rect 7151 9336 7196 9364
rect 5408 9324 5414 9336
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 8294 9364 8300 9376
rect 7340 9336 7385 9364
rect 8255 9336 8300 9364
rect 7340 9324 7346 9336
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 9677 9367 9735 9373
rect 9677 9333 9689 9367
rect 9723 9364 9735 9367
rect 9858 9364 9864 9376
rect 9723 9336 9864 9364
rect 9723 9333 9735 9336
rect 9677 9327 9735 9333
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 10045 9367 10103 9373
rect 10045 9364 10057 9367
rect 10008 9336 10057 9364
rect 10008 9324 10014 9336
rect 10045 9333 10057 9336
rect 10091 9333 10103 9367
rect 10045 9327 10103 9333
rect 10134 9324 10140 9376
rect 10192 9364 10198 9376
rect 10502 9364 10508 9376
rect 10192 9336 10237 9364
rect 10463 9336 10508 9364
rect 10192 9324 10198 9336
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 11330 9364 11336 9376
rect 11291 9336 11336 9364
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 11624 9364 11652 9404
rect 11701 9401 11713 9435
rect 11747 9432 11759 9435
rect 12253 9435 12311 9441
rect 12253 9432 12265 9435
rect 11747 9404 12265 9432
rect 11747 9401 11759 9404
rect 11701 9395 11759 9401
rect 12253 9401 12265 9404
rect 12299 9401 12311 9435
rect 14182 9432 14188 9444
rect 12253 9395 12311 9401
rect 12544 9404 14188 9432
rect 12544 9364 12572 9404
rect 14182 9392 14188 9404
rect 14240 9392 14246 9444
rect 14642 9392 14648 9444
rect 14700 9432 14706 9444
rect 14921 9435 14979 9441
rect 14921 9432 14933 9435
rect 14700 9404 14933 9432
rect 14700 9392 14706 9404
rect 14921 9401 14933 9404
rect 14967 9401 14979 9435
rect 14921 9395 14979 9401
rect 11624 9336 12572 9364
rect 12710 9324 12716 9376
rect 12768 9364 12774 9376
rect 12805 9367 12863 9373
rect 12805 9364 12817 9367
rect 12768 9336 12817 9364
rect 12768 9324 12774 9336
rect 12805 9333 12817 9336
rect 12851 9333 12863 9367
rect 12805 9327 12863 9333
rect 13357 9367 13415 9373
rect 13357 9333 13369 9367
rect 13403 9364 13415 9367
rect 13449 9367 13507 9373
rect 13449 9364 13461 9367
rect 13403 9336 13461 9364
rect 13403 9333 13415 9336
rect 13357 9327 13415 9333
rect 13449 9333 13461 9336
rect 13495 9333 13507 9367
rect 13449 9327 13507 9333
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 13817 9367 13875 9373
rect 13817 9364 13829 9367
rect 13780 9336 13829 9364
rect 13780 9324 13786 9336
rect 13817 9333 13829 9336
rect 13863 9333 13875 9367
rect 13817 9327 13875 9333
rect 13909 9367 13967 9373
rect 13909 9333 13921 9367
rect 13955 9364 13967 9367
rect 13998 9364 14004 9376
rect 13955 9336 14004 9364
rect 13955 9333 13967 9336
rect 13909 9327 13967 9333
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 14458 9364 14464 9376
rect 14419 9336 14464 9364
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 14550 9324 14556 9376
rect 14608 9364 14614 9376
rect 14829 9367 14887 9373
rect 14829 9364 14841 9367
rect 14608 9336 14841 9364
rect 14608 9324 14614 9336
rect 14829 9333 14841 9336
rect 14875 9333 14887 9367
rect 14829 9327 14887 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 1854 9160 1860 9172
rect 1815 9132 1860 9160
rect 1854 9120 1860 9132
rect 1912 9120 1918 9172
rect 2498 9120 2504 9172
rect 2556 9160 2562 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 2556 9132 4077 9160
rect 2556 9120 2562 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 7101 9163 7159 9169
rect 7101 9129 7113 9163
rect 7147 9160 7159 9163
rect 7374 9160 7380 9172
rect 7147 9132 7380 9160
rect 7147 9129 7159 9132
rect 7101 9123 7159 9129
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 7929 9163 7987 9169
rect 7929 9129 7941 9163
rect 7975 9160 7987 9163
rect 8294 9160 8300 9172
rect 7975 9132 8300 9160
rect 7975 9129 7987 9132
rect 7929 9123 7987 9129
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 8389 9163 8447 9169
rect 8389 9129 8401 9163
rect 8435 9160 8447 9163
rect 8757 9163 8815 9169
rect 8757 9160 8769 9163
rect 8435 9132 8769 9160
rect 8435 9129 8447 9132
rect 8389 9123 8447 9129
rect 8757 9129 8769 9132
rect 8803 9160 8815 9163
rect 10870 9160 10876 9172
rect 8803 9132 10876 9160
rect 8803 9129 8815 9132
rect 8757 9123 8815 9129
rect 10870 9120 10876 9132
rect 10928 9120 10934 9172
rect 10962 9120 10968 9172
rect 11020 9160 11026 9172
rect 12158 9160 12164 9172
rect 11020 9132 11065 9160
rect 12119 9132 12164 9160
rect 11020 9120 11026 9132
rect 12158 9120 12164 9132
rect 12216 9120 12222 9172
rect 12710 9160 12716 9172
rect 12671 9132 12716 9160
rect 12710 9120 12716 9132
rect 12768 9120 12774 9172
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 13725 9163 13783 9169
rect 13725 9160 13737 9163
rect 13044 9132 13737 9160
rect 13044 9120 13050 9132
rect 13725 9129 13737 9132
rect 13771 9129 13783 9163
rect 13725 9123 13783 9129
rect 14093 9163 14151 9169
rect 14093 9129 14105 9163
rect 14139 9160 14151 9163
rect 14274 9160 14280 9172
rect 14139 9132 14280 9160
rect 14139 9129 14151 9132
rect 14093 9123 14151 9129
rect 14274 9120 14280 9132
rect 14332 9120 14338 9172
rect 2130 9052 2136 9104
rect 2188 9092 2194 9104
rect 2225 9095 2283 9101
rect 2225 9092 2237 9095
rect 2188 9064 2237 9092
rect 2188 9052 2194 9064
rect 2225 9061 2237 9064
rect 2271 9061 2283 9095
rect 2225 9055 2283 9061
rect 4246 9052 4252 9104
rect 4304 9092 4310 9104
rect 4982 9092 4988 9104
rect 4304 9064 4988 9092
rect 4304 9052 4310 9064
rect 4982 9052 4988 9064
rect 5040 9092 5046 9104
rect 5445 9095 5503 9101
rect 5445 9092 5457 9095
rect 5040 9064 5457 9092
rect 5040 9052 5046 9064
rect 5445 9061 5457 9064
rect 5491 9061 5503 9095
rect 5445 9055 5503 9061
rect 6089 9095 6147 9101
rect 6089 9061 6101 9095
rect 6135 9092 6147 9095
rect 10137 9095 10195 9101
rect 6135 9064 9260 9092
rect 6135 9061 6147 9064
rect 6089 9055 6147 9061
rect 3237 9027 3295 9033
rect 3237 8993 3249 9027
rect 3283 9024 3295 9027
rect 3878 9024 3884 9036
rect 3283 8996 3884 9024
rect 3283 8993 3295 8996
rect 3237 8987 3295 8993
rect 3878 8984 3884 8996
rect 3936 8984 3942 9036
rect 4154 8984 4160 9036
rect 4212 9024 4218 9036
rect 4433 9027 4491 9033
rect 4433 9024 4445 9027
rect 4212 8996 4445 9024
rect 4212 8984 4218 8996
rect 4433 8993 4445 8996
rect 4479 8993 4491 9027
rect 6362 9024 6368 9036
rect 4433 8987 4491 8993
rect 4540 8996 6368 9024
rect 1946 8916 1952 8968
rect 2004 8956 2010 8968
rect 2317 8959 2375 8965
rect 2317 8956 2329 8959
rect 2004 8928 2329 8956
rect 2004 8916 2010 8928
rect 2317 8925 2329 8928
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8956 2559 8959
rect 2866 8956 2872 8968
rect 2547 8928 2872 8956
rect 2547 8925 2559 8928
rect 2501 8919 2559 8925
rect 2866 8916 2872 8928
rect 2924 8956 2930 8968
rect 3142 8956 3148 8968
rect 2924 8928 3148 8956
rect 2924 8916 2930 8928
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 3326 8956 3332 8968
rect 3287 8928 3332 8956
rect 3326 8916 3332 8928
rect 3384 8916 3390 8968
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 3436 8888 3464 8919
rect 3602 8916 3608 8968
rect 3660 8956 3666 8968
rect 4540 8965 4568 8996
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 9024 7251 9027
rect 7239 8996 7604 9024
rect 7239 8993 7251 8996
rect 7193 8987 7251 8993
rect 4525 8959 4583 8965
rect 4525 8956 4537 8959
rect 3660 8928 4537 8956
rect 3660 8916 3666 8928
rect 4525 8925 4537 8928
rect 4571 8925 4583 8959
rect 4706 8956 4712 8968
rect 4667 8928 4712 8956
rect 4525 8919 4583 8925
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 4798 8916 4804 8968
rect 4856 8956 4862 8968
rect 5166 8956 5172 8968
rect 4856 8928 5172 8956
rect 4856 8916 4862 8928
rect 5166 8916 5172 8928
rect 5224 8956 5230 8968
rect 5537 8959 5595 8965
rect 5537 8956 5549 8959
rect 5224 8928 5549 8956
rect 5224 8916 5230 8928
rect 5537 8925 5549 8928
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 5721 8959 5779 8965
rect 5721 8925 5733 8959
rect 5767 8956 5779 8959
rect 6730 8956 6736 8968
rect 5767 8928 6736 8956
rect 5767 8925 5779 8928
rect 5721 8919 5779 8925
rect 6730 8916 6736 8928
rect 6788 8916 6794 8968
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 7466 8956 7472 8968
rect 7423 8928 7472 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 7576 8956 7604 8996
rect 7650 8984 7656 9036
rect 7708 9024 7714 9036
rect 7834 9024 7840 9036
rect 7708 8996 7840 9024
rect 7708 8984 7714 8996
rect 7834 8984 7840 8996
rect 7892 8984 7898 9036
rect 8297 9027 8355 9033
rect 8297 8993 8309 9027
rect 8343 9024 8355 9027
rect 8754 9024 8760 9036
rect 8343 8996 8760 9024
rect 8343 8993 8355 8996
rect 8297 8987 8355 8993
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 9125 9027 9183 9033
rect 9125 8993 9137 9027
rect 9171 8993 9183 9027
rect 9232 9024 9260 9064
rect 10137 9061 10149 9095
rect 10183 9092 10195 9095
rect 13081 9095 13139 9101
rect 13081 9092 13093 9095
rect 10183 9064 13093 9092
rect 10183 9061 10195 9064
rect 10137 9055 10195 9061
rect 13081 9061 13093 9064
rect 13127 9061 13139 9095
rect 13081 9055 13139 9061
rect 13173 9095 13231 9101
rect 13173 9061 13185 9095
rect 13219 9092 13231 9095
rect 13354 9092 13360 9104
rect 13219 9064 13360 9092
rect 13219 9061 13231 9064
rect 13173 9055 13231 9061
rect 13354 9052 13360 9064
rect 13412 9052 13418 9104
rect 10594 9024 10600 9036
rect 9232 8996 10600 9024
rect 9125 8987 9183 8993
rect 8386 8956 8392 8968
rect 7576 8928 8392 8956
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 8478 8916 8484 8968
rect 8536 8956 8542 8968
rect 9140 8956 9168 8987
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 10778 8984 10784 9036
rect 10836 9024 10842 9036
rect 11057 9027 11115 9033
rect 11057 9024 11069 9027
rect 10836 8996 11069 9024
rect 10836 8984 10842 8996
rect 11057 8993 11069 8996
rect 11103 9024 11115 9027
rect 12066 9024 12072 9036
rect 11103 8996 11744 9024
rect 12027 8996 12072 9024
rect 11103 8993 11115 8996
rect 11057 8987 11115 8993
rect 10410 8956 10416 8968
rect 8536 8928 8581 8956
rect 9140 8928 10416 8956
rect 8536 8916 8542 8928
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 11716 8956 11744 8996
rect 12066 8984 12072 8996
rect 12124 8984 12130 9036
rect 14366 9024 14372 9036
rect 12176 8996 14372 9024
rect 12176 8956 12204 8996
rect 14366 8984 14372 8996
rect 14424 8984 14430 9036
rect 11204 8928 11249 8956
rect 11716 8928 12204 8956
rect 12345 8959 12403 8965
rect 11204 8916 11210 8928
rect 12345 8925 12357 8959
rect 12391 8956 12403 8959
rect 12434 8956 12440 8968
rect 12391 8928 12440 8956
rect 12391 8925 12403 8928
rect 12345 8919 12403 8925
rect 12434 8916 12440 8928
rect 12492 8916 12498 8968
rect 13262 8956 13268 8968
rect 13223 8928 13268 8956
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 14182 8956 14188 8968
rect 14143 8928 14188 8956
rect 14182 8916 14188 8928
rect 14240 8916 14246 8968
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8956 14335 8959
rect 15010 8956 15016 8968
rect 14323 8928 15016 8956
rect 14323 8925 14335 8928
rect 14277 8919 14335 8925
rect 2464 8860 3464 8888
rect 2464 8848 2470 8860
rect 4062 8848 4068 8900
rect 4120 8888 4126 8900
rect 10134 8888 10140 8900
rect 4120 8860 10140 8888
rect 4120 8848 4126 8860
rect 10134 8848 10140 8860
rect 10192 8888 10198 8900
rect 10502 8888 10508 8900
rect 10192 8860 10508 8888
rect 10192 8848 10198 8860
rect 10502 8848 10508 8860
rect 10560 8848 10566 8900
rect 10597 8891 10655 8897
rect 10597 8857 10609 8891
rect 10643 8888 10655 8891
rect 12894 8888 12900 8900
rect 10643 8860 12900 8888
rect 10643 8857 10655 8860
rect 10597 8851 10655 8857
rect 12894 8848 12900 8860
rect 12952 8848 12958 8900
rect 12986 8848 12992 8900
rect 13044 8888 13050 8900
rect 14292 8888 14320 8919
rect 15010 8916 15016 8928
rect 15068 8916 15074 8968
rect 13044 8860 14320 8888
rect 13044 8848 13050 8860
rect 2869 8823 2927 8829
rect 2869 8789 2881 8823
rect 2915 8820 2927 8823
rect 3970 8820 3976 8832
rect 2915 8792 3976 8820
rect 2915 8789 2927 8792
rect 2869 8783 2927 8789
rect 3970 8780 3976 8792
rect 4028 8780 4034 8832
rect 5077 8823 5135 8829
rect 5077 8789 5089 8823
rect 5123 8820 5135 8823
rect 6638 8820 6644 8832
rect 5123 8792 6644 8820
rect 5123 8789 5135 8792
rect 5077 8783 5135 8789
rect 6638 8780 6644 8792
rect 6696 8780 6702 8832
rect 6733 8823 6791 8829
rect 6733 8789 6745 8823
rect 6779 8820 6791 8823
rect 7650 8820 7656 8832
rect 6779 8792 7656 8820
rect 6779 8789 6791 8792
rect 6733 8783 6791 8789
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 7834 8780 7840 8832
rect 7892 8820 7898 8832
rect 8757 8823 8815 8829
rect 8757 8820 8769 8823
rect 7892 8792 8769 8820
rect 7892 8780 7898 8792
rect 8757 8789 8769 8792
rect 8803 8789 8815 8823
rect 8757 8783 8815 8789
rect 8941 8823 8999 8829
rect 8941 8789 8953 8823
rect 8987 8820 8999 8823
rect 9674 8820 9680 8832
rect 8987 8792 9680 8820
rect 8987 8789 8999 8792
rect 8941 8783 8999 8789
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 10778 8820 10784 8832
rect 9824 8792 10784 8820
rect 9824 8780 9830 8792
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 11701 8823 11759 8829
rect 11701 8789 11713 8823
rect 11747 8820 11759 8823
rect 12618 8820 12624 8832
rect 11747 8792 12624 8820
rect 11747 8789 11759 8792
rect 11701 8783 11759 8789
rect 12618 8780 12624 8792
rect 12676 8780 12682 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 2406 8576 2412 8628
rect 2464 8616 2470 8628
rect 3605 8619 3663 8625
rect 3605 8616 3617 8619
rect 2464 8588 3617 8616
rect 2464 8576 2470 8588
rect 3605 8585 3617 8588
rect 3651 8585 3663 8619
rect 3878 8616 3884 8628
rect 3839 8588 3884 8616
rect 3605 8579 3663 8585
rect 3878 8576 3884 8588
rect 3936 8576 3942 8628
rect 5442 8616 5448 8628
rect 5092 8588 5448 8616
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 4706 8480 4712 8492
rect 4479 8452 4712 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 1486 8412 1492 8424
rect 1447 8384 1492 8412
rect 1486 8372 1492 8384
rect 1544 8372 1550 8424
rect 1670 8372 1676 8424
rect 1728 8412 1734 8424
rect 2225 8415 2283 8421
rect 2225 8412 2237 8415
rect 1728 8384 2237 8412
rect 1728 8372 1734 8384
rect 2225 8381 2237 8384
rect 2271 8381 2283 8415
rect 2225 8375 2283 8381
rect 2492 8415 2550 8421
rect 2492 8381 2504 8415
rect 2538 8412 2550 8415
rect 2866 8412 2872 8424
rect 2538 8384 2872 8412
rect 2538 8381 2550 8384
rect 2492 8375 2550 8381
rect 2866 8372 2872 8384
rect 2924 8412 2930 8424
rect 4448 8412 4476 8443
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 5092 8489 5120 8588
rect 5442 8576 5448 8588
rect 5500 8616 5506 8628
rect 6454 8616 6460 8628
rect 5500 8588 6132 8616
rect 6367 8588 6460 8616
rect 5500 8576 5506 8588
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8449 5135 8483
rect 6104 8480 6132 8588
rect 6454 8576 6460 8588
rect 6512 8616 6518 8628
rect 10042 8616 10048 8628
rect 6512 8588 9628 8616
rect 10003 8588 10048 8616
rect 6512 8576 6518 8588
rect 9600 8548 9628 8588
rect 10042 8576 10048 8588
rect 10100 8576 10106 8628
rect 12986 8616 12992 8628
rect 10152 8588 12992 8616
rect 10152 8548 10180 8588
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 13814 8616 13820 8628
rect 13372 8588 13820 8616
rect 10410 8548 10416 8560
rect 9600 8520 10180 8548
rect 10371 8520 10416 8548
rect 10410 8508 10416 8520
rect 10468 8508 10474 8560
rect 12069 8551 12127 8557
rect 12069 8517 12081 8551
rect 12115 8517 12127 8551
rect 12069 8511 12127 8517
rect 12437 8551 12495 8557
rect 12437 8517 12449 8551
rect 12483 8548 12495 8551
rect 13372 8548 13400 8588
rect 13814 8576 13820 8588
rect 13872 8576 13878 8628
rect 14182 8576 14188 8628
rect 14240 8616 14246 8628
rect 14461 8619 14519 8625
rect 14461 8616 14473 8619
rect 14240 8588 14473 8616
rect 14240 8576 14246 8588
rect 14461 8585 14473 8588
rect 14507 8585 14519 8619
rect 14461 8579 14519 8585
rect 12483 8520 13400 8548
rect 13449 8551 13507 8557
rect 12483 8517 12495 8520
rect 12437 8511 12495 8517
rect 13449 8517 13461 8551
rect 13495 8548 13507 8551
rect 16482 8548 16488 8560
rect 13495 8520 16488 8548
rect 13495 8517 13507 8520
rect 13449 8511 13507 8517
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 6104 8452 7021 8480
rect 5077 8443 5135 8449
rect 7009 8449 7021 8452
rect 7055 8449 7067 8483
rect 10689 8483 10747 8489
rect 10689 8480 10701 8483
rect 7009 8443 7067 8449
rect 9692 8452 10701 8480
rect 9692 8424 9720 8452
rect 10689 8449 10701 8452
rect 10735 8449 10747 8483
rect 12084 8480 12112 8511
rect 16482 8508 16488 8520
rect 16540 8508 16546 8560
rect 12710 8480 12716 8492
rect 12084 8452 12716 8480
rect 10689 8443 10747 8449
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 12894 8480 12900 8492
rect 12855 8452 12900 8480
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 12986 8440 12992 8492
rect 13044 8480 13050 8492
rect 13044 8452 13089 8480
rect 13044 8440 13050 8452
rect 13170 8440 13176 8492
rect 13228 8480 13234 8492
rect 13909 8483 13967 8489
rect 13909 8480 13921 8483
rect 13228 8452 13921 8480
rect 13228 8440 13234 8452
rect 13909 8449 13921 8452
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8449 14151 8483
rect 15010 8480 15016 8492
rect 14971 8452 15016 8480
rect 14093 8443 14151 8449
rect 2924 8384 4476 8412
rect 5344 8415 5402 8421
rect 2924 8372 2930 8384
rect 5344 8381 5356 8415
rect 5390 8412 5402 8415
rect 5626 8412 5632 8424
rect 5390 8384 5632 8412
rect 5390 8381 5402 8384
rect 5344 8375 5402 8381
rect 5626 8372 5632 8384
rect 5684 8372 5690 8424
rect 8665 8415 8723 8421
rect 8665 8381 8677 8415
rect 8711 8412 8723 8415
rect 9674 8412 9680 8424
rect 8711 8384 9680 8412
rect 8711 8381 8723 8384
rect 8665 8375 8723 8381
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 10597 8415 10655 8421
rect 10597 8381 10609 8415
rect 10643 8381 10655 8415
rect 12526 8412 12532 8424
rect 10597 8375 10655 8381
rect 10888 8384 12532 8412
rect 1765 8347 1823 8353
rect 1765 8313 1777 8347
rect 1811 8344 1823 8347
rect 3510 8344 3516 8356
rect 1811 8316 3516 8344
rect 1811 8313 1823 8316
rect 1765 8307 1823 8313
rect 3510 8304 3516 8316
rect 3568 8304 3574 8356
rect 4341 8347 4399 8353
rect 4341 8313 4353 8347
rect 4387 8344 4399 8347
rect 7098 8344 7104 8356
rect 4387 8316 7104 8344
rect 4387 8313 4399 8316
rect 4341 8307 4399 8313
rect 5644 8288 5672 8316
rect 7098 8304 7104 8316
rect 7156 8304 7162 8356
rect 7276 8347 7334 8353
rect 7276 8313 7288 8347
rect 7322 8344 7334 8347
rect 7466 8344 7472 8356
rect 7322 8316 7472 8344
rect 7322 8313 7334 8316
rect 7276 8307 7334 8313
rect 7466 8304 7472 8316
rect 7524 8304 7530 8356
rect 8910 8347 8968 8353
rect 8910 8344 8922 8347
rect 8404 8316 8922 8344
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 4249 8279 4307 8285
rect 4249 8276 4261 8279
rect 4120 8248 4261 8276
rect 4120 8236 4126 8248
rect 4249 8245 4261 8248
rect 4295 8276 4307 8279
rect 5350 8276 5356 8288
rect 4295 8248 5356 8276
rect 4295 8245 4307 8248
rect 4249 8239 4307 8245
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 5626 8236 5632 8288
rect 5684 8236 5690 8288
rect 6270 8236 6276 8288
rect 6328 8276 6334 8288
rect 6546 8276 6552 8288
rect 6328 8248 6552 8276
rect 6328 8236 6334 8248
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 8294 8236 8300 8288
rect 8352 8276 8358 8288
rect 8404 8285 8432 8316
rect 8910 8313 8922 8316
rect 8956 8313 8968 8347
rect 10612 8344 10640 8375
rect 10888 8344 10916 8384
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12676 8384 12817 8412
rect 12676 8372 12682 8384
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 14108 8412 14136 8443
rect 15010 8440 15016 8452
rect 15068 8440 15074 8492
rect 14108 8384 15056 8412
rect 12805 8375 12863 8381
rect 15028 8356 15056 8384
rect 10612 8316 10916 8344
rect 10956 8347 11014 8353
rect 8910 8307 8968 8313
rect 10956 8313 10968 8347
rect 11002 8344 11014 8347
rect 11146 8344 11152 8356
rect 11002 8316 11152 8344
rect 11002 8313 11014 8316
rect 10956 8307 11014 8313
rect 11146 8304 11152 8316
rect 11204 8344 11210 8356
rect 11606 8344 11612 8356
rect 11204 8316 11612 8344
rect 11204 8304 11210 8316
rect 11606 8304 11612 8316
rect 11664 8344 11670 8356
rect 12434 8344 12440 8356
rect 11664 8316 12440 8344
rect 11664 8304 11670 8316
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 12894 8304 12900 8356
rect 12952 8344 12958 8356
rect 12952 8316 14964 8344
rect 12952 8304 12958 8316
rect 8389 8279 8447 8285
rect 8389 8276 8401 8279
rect 8352 8248 8401 8276
rect 8352 8236 8358 8248
rect 8389 8245 8401 8248
rect 8435 8245 8447 8279
rect 8389 8239 8447 8245
rect 8570 8236 8576 8288
rect 8628 8276 8634 8288
rect 13817 8279 13875 8285
rect 13817 8276 13829 8279
rect 8628 8248 13829 8276
rect 8628 8236 8634 8248
rect 13817 8245 13829 8248
rect 13863 8245 13875 8279
rect 13817 8239 13875 8245
rect 14090 8236 14096 8288
rect 14148 8276 14154 8288
rect 14936 8285 14964 8316
rect 15010 8304 15016 8356
rect 15068 8304 15074 8356
rect 14829 8279 14887 8285
rect 14829 8276 14841 8279
rect 14148 8248 14841 8276
rect 14148 8236 14154 8248
rect 14829 8245 14841 8248
rect 14875 8245 14887 8279
rect 14829 8239 14887 8245
rect 14921 8279 14979 8285
rect 14921 8245 14933 8279
rect 14967 8276 14979 8279
rect 15194 8276 15200 8288
rect 14967 8248 15200 8276
rect 14967 8245 14979 8248
rect 14921 8239 14979 8245
rect 15194 8236 15200 8248
rect 15252 8276 15258 8288
rect 16666 8276 16672 8288
rect 15252 8248 16672 8276
rect 15252 8236 15258 8248
rect 16666 8236 16672 8248
rect 16724 8236 16730 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 3326 8032 3332 8084
rect 3384 8072 3390 8084
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 3384 8044 4077 8072
rect 3384 8032 3390 8044
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 4154 8032 4160 8084
rect 4212 8032 4218 8084
rect 5537 8075 5595 8081
rect 5537 8041 5549 8075
rect 5583 8072 5595 8075
rect 6181 8075 6239 8081
rect 6181 8072 6193 8075
rect 5583 8044 6193 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 6181 8041 6193 8044
rect 6227 8041 6239 8075
rect 6638 8072 6644 8084
rect 6599 8044 6644 8072
rect 6181 8035 6239 8041
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 7282 8032 7288 8084
rect 7340 8072 7346 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7340 8044 7757 8072
rect 7340 8032 7346 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 11882 8072 11888 8084
rect 10836 8044 11888 8072
rect 10836 8032 10842 8044
rect 11882 8032 11888 8044
rect 11940 8032 11946 8084
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 13998 8072 14004 8084
rect 12676 8044 14004 8072
rect 12676 8032 12682 8044
rect 13998 8032 14004 8044
rect 14056 8032 14062 8084
rect 1664 8007 1722 8013
rect 1664 7973 1676 8007
rect 1710 8004 1722 8007
rect 2406 8004 2412 8016
rect 1710 7976 2412 8004
rect 1710 7973 1722 7976
rect 1664 7967 1722 7973
rect 2406 7964 2412 7976
rect 2464 7964 2470 8016
rect 3053 8007 3111 8013
rect 3053 7973 3065 8007
rect 3099 8004 3111 8007
rect 4172 8004 4200 8032
rect 3099 7976 4200 8004
rect 4525 8007 4583 8013
rect 3099 7973 3111 7976
rect 3053 7967 3111 7973
rect 4525 7973 4537 8007
rect 4571 8004 4583 8007
rect 7558 8004 7564 8016
rect 4571 7976 7564 8004
rect 4571 7973 4583 7976
rect 4525 7967 4583 7973
rect 7558 7964 7564 7976
rect 7616 7964 7622 8016
rect 7650 7964 7656 8016
rect 7708 8004 7714 8016
rect 8113 8007 8171 8013
rect 8113 8004 8125 8007
rect 7708 7976 8125 8004
rect 7708 7964 7714 7976
rect 8113 7973 8125 7976
rect 8159 7973 8171 8007
rect 8113 7967 8171 7973
rect 9944 8007 10002 8013
rect 9944 7973 9956 8007
rect 9990 8004 10002 8007
rect 10042 8004 10048 8016
rect 9990 7976 10048 8004
rect 9990 7973 10002 7976
rect 9944 7967 10002 7973
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 11692 8007 11750 8013
rect 11692 7973 11704 8007
rect 11738 8004 11750 8007
rect 12710 8004 12716 8016
rect 11738 7976 12716 8004
rect 11738 7973 11750 7976
rect 11692 7967 11750 7973
rect 12710 7964 12716 7976
rect 12768 8004 12774 8016
rect 12986 8004 12992 8016
rect 12768 7976 12992 8004
rect 12768 7964 12774 7976
rect 12986 7964 12992 7976
rect 13044 7964 13050 8016
rect 13538 8004 13544 8016
rect 13096 7976 13544 8004
rect 3878 7896 3884 7948
rect 3936 7936 3942 7948
rect 4433 7939 4491 7945
rect 4433 7936 4445 7939
rect 3936 7908 4445 7936
rect 3936 7896 3942 7908
rect 4433 7905 4445 7908
rect 4479 7905 4491 7939
rect 4433 7899 4491 7905
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7936 5687 7939
rect 6270 7936 6276 7948
rect 5675 7908 6276 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 6549 7939 6607 7945
rect 6549 7905 6561 7939
rect 6595 7936 6607 7939
rect 6822 7936 6828 7948
rect 6595 7908 6828 7936
rect 6595 7905 6607 7908
rect 6549 7899 6607 7905
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 7742 7896 7748 7948
rect 7800 7936 7806 7948
rect 8205 7939 8263 7945
rect 8205 7936 8217 7939
rect 7800 7908 8217 7936
rect 7800 7896 7806 7908
rect 8205 7905 8217 7908
rect 8251 7905 8263 7939
rect 8205 7899 8263 7905
rect 11425 7939 11483 7945
rect 11425 7905 11437 7939
rect 11471 7936 11483 7939
rect 12158 7936 12164 7948
rect 11471 7908 12164 7936
rect 11471 7905 11483 7908
rect 11425 7899 11483 7905
rect 12158 7896 12164 7908
rect 12216 7936 12222 7948
rect 13096 7945 13124 7976
rect 13538 7964 13544 7976
rect 13596 7964 13602 8016
rect 13354 7945 13360 7948
rect 13081 7939 13139 7945
rect 13081 7936 13093 7939
rect 12216 7908 13093 7936
rect 12216 7896 12222 7908
rect 13081 7905 13093 7908
rect 13127 7905 13139 7939
rect 13348 7936 13360 7945
rect 13315 7908 13360 7936
rect 13081 7899 13139 7905
rect 13348 7899 13360 7908
rect 13354 7896 13360 7899
rect 13412 7896 13418 7948
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7837 1455 7871
rect 4706 7868 4712 7880
rect 4667 7840 4712 7868
rect 1397 7831 1455 7837
rect 1412 7732 1440 7831
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 5810 7868 5816 7880
rect 5771 7840 5816 7868
rect 5810 7828 5816 7840
rect 5868 7828 5874 7880
rect 5902 7828 5908 7880
rect 5960 7868 5966 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 5960 7840 6745 7868
rect 5960 7828 5966 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 8294 7868 8300 7880
rect 8255 7840 8300 7868
rect 6733 7831 6791 7837
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 8386 7828 8392 7880
rect 8444 7868 8450 7880
rect 8757 7871 8815 7877
rect 8757 7868 8769 7871
rect 8444 7840 8769 7868
rect 8444 7828 8450 7840
rect 8757 7837 8769 7840
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 9674 7828 9680 7880
rect 9732 7868 9738 7880
rect 9732 7840 9777 7868
rect 9732 7828 9738 7840
rect 1670 7732 1676 7744
rect 1412 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 2777 7735 2835 7741
rect 2777 7701 2789 7735
rect 2823 7732 2835 7735
rect 2866 7732 2872 7744
rect 2823 7704 2872 7732
rect 2823 7701 2835 7704
rect 2777 7695 2835 7701
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 5169 7735 5227 7741
rect 5169 7701 5181 7735
rect 5215 7732 5227 7735
rect 10594 7732 10600 7744
rect 5215 7704 10600 7732
rect 5215 7701 5227 7704
rect 5169 7695 5227 7701
rect 10594 7692 10600 7704
rect 10652 7692 10658 7744
rect 10870 7692 10876 7744
rect 10928 7732 10934 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 10928 7704 11069 7732
rect 10928 7692 10934 7704
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11057 7695 11115 7701
rect 12805 7735 12863 7741
rect 12805 7701 12817 7735
rect 12851 7732 12863 7735
rect 13354 7732 13360 7744
rect 12851 7704 13360 7732
rect 12851 7701 12863 7704
rect 12805 7695 12863 7701
rect 13354 7692 13360 7704
rect 13412 7692 13418 7744
rect 14461 7735 14519 7741
rect 14461 7701 14473 7735
rect 14507 7732 14519 7735
rect 14550 7732 14556 7744
rect 14507 7704 14556 7732
rect 14507 7701 14519 7704
rect 14461 7695 14519 7701
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 3513 7531 3571 7537
rect 3513 7497 3525 7531
rect 3559 7528 3571 7531
rect 3786 7528 3792 7540
rect 3559 7500 3792 7528
rect 3559 7497 3571 7500
rect 3513 7491 3571 7497
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 5500 7500 5672 7528
rect 5500 7488 5506 7500
rect 5644 7460 5672 7500
rect 5810 7488 5816 7540
rect 5868 7528 5874 7540
rect 6089 7531 6147 7537
rect 6089 7528 6101 7531
rect 5868 7500 6101 7528
rect 5868 7488 5874 7500
rect 6089 7497 6101 7500
rect 6135 7497 6147 7531
rect 6822 7528 6828 7540
rect 6783 7500 6828 7528
rect 6089 7491 6147 7497
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 10778 7528 10784 7540
rect 10739 7500 10784 7528
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 13262 7528 13268 7540
rect 11440 7500 13268 7528
rect 6365 7463 6423 7469
rect 6365 7460 6377 7463
rect 5644 7432 6377 7460
rect 6365 7429 6377 7432
rect 6411 7429 6423 7463
rect 7745 7463 7803 7469
rect 7745 7460 7757 7463
rect 6365 7423 6423 7429
rect 6656 7432 7757 7460
rect 3970 7392 3976 7404
rect 3931 7364 3976 7392
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 4065 7395 4123 7401
rect 4065 7361 4077 7395
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 1670 7284 1676 7336
rect 1728 7324 1734 7336
rect 1857 7327 1915 7333
rect 1857 7324 1869 7327
rect 1728 7296 1869 7324
rect 1728 7284 1734 7296
rect 1857 7293 1869 7296
rect 1903 7293 1915 7327
rect 1857 7287 1915 7293
rect 2124 7327 2182 7333
rect 2124 7293 2136 7327
rect 2170 7324 2182 7327
rect 2866 7324 2872 7336
rect 2170 7296 2872 7324
rect 2170 7293 2182 7296
rect 2124 7287 2182 7293
rect 2866 7284 2872 7296
rect 2924 7324 2930 7336
rect 4080 7324 4108 7355
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 6656 7392 6684 7432
rect 7745 7429 7757 7432
rect 7791 7429 7803 7463
rect 7745 7423 7803 7429
rect 7837 7463 7895 7469
rect 7837 7429 7849 7463
rect 7883 7460 7895 7463
rect 8478 7460 8484 7472
rect 7883 7432 8484 7460
rect 7883 7429 7895 7432
rect 7837 7423 7895 7429
rect 8478 7420 8484 7432
rect 8536 7420 8542 7472
rect 9769 7463 9827 7469
rect 9769 7429 9781 7463
rect 9815 7460 9827 7463
rect 10689 7463 10747 7469
rect 10689 7460 10701 7463
rect 9815 7432 10701 7460
rect 9815 7429 9827 7432
rect 9769 7423 9827 7429
rect 10689 7429 10701 7432
rect 10735 7429 10747 7463
rect 10689 7423 10747 7429
rect 6052 7364 6684 7392
rect 6052 7352 6058 7364
rect 6730 7352 6736 7404
rect 6788 7392 6794 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 6788 7364 7389 7392
rect 6788 7352 6794 7364
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 8389 7395 8447 7401
rect 8389 7392 8401 7395
rect 7524 7364 8401 7392
rect 7524 7352 7530 7364
rect 8389 7361 8401 7364
rect 8435 7361 8447 7395
rect 8389 7355 8447 7361
rect 10413 7395 10471 7401
rect 10413 7361 10425 7395
rect 10459 7392 10471 7395
rect 10962 7392 10968 7404
rect 10459 7364 10968 7392
rect 10459 7361 10471 7364
rect 10413 7355 10471 7361
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 11440 7401 11468 7500
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 11514 7420 11520 7472
rect 11572 7460 11578 7472
rect 11572 7432 15056 7460
rect 11572 7420 11578 7432
rect 15028 7404 15056 7432
rect 11425 7395 11483 7401
rect 11425 7361 11437 7395
rect 11471 7361 11483 7395
rect 11425 7355 11483 7361
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7392 11943 7395
rect 12066 7392 12072 7404
rect 11931 7364 12072 7392
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 12986 7392 12992 7404
rect 12947 7364 12992 7392
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 13354 7352 13360 7404
rect 13412 7392 13418 7404
rect 14001 7395 14059 7401
rect 14001 7392 14013 7395
rect 13412 7364 14013 7392
rect 13412 7352 13418 7364
rect 14001 7361 14013 7364
rect 14047 7361 14059 7395
rect 15010 7392 15016 7404
rect 14971 7364 15016 7392
rect 14001 7355 14059 7361
rect 15010 7352 15016 7364
rect 15068 7392 15074 7404
rect 16025 7395 16083 7401
rect 16025 7392 16037 7395
rect 15068 7364 16037 7392
rect 15068 7352 15074 7364
rect 16025 7361 16037 7364
rect 16071 7361 16083 7395
rect 16025 7355 16083 7361
rect 2924 7296 4108 7324
rect 4709 7327 4767 7333
rect 2924 7284 2930 7296
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 5442 7324 5448 7336
rect 4755 7296 5448 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 5442 7284 5448 7296
rect 5500 7284 5506 7336
rect 5718 7284 5724 7336
rect 5776 7324 5782 7336
rect 6549 7327 6607 7333
rect 6549 7324 6561 7327
rect 5776 7296 6561 7324
rect 5776 7284 5782 7296
rect 6549 7293 6561 7296
rect 6595 7293 6607 7327
rect 6549 7287 6607 7293
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7285 7327 7343 7333
rect 7285 7324 7297 7327
rect 6972 7296 7297 7324
rect 6972 7284 6978 7296
rect 7285 7293 7297 7296
rect 7331 7293 7343 7327
rect 7285 7287 7343 7293
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7324 7803 7327
rect 8205 7327 8263 7333
rect 8205 7324 8217 7327
rect 7791 7296 8217 7324
rect 7791 7293 7803 7296
rect 7745 7287 7803 7293
rect 8205 7293 8217 7296
rect 8251 7324 8263 7327
rect 8251 7296 9168 7324
rect 8251 7293 8263 7296
rect 8205 7287 8263 7293
rect 2774 7216 2780 7268
rect 2832 7256 2838 7268
rect 3881 7259 3939 7265
rect 3881 7256 3893 7259
rect 2832 7228 3893 7256
rect 2832 7216 2838 7228
rect 3881 7225 3893 7228
rect 3927 7225 3939 7259
rect 3881 7219 3939 7225
rect 4976 7259 5034 7265
rect 4976 7225 4988 7259
rect 5022 7256 5034 7259
rect 5902 7256 5908 7268
rect 5022 7228 5908 7256
rect 5022 7225 5034 7228
rect 4976 7219 5034 7225
rect 5902 7216 5908 7228
rect 5960 7216 5966 7268
rect 8297 7259 8355 7265
rect 8297 7256 8309 7259
rect 6288 7228 8309 7256
rect 3237 7191 3295 7197
rect 3237 7157 3249 7191
rect 3283 7188 3295 7191
rect 3326 7188 3332 7200
rect 3283 7160 3332 7188
rect 3283 7157 3295 7160
rect 3237 7151 3295 7157
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 4062 7148 4068 7200
rect 4120 7188 4126 7200
rect 6288 7188 6316 7228
rect 8297 7225 8309 7228
rect 8343 7256 8355 7259
rect 8570 7256 8576 7268
rect 8343 7228 8576 7256
rect 8343 7225 8355 7228
rect 8297 7219 8355 7225
rect 8570 7216 8576 7228
rect 8628 7216 8634 7268
rect 9140 7256 9168 7296
rect 9214 7284 9220 7336
rect 9272 7324 9278 7336
rect 10137 7327 10195 7333
rect 10137 7324 10149 7327
rect 9272 7296 10149 7324
rect 9272 7284 9278 7296
rect 10137 7293 10149 7296
rect 10183 7293 10195 7327
rect 10137 7287 10195 7293
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 12805 7327 12863 7333
rect 12805 7324 12817 7327
rect 11204 7296 12817 7324
rect 11204 7284 11210 7296
rect 12805 7293 12817 7296
rect 12851 7293 12863 7327
rect 13814 7324 13820 7336
rect 13775 7296 13820 7324
rect 12805 7287 12863 7293
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 14829 7327 14887 7333
rect 14829 7293 14841 7327
rect 14875 7324 14887 7327
rect 16298 7324 16304 7336
rect 14875 7296 16304 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 10042 7256 10048 7268
rect 9140 7228 10048 7256
rect 10042 7216 10048 7228
rect 10100 7216 10106 7268
rect 10689 7259 10747 7265
rect 10689 7225 10701 7259
rect 10735 7256 10747 7259
rect 12250 7256 12256 7268
rect 10735 7228 12256 7256
rect 10735 7225 10747 7228
rect 10689 7219 10747 7225
rect 12250 7216 12256 7228
rect 12308 7216 12314 7268
rect 13909 7259 13967 7265
rect 13909 7256 13921 7259
rect 12452 7228 13921 7256
rect 4120 7160 6316 7188
rect 4120 7148 4126 7160
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 7193 7191 7251 7197
rect 7193 7188 7205 7191
rect 6512 7160 7205 7188
rect 6512 7148 6518 7160
rect 7193 7157 7205 7160
rect 7239 7157 7251 7191
rect 7193 7151 7251 7157
rect 9030 7148 9036 7200
rect 9088 7188 9094 7200
rect 10229 7191 10287 7197
rect 10229 7188 10241 7191
rect 9088 7160 10241 7188
rect 9088 7148 9094 7160
rect 10229 7157 10241 7160
rect 10275 7157 10287 7191
rect 10229 7151 10287 7157
rect 10502 7148 10508 7200
rect 10560 7188 10566 7200
rect 11149 7191 11207 7197
rect 11149 7188 11161 7191
rect 10560 7160 11161 7188
rect 10560 7148 10566 7160
rect 11149 7157 11161 7160
rect 11195 7157 11207 7191
rect 11149 7151 11207 7157
rect 11238 7148 11244 7200
rect 11296 7188 11302 7200
rect 12452 7197 12480 7228
rect 13909 7225 13921 7228
rect 13955 7225 13967 7259
rect 13909 7219 13967 7225
rect 13998 7216 14004 7268
rect 14056 7256 14062 7268
rect 15841 7259 15899 7265
rect 15841 7256 15853 7259
rect 14056 7228 15853 7256
rect 14056 7216 14062 7228
rect 15841 7225 15853 7228
rect 15887 7225 15899 7259
rect 15841 7219 15899 7225
rect 15930 7216 15936 7268
rect 15988 7256 15994 7268
rect 15988 7228 16033 7256
rect 15988 7216 15994 7228
rect 12437 7191 12495 7197
rect 11296 7160 11341 7188
rect 11296 7148 11302 7160
rect 12437 7157 12449 7191
rect 12483 7157 12495 7191
rect 12437 7151 12495 7157
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 12897 7191 12955 7197
rect 12897 7188 12909 7191
rect 12584 7160 12909 7188
rect 12584 7148 12590 7160
rect 12897 7157 12909 7160
rect 12943 7157 12955 7191
rect 12897 7151 12955 7157
rect 13449 7191 13507 7197
rect 13449 7157 13461 7191
rect 13495 7188 13507 7191
rect 14182 7188 14188 7200
rect 13495 7160 14188 7188
rect 13495 7157 13507 7160
rect 13449 7151 13507 7157
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 14458 7188 14464 7200
rect 14419 7160 14464 7188
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 14921 7191 14979 7197
rect 14921 7157 14933 7191
rect 14967 7188 14979 7191
rect 15194 7188 15200 7200
rect 14967 7160 15200 7188
rect 14967 7157 14979 7160
rect 14921 7151 14979 7157
rect 15194 7148 15200 7160
rect 15252 7148 15258 7200
rect 15473 7191 15531 7197
rect 15473 7157 15485 7191
rect 15519 7188 15531 7191
rect 16574 7188 16580 7200
rect 15519 7160 16580 7188
rect 15519 7157 15531 7160
rect 15473 7151 15531 7157
rect 16574 7148 16580 7160
rect 16632 7148 16638 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 3234 6944 3240 6996
rect 3292 6984 3298 6996
rect 3329 6987 3387 6993
rect 3329 6984 3341 6987
rect 3292 6956 3341 6984
rect 3292 6944 3298 6956
rect 3329 6953 3341 6956
rect 3375 6953 3387 6987
rect 3329 6947 3387 6953
rect 4433 6987 4491 6993
rect 4433 6953 4445 6987
rect 4479 6984 4491 6987
rect 5074 6984 5080 6996
rect 4479 6956 5080 6984
rect 4479 6953 4491 6956
rect 4433 6947 4491 6953
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 7285 6987 7343 6993
rect 7285 6953 7297 6987
rect 7331 6984 7343 6987
rect 8202 6984 8208 6996
rect 7331 6956 8208 6984
rect 7331 6953 7343 6956
rect 7285 6947 7343 6953
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 8386 6984 8392 6996
rect 8347 6956 8392 6984
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 10042 6944 10048 6996
rect 10100 6984 10106 6996
rect 11057 6987 11115 6993
rect 11057 6984 11069 6987
rect 10100 6956 11069 6984
rect 10100 6944 10106 6956
rect 11057 6953 11069 6956
rect 11103 6984 11115 6987
rect 11514 6984 11520 6996
rect 11103 6956 11520 6984
rect 11103 6953 11115 6956
rect 11057 6947 11115 6953
rect 11514 6944 11520 6956
rect 11572 6944 11578 6996
rect 11793 6987 11851 6993
rect 11793 6953 11805 6987
rect 11839 6984 11851 6987
rect 11974 6984 11980 6996
rect 11839 6956 11980 6984
rect 11839 6953 11851 6956
rect 11793 6947 11851 6953
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 12437 6987 12495 6993
rect 12437 6953 12449 6987
rect 12483 6984 12495 6987
rect 12526 6984 12532 6996
rect 12483 6956 12532 6984
rect 12483 6953 12495 6956
rect 12437 6947 12495 6953
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 12805 6987 12863 6993
rect 12805 6953 12817 6987
rect 12851 6984 12863 6987
rect 13446 6984 13452 6996
rect 12851 6956 13452 6984
rect 12851 6953 12863 6956
rect 12805 6947 12863 6953
rect 13446 6944 13452 6956
rect 13504 6984 13510 6996
rect 15838 6984 15844 6996
rect 13504 6956 15844 6984
rect 13504 6944 13510 6956
rect 15838 6944 15844 6956
rect 15896 6944 15902 6996
rect 5810 6876 5816 6928
rect 5868 6916 5874 6928
rect 6150 6919 6208 6925
rect 6150 6916 6162 6919
rect 5868 6888 6162 6916
rect 5868 6876 5874 6888
rect 6150 6885 6162 6888
rect 6196 6885 6208 6919
rect 8220 6916 8248 6944
rect 9214 6916 9220 6928
rect 8220 6888 9220 6916
rect 6150 6879 6208 6885
rect 9214 6876 9220 6888
rect 9272 6876 9278 6928
rect 9944 6919 10002 6925
rect 9944 6885 9956 6919
rect 9990 6916 10002 6919
rect 10870 6916 10876 6928
rect 9990 6888 10876 6916
rect 9990 6885 10002 6888
rect 9944 6879 10002 6885
rect 10870 6876 10876 6888
rect 10928 6876 10934 6928
rect 11885 6919 11943 6925
rect 11885 6885 11897 6919
rect 11931 6916 11943 6919
rect 12618 6916 12624 6928
rect 11931 6888 12624 6916
rect 11931 6885 11943 6888
rect 11885 6879 11943 6885
rect 2216 6851 2274 6857
rect 2216 6817 2228 6851
rect 2262 6848 2274 6851
rect 3142 6848 3148 6860
rect 2262 6820 3148 6848
rect 2262 6817 2274 6820
rect 2216 6811 2274 6817
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 5169 6851 5227 6857
rect 5169 6817 5181 6851
rect 5215 6848 5227 6851
rect 6454 6848 6460 6860
rect 5215 6820 6460 6848
rect 5215 6817 5227 6820
rect 5169 6811 5227 6817
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 8478 6848 8484 6860
rect 8439 6820 8484 6848
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 9766 6848 9772 6860
rect 8956 6820 9772 6848
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 1964 6644 1992 6743
rect 2958 6740 2964 6792
rect 3016 6780 3022 6792
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 3016 6752 4537 6780
rect 3016 6740 3022 6752
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 4706 6780 4712 6792
rect 4667 6752 4712 6780
rect 4525 6743 4583 6749
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 5442 6740 5448 6792
rect 5500 6780 5506 6792
rect 5905 6783 5963 6789
rect 5905 6780 5917 6783
rect 5500 6752 5917 6780
rect 5500 6740 5506 6752
rect 5905 6749 5917 6752
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 7116 6752 8248 6780
rect 3786 6672 3792 6724
rect 3844 6712 3850 6724
rect 3844 6684 5948 6712
rect 3844 6672 3850 6684
rect 3694 6644 3700 6656
rect 1964 6616 3700 6644
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 4062 6644 4068 6656
rect 4023 6616 4068 6644
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 5920 6644 5948 6684
rect 7116 6644 7144 6752
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 8021 6715 8079 6721
rect 8021 6712 8033 6715
rect 7248 6684 8033 6712
rect 7248 6672 7254 6684
rect 8021 6681 8033 6684
rect 8067 6681 8079 6715
rect 8220 6712 8248 6752
rect 8294 6740 8300 6792
rect 8352 6780 8358 6792
rect 8573 6783 8631 6789
rect 8573 6780 8585 6783
rect 8352 6752 8585 6780
rect 8352 6740 8358 6752
rect 8573 6749 8585 6752
rect 8619 6749 8631 6783
rect 8573 6743 8631 6749
rect 8956 6712 8984 6820
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 11900 6848 11928 6879
rect 12618 6876 12624 6888
rect 12676 6876 12682 6928
rect 12897 6919 12955 6925
rect 12897 6885 12909 6919
rect 12943 6885 12955 6919
rect 12897 6879 12955 6885
rect 11808 6820 11928 6848
rect 9033 6783 9091 6789
rect 9033 6749 9045 6783
rect 9079 6749 9091 6783
rect 9033 6743 9091 6749
rect 8220 6684 8984 6712
rect 8021 6675 8079 6681
rect 5920 6616 7144 6644
rect 9048 6644 9076 6743
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 9732 6752 9777 6780
rect 9732 6740 9738 6752
rect 10778 6740 10784 6792
rect 10836 6780 10842 6792
rect 11808 6780 11836 6820
rect 10836 6752 11836 6780
rect 10836 6740 10842 6752
rect 12066 6740 12072 6792
rect 12124 6780 12130 6792
rect 12912 6780 12940 6879
rect 13814 6848 13820 6860
rect 13775 6820 13820 6848
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 13906 6808 13912 6860
rect 13964 6848 13970 6860
rect 14737 6851 14795 6857
rect 13964 6820 14009 6848
rect 13964 6808 13970 6820
rect 14737 6817 14749 6851
rect 14783 6848 14795 6851
rect 15657 6851 15715 6857
rect 15657 6848 15669 6851
rect 14783 6820 15669 6848
rect 14783 6817 14795 6820
rect 14737 6811 14795 6817
rect 15657 6817 15669 6820
rect 15703 6817 15715 6851
rect 15657 6811 15715 6817
rect 12986 6780 12992 6792
rect 12124 6752 12169 6780
rect 12912 6752 12992 6780
rect 12124 6740 12130 6752
rect 12986 6740 12992 6752
rect 13044 6740 13050 6792
rect 13081 6783 13139 6789
rect 13081 6749 13093 6783
rect 13127 6780 13139 6783
rect 13354 6780 13360 6792
rect 13127 6752 13360 6780
rect 13127 6749 13139 6752
rect 13081 6743 13139 6749
rect 13354 6740 13360 6752
rect 13412 6740 13418 6792
rect 13998 6780 14004 6792
rect 13959 6752 14004 6780
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 11054 6672 11060 6724
rect 11112 6712 11118 6724
rect 11238 6712 11244 6724
rect 11112 6684 11244 6712
rect 11112 6672 11118 6684
rect 11238 6672 11244 6684
rect 11296 6672 11302 6724
rect 12250 6672 12256 6724
rect 12308 6712 12314 6724
rect 15764 6712 15792 6743
rect 12308 6684 15792 6712
rect 12308 6672 12314 6684
rect 9950 6644 9956 6656
rect 9048 6616 9956 6644
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 11425 6647 11483 6653
rect 11425 6613 11437 6647
rect 11471 6644 11483 6647
rect 11790 6644 11796 6656
rect 11471 6616 11796 6644
rect 11471 6613 11483 6616
rect 11425 6607 11483 6613
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 13170 6604 13176 6656
rect 13228 6644 13234 6656
rect 13449 6647 13507 6653
rect 13449 6644 13461 6647
rect 13228 6616 13461 6644
rect 13228 6604 13234 6616
rect 13449 6613 13461 6616
rect 13495 6613 13507 6647
rect 15286 6644 15292 6656
rect 15247 6616 15292 6644
rect 13449 6607 13507 6613
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 15562 6604 15568 6656
rect 15620 6644 15626 6656
rect 15856 6644 15884 6743
rect 15620 6616 15884 6644
rect 15620 6604 15626 6616
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 3142 6440 3148 6452
rect 3103 6412 3148 6440
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 3970 6400 3976 6452
rect 4028 6440 4034 6452
rect 10778 6440 10784 6452
rect 4028 6412 10784 6440
rect 4028 6400 4034 6412
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 10873 6443 10931 6449
rect 10873 6409 10885 6443
rect 10919 6440 10931 6443
rect 11146 6440 11152 6452
rect 10919 6412 11152 6440
rect 10919 6409 10931 6412
rect 10873 6403 10931 6409
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 11606 6400 11612 6452
rect 11664 6440 11670 6452
rect 13354 6440 13360 6452
rect 11664 6412 13360 6440
rect 11664 6400 11670 6412
rect 13354 6400 13360 6412
rect 13412 6440 13418 6452
rect 13817 6443 13875 6449
rect 13817 6440 13829 6443
rect 13412 6412 13829 6440
rect 13412 6400 13418 6412
rect 13817 6409 13829 6412
rect 13863 6409 13875 6443
rect 13817 6403 13875 6409
rect 10410 6332 10416 6384
rect 10468 6372 10474 6384
rect 10468 6344 12296 6372
rect 10468 6332 10474 6344
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 11333 6307 11391 6313
rect 11333 6304 11345 6307
rect 11204 6276 11345 6304
rect 11204 6264 11210 6276
rect 11333 6273 11345 6276
rect 11379 6273 11391 6307
rect 11333 6267 11391 6273
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6304 11575 6307
rect 11606 6304 11612 6316
rect 11563 6276 11612 6304
rect 11563 6273 11575 6276
rect 11517 6267 11575 6273
rect 11606 6264 11612 6276
rect 11664 6264 11670 6316
rect 1670 6196 1676 6248
rect 1728 6236 1734 6248
rect 1765 6239 1823 6245
rect 1765 6236 1777 6239
rect 1728 6208 1777 6236
rect 1728 6196 1734 6208
rect 1765 6205 1777 6208
rect 1811 6205 1823 6239
rect 1765 6199 1823 6205
rect 3694 6196 3700 6248
rect 3752 6236 3758 6248
rect 4246 6236 4252 6248
rect 3752 6208 4252 6236
rect 3752 6196 3758 6208
rect 4246 6196 4252 6208
rect 4304 6236 4310 6248
rect 4341 6239 4399 6245
rect 4341 6236 4353 6239
rect 4304 6208 4353 6236
rect 4304 6196 4310 6208
rect 4341 6205 4353 6208
rect 4387 6205 4399 6239
rect 4341 6199 4399 6205
rect 4608 6239 4666 6245
rect 4608 6205 4620 6239
rect 4654 6236 4666 6239
rect 6730 6236 6736 6248
rect 4654 6208 6736 6236
rect 4654 6205 4666 6208
rect 4608 6199 4666 6205
rect 6730 6196 6736 6208
rect 6788 6196 6794 6248
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 7561 6239 7619 6245
rect 7561 6236 7573 6239
rect 7156 6208 7573 6236
rect 7156 6196 7162 6208
rect 7561 6205 7573 6208
rect 7607 6205 7619 6239
rect 9030 6236 9036 6248
rect 7561 6199 7619 6205
rect 7760 6208 9036 6236
rect 2032 6171 2090 6177
rect 2032 6137 2044 6171
rect 2078 6168 2090 6171
rect 4706 6168 4712 6180
rect 2078 6140 4712 6168
rect 2078 6137 2090 6140
rect 2032 6131 2090 6137
rect 4706 6128 4712 6140
rect 4764 6128 4770 6180
rect 7760 6168 7788 6208
rect 9030 6196 9036 6208
rect 9088 6196 9094 6248
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6236 9183 6239
rect 9217 6239 9275 6245
rect 9217 6236 9229 6239
rect 9171 6208 9229 6236
rect 9171 6205 9183 6208
rect 9125 6199 9183 6205
rect 9217 6205 9229 6208
rect 9263 6205 9275 6239
rect 9217 6199 9275 6205
rect 9484 6239 9542 6245
rect 9484 6205 9496 6239
rect 9530 6236 9542 6239
rect 10042 6236 10048 6248
rect 9530 6208 10048 6236
rect 9530 6205 9542 6208
rect 9484 6199 9542 6205
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 12268 6245 12296 6344
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 13872 6276 14105 6304
rect 13872 6264 13878 6276
rect 14093 6273 14105 6276
rect 14139 6273 14151 6307
rect 16758 6304 16764 6316
rect 16719 6276 16764 6304
rect 14093 6267 14151 6273
rect 16758 6264 16764 6276
rect 16816 6264 16822 6316
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6205 12311 6239
rect 12253 6199 12311 6205
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6205 12495 6239
rect 12437 6199 12495 6205
rect 5644 6140 7788 6168
rect 7828 6171 7886 6177
rect 3418 6100 3424 6112
rect 3379 6072 3424 6100
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 3602 6060 3608 6112
rect 3660 6100 3666 6112
rect 5644 6100 5672 6140
rect 7828 6137 7840 6171
rect 7874 6168 7886 6171
rect 11422 6168 11428 6180
rect 7874 6140 11428 6168
rect 7874 6137 7886 6140
rect 7828 6131 7886 6137
rect 3660 6072 5672 6100
rect 5721 6103 5779 6109
rect 3660 6060 3666 6072
rect 5721 6069 5733 6103
rect 5767 6100 5779 6103
rect 5810 6100 5816 6112
rect 5767 6072 5816 6100
rect 5767 6069 5779 6072
rect 5721 6063 5779 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 8938 6100 8944 6112
rect 8899 6072 8944 6100
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 9125 6103 9183 6109
rect 9125 6069 9137 6103
rect 9171 6100 9183 6103
rect 9766 6100 9772 6112
rect 9171 6072 9772 6100
rect 9171 6069 9183 6072
rect 9125 6063 9183 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10410 6060 10416 6112
rect 10468 6100 10474 6112
rect 10612 6109 10640 6140
rect 11422 6128 11428 6140
rect 11480 6128 11486 6180
rect 12452 6112 12480 6199
rect 14458 6196 14464 6248
rect 14516 6236 14522 6248
rect 14553 6239 14611 6245
rect 14553 6236 14565 6239
rect 14516 6208 14565 6236
rect 14516 6196 14522 6208
rect 14553 6205 14565 6208
rect 14599 6205 14611 6239
rect 14553 6199 14611 6205
rect 16482 6196 16488 6248
rect 16540 6236 16546 6248
rect 16669 6239 16727 6245
rect 16669 6236 16681 6239
rect 16540 6208 16681 6236
rect 16540 6196 16546 6208
rect 16669 6205 16681 6208
rect 16715 6205 16727 6239
rect 16669 6199 16727 6205
rect 12710 6177 12716 6180
rect 12704 6168 12716 6177
rect 12671 6140 12716 6168
rect 12704 6131 12716 6140
rect 12710 6128 12716 6131
rect 12768 6128 12774 6180
rect 14820 6171 14878 6177
rect 14820 6137 14832 6171
rect 14866 6168 14878 6171
rect 15562 6168 15568 6180
rect 14866 6140 15568 6168
rect 14866 6137 14878 6140
rect 14820 6131 14878 6137
rect 15562 6128 15568 6140
rect 15620 6128 15626 6180
rect 16574 6168 16580 6180
rect 15672 6140 16252 6168
rect 16535 6140 16580 6168
rect 10597 6103 10655 6109
rect 10597 6100 10609 6103
rect 10468 6072 10609 6100
rect 10468 6060 10474 6072
rect 10597 6069 10609 6072
rect 10643 6069 10655 6103
rect 10597 6063 10655 6069
rect 10778 6060 10784 6112
rect 10836 6100 10842 6112
rect 11241 6103 11299 6109
rect 11241 6100 11253 6103
rect 10836 6072 11253 6100
rect 10836 6060 10842 6072
rect 11241 6069 11253 6072
rect 11287 6069 11299 6103
rect 11241 6063 11299 6069
rect 11330 6060 11336 6112
rect 11388 6100 11394 6112
rect 12069 6103 12127 6109
rect 12069 6100 12081 6103
rect 11388 6072 12081 6100
rect 11388 6060 11394 6072
rect 12069 6069 12081 6072
rect 12115 6100 12127 6103
rect 12158 6100 12164 6112
rect 12115 6072 12164 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12158 6060 12164 6072
rect 12216 6100 12222 6112
rect 12434 6100 12440 6112
rect 12216 6072 12440 6100
rect 12216 6060 12222 6072
rect 12434 6060 12440 6072
rect 12492 6060 12498 6112
rect 12618 6060 12624 6112
rect 12676 6100 12682 6112
rect 15672 6100 15700 6140
rect 15930 6100 15936 6112
rect 12676 6072 15700 6100
rect 15891 6072 15936 6100
rect 12676 6060 12682 6072
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 16224 6109 16252 6140
rect 16574 6128 16580 6140
rect 16632 6128 16638 6180
rect 16209 6103 16267 6109
rect 16209 6069 16221 6103
rect 16255 6069 16267 6103
rect 16209 6063 16267 6069
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 2685 5899 2743 5905
rect 2685 5865 2697 5899
rect 2731 5896 2743 5899
rect 3418 5896 3424 5908
rect 2731 5868 3424 5896
rect 2731 5865 2743 5868
rect 2685 5859 2743 5865
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 4356 5868 19012 5896
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5828 2835 5831
rect 4062 5828 4068 5840
rect 2823 5800 4068 5828
rect 2823 5797 2835 5800
rect 2777 5791 2835 5797
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 1854 5720 1860 5772
rect 1912 5760 1918 5772
rect 4356 5760 4384 5868
rect 4706 5788 4712 5840
rect 4764 5828 4770 5840
rect 9674 5828 9680 5840
rect 4764 5800 9680 5828
rect 4764 5788 4770 5800
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 10042 5828 10048 5840
rect 10003 5800 10048 5828
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 10137 5831 10195 5837
rect 10137 5797 10149 5831
rect 10183 5828 10195 5831
rect 10502 5828 10508 5840
rect 10183 5800 10508 5828
rect 10183 5797 10195 5800
rect 10137 5791 10195 5797
rect 10502 5788 10508 5800
rect 10560 5788 10566 5840
rect 10870 5788 10876 5840
rect 10928 5828 10934 5840
rect 10928 5800 12388 5828
rect 10928 5788 10934 5800
rect 1912 5732 4384 5760
rect 4433 5763 4491 5769
rect 1912 5720 1918 5732
rect 4433 5729 4445 5763
rect 4479 5729 4491 5763
rect 4433 5723 4491 5729
rect 4525 5763 4583 5769
rect 4525 5729 4537 5763
rect 4571 5760 4583 5763
rect 5350 5760 5356 5772
rect 4571 5732 5356 5760
rect 4571 5729 4583 5732
rect 4525 5723 4583 5729
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 3142 5692 3148 5704
rect 3007 5664 3148 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 4448 5692 4476 5723
rect 5350 5720 5356 5732
rect 5408 5720 5414 5772
rect 5712 5763 5770 5769
rect 5712 5729 5724 5763
rect 5758 5760 5770 5763
rect 7368 5763 7426 5769
rect 5758 5732 7052 5760
rect 5758 5729 5770 5732
rect 5712 5723 5770 5729
rect 4706 5692 4712 5704
rect 4356 5664 4476 5692
rect 4667 5664 4712 5692
rect 3050 5584 3056 5636
rect 3108 5624 3114 5636
rect 4356 5624 4384 5664
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 5442 5692 5448 5704
rect 5355 5664 5448 5692
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 3108 5596 4384 5624
rect 3108 5584 3114 5596
rect 2314 5556 2320 5568
rect 2275 5528 2320 5556
rect 2314 5516 2320 5528
rect 2372 5516 2378 5568
rect 4062 5556 4068 5568
rect 4023 5528 4068 5556
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 5460 5556 5488 5652
rect 6730 5584 6736 5636
rect 6788 5624 6794 5636
rect 6825 5627 6883 5633
rect 6825 5624 6837 5627
rect 6788 5596 6837 5624
rect 6788 5584 6794 5596
rect 6825 5593 6837 5596
rect 6871 5593 6883 5627
rect 6825 5587 6883 5593
rect 6914 5556 6920 5568
rect 5460 5528 6920 5556
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 7024 5556 7052 5732
rect 7368 5729 7380 5763
rect 7414 5760 7426 5763
rect 8938 5760 8944 5772
rect 7414 5732 8944 5760
rect 7414 5729 7426 5732
rect 7368 5723 7426 5729
rect 8938 5720 8944 5732
rect 8996 5720 9002 5772
rect 9030 5720 9036 5772
rect 9088 5760 9094 5772
rect 10778 5760 10784 5772
rect 9088 5732 10784 5760
rect 9088 5720 9094 5732
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 11238 5760 11244 5772
rect 11199 5732 11244 5760
rect 11238 5720 11244 5732
rect 11296 5720 11302 5772
rect 11497 5763 11555 5769
rect 11497 5760 11509 5763
rect 11348 5732 11509 5760
rect 7098 5652 7104 5704
rect 7156 5692 7162 5704
rect 10321 5695 10379 5701
rect 7156 5664 7201 5692
rect 7156 5652 7162 5664
rect 10321 5661 10333 5695
rect 10367 5692 10379 5695
rect 10410 5692 10416 5704
rect 10367 5664 10416 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 11348 5692 11376 5732
rect 11497 5729 11509 5732
rect 11543 5760 11555 5763
rect 12066 5760 12072 5772
rect 11543 5732 12072 5760
rect 11543 5729 11555 5732
rect 11497 5723 11555 5729
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 10928 5664 11376 5692
rect 12360 5692 12388 5800
rect 12434 5788 12440 5840
rect 12492 5828 12498 5840
rect 14458 5828 14464 5840
rect 12492 5800 14464 5828
rect 12492 5788 12498 5800
rect 12897 5763 12955 5769
rect 12897 5729 12909 5763
rect 12943 5760 12955 5763
rect 13170 5760 13176 5772
rect 12943 5732 13176 5760
rect 12943 5729 12955 5732
rect 12897 5723 12955 5729
rect 13170 5720 13176 5732
rect 13228 5720 13234 5772
rect 13556 5769 13584 5800
rect 14458 5788 14464 5800
rect 14516 5828 14522 5840
rect 14516 5800 15332 5828
rect 14516 5788 14522 5800
rect 13814 5769 13820 5772
rect 13541 5763 13599 5769
rect 13541 5729 13553 5763
rect 13587 5729 13599 5763
rect 13808 5760 13820 5769
rect 13775 5732 13820 5760
rect 13541 5723 13599 5729
rect 13808 5723 13820 5732
rect 13814 5720 13820 5723
rect 13872 5720 13878 5772
rect 15304 5769 15332 5800
rect 15470 5788 15476 5840
rect 15528 5788 15534 5840
rect 16022 5788 16028 5840
rect 16080 5828 16086 5840
rect 16080 5800 17172 5828
rect 16080 5788 16086 5800
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5729 15347 5763
rect 15488 5760 15516 5788
rect 15556 5763 15614 5769
rect 15556 5760 15568 5763
rect 15488 5732 15568 5760
rect 15289 5723 15347 5729
rect 15556 5729 15568 5732
rect 15602 5760 15614 5763
rect 15930 5760 15936 5772
rect 15602 5732 15936 5760
rect 15602 5729 15614 5732
rect 15556 5723 15614 5729
rect 15930 5720 15936 5732
rect 15988 5720 15994 5772
rect 17144 5769 17172 5800
rect 18984 5769 19012 5868
rect 17129 5763 17187 5769
rect 17129 5729 17141 5763
rect 17175 5729 17187 5763
rect 17129 5723 17187 5729
rect 18969 5763 19027 5769
rect 18969 5729 18981 5763
rect 19015 5729 19027 5763
rect 18969 5723 19027 5729
rect 13354 5692 13360 5704
rect 12360 5664 13360 5692
rect 10928 5652 10934 5664
rect 13354 5652 13360 5664
rect 13412 5652 13418 5704
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5692 17463 5695
rect 17954 5692 17960 5704
rect 17451 5664 17960 5692
rect 17451 5661 17463 5664
rect 17405 5655 17463 5661
rect 17954 5652 17960 5664
rect 18012 5652 18018 5704
rect 19245 5695 19303 5701
rect 19245 5661 19257 5695
rect 19291 5692 19303 5695
rect 19794 5692 19800 5704
rect 19291 5664 19800 5692
rect 19291 5661 19303 5664
rect 19245 5655 19303 5661
rect 19794 5652 19800 5664
rect 19852 5652 19858 5704
rect 16390 5584 16396 5636
rect 16448 5624 16454 5636
rect 16669 5627 16727 5633
rect 16669 5624 16681 5627
rect 16448 5596 16681 5624
rect 16448 5584 16454 5596
rect 16669 5593 16681 5596
rect 16715 5593 16727 5627
rect 16669 5587 16727 5593
rect 8202 5556 8208 5568
rect 7024 5528 8208 5556
rect 8202 5516 8208 5528
rect 8260 5556 8266 5568
rect 8481 5559 8539 5565
rect 8481 5556 8493 5559
rect 8260 5528 8493 5556
rect 8260 5516 8266 5528
rect 8481 5525 8493 5528
rect 8527 5525 8539 5559
rect 9674 5556 9680 5568
rect 9635 5528 9680 5556
rect 8481 5519 8539 5525
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 10042 5516 10048 5568
rect 10100 5556 10106 5568
rect 11974 5556 11980 5568
rect 10100 5528 11980 5556
rect 10100 5516 10106 5528
rect 11974 5516 11980 5528
rect 12032 5516 12038 5568
rect 12526 5516 12532 5568
rect 12584 5556 12590 5568
rect 12621 5559 12679 5565
rect 12621 5556 12633 5559
rect 12584 5528 12633 5556
rect 12584 5516 12590 5528
rect 12621 5525 12633 5528
rect 12667 5525 12679 5559
rect 12621 5519 12679 5525
rect 13081 5559 13139 5565
rect 13081 5525 13093 5559
rect 13127 5556 13139 5559
rect 13538 5556 13544 5568
rect 13127 5528 13544 5556
rect 13127 5525 13139 5528
rect 13081 5519 13139 5525
rect 13538 5516 13544 5528
rect 13596 5516 13602 5568
rect 14921 5559 14979 5565
rect 14921 5525 14933 5559
rect 14967 5556 14979 5559
rect 15562 5556 15568 5568
rect 14967 5528 15568 5556
rect 14967 5525 14979 5528
rect 14921 5519 14979 5525
rect 15562 5516 15568 5528
rect 15620 5516 15626 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 1854 5352 1860 5364
rect 1815 5324 1860 5352
rect 1854 5312 1860 5324
rect 1912 5312 1918 5364
rect 3234 5352 3240 5364
rect 2424 5324 3240 5352
rect 2424 5225 2452 5324
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 3786 5312 3792 5364
rect 3844 5352 3850 5364
rect 6178 5352 6184 5364
rect 3844 5324 6040 5352
rect 6139 5324 6184 5352
rect 3844 5312 3850 5324
rect 6012 5284 6040 5324
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 6270 5312 6276 5364
rect 6328 5352 6334 5364
rect 6825 5355 6883 5361
rect 6825 5352 6837 5355
rect 6328 5324 6837 5352
rect 6328 5312 6334 5324
rect 6825 5321 6837 5324
rect 6871 5321 6883 5355
rect 7374 5352 7380 5364
rect 6825 5315 6883 5321
rect 7300 5324 7380 5352
rect 7300 5284 7328 5324
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 12618 5352 12624 5364
rect 8680 5324 12624 5352
rect 6012 5256 7328 5284
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5185 2467 5219
rect 2409 5179 2467 5185
rect 3142 5176 3148 5228
rect 3200 5216 3206 5228
rect 3421 5219 3479 5225
rect 3421 5216 3433 5219
rect 3200 5188 3433 5216
rect 3200 5176 3206 5188
rect 3421 5185 3433 5188
rect 3467 5185 3479 5219
rect 3421 5179 3479 5185
rect 5810 5176 5816 5228
rect 5868 5216 5874 5228
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 5868 5188 7389 5216
rect 5868 5176 5874 5188
rect 7377 5185 7389 5188
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 2225 5151 2283 5157
rect 2225 5117 2237 5151
rect 2271 5148 2283 5151
rect 2314 5148 2320 5160
rect 2271 5120 2320 5148
rect 2271 5117 2283 5120
rect 2225 5111 2283 5117
rect 2314 5108 2320 5120
rect 2372 5108 2378 5160
rect 3237 5151 3295 5157
rect 3237 5117 3249 5151
rect 3283 5148 3295 5151
rect 4062 5148 4068 5160
rect 3283 5120 4068 5148
rect 3283 5117 3295 5120
rect 3237 5111 3295 5117
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 4246 5108 4252 5160
rect 4304 5148 4310 5160
rect 4614 5148 4620 5160
rect 4304 5120 4620 5148
rect 4304 5108 4310 5120
rect 4614 5108 4620 5120
rect 4672 5148 4678 5160
rect 4801 5151 4859 5157
rect 4801 5148 4813 5151
rect 4672 5120 4813 5148
rect 4672 5108 4678 5120
rect 4801 5117 4813 5120
rect 4847 5148 4859 5151
rect 5442 5148 5448 5160
rect 4847 5120 5448 5148
rect 4847 5117 4859 5120
rect 4801 5111 4859 5117
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 5534 5108 5540 5160
rect 5592 5148 5598 5160
rect 8680 5157 8708 5324
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 12710 5312 12716 5364
rect 12768 5352 12774 5364
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 12768 5324 13829 5352
rect 12768 5312 12774 5324
rect 13817 5321 13829 5324
rect 13863 5321 13875 5355
rect 13817 5315 13875 5321
rect 13906 5312 13912 5364
rect 13964 5352 13970 5364
rect 14550 5352 14556 5364
rect 13964 5324 14556 5352
rect 13964 5312 13970 5324
rect 14550 5312 14556 5324
rect 14608 5352 14614 5364
rect 14734 5352 14740 5364
rect 14608 5324 14740 5352
rect 14608 5312 14614 5324
rect 14734 5312 14740 5324
rect 14792 5312 14798 5364
rect 14829 5355 14887 5361
rect 14829 5321 14841 5355
rect 14875 5352 14887 5355
rect 16022 5352 16028 5364
rect 14875 5324 16028 5352
rect 14875 5321 14887 5324
rect 14829 5315 14887 5321
rect 16022 5312 16028 5324
rect 16080 5312 16086 5364
rect 11333 5287 11391 5293
rect 11333 5253 11345 5287
rect 11379 5253 11391 5287
rect 11333 5247 11391 5253
rect 8938 5216 8944 5228
rect 8899 5188 8944 5216
rect 8938 5176 8944 5188
rect 8996 5176 9002 5228
rect 9582 5176 9588 5228
rect 9640 5216 9646 5228
rect 10505 5219 10563 5225
rect 10505 5216 10517 5219
rect 9640 5188 10517 5216
rect 9640 5176 9646 5188
rect 10505 5185 10517 5188
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5216 10747 5219
rect 10962 5216 10968 5228
rect 10735 5188 10968 5216
rect 10735 5185 10747 5188
rect 10689 5179 10747 5185
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 7193 5151 7251 5157
rect 7193 5148 7205 5151
rect 5592 5120 7205 5148
rect 5592 5108 5598 5120
rect 7193 5117 7205 5120
rect 7239 5117 7251 5151
rect 7193 5111 7251 5117
rect 8665 5151 8723 5157
rect 8665 5117 8677 5151
rect 8711 5117 8723 5151
rect 8665 5111 8723 5117
rect 8757 5151 8815 5157
rect 8757 5117 8769 5151
rect 8803 5148 8815 5151
rect 9674 5148 9680 5160
rect 8803 5120 9680 5148
rect 8803 5117 8815 5120
rect 8757 5111 8815 5117
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 11348 5148 11376 5247
rect 12250 5244 12256 5296
rect 12308 5284 12314 5296
rect 12434 5284 12440 5296
rect 12308 5256 12440 5284
rect 12308 5244 12314 5256
rect 12434 5244 12440 5256
rect 12492 5244 12498 5296
rect 13446 5244 13452 5296
rect 13504 5284 13510 5296
rect 13504 5256 17264 5284
rect 13504 5244 13510 5256
rect 11790 5216 11796 5228
rect 11751 5188 11796 5216
rect 11790 5176 11796 5188
rect 11848 5176 11854 5228
rect 11882 5176 11888 5228
rect 11940 5216 11946 5228
rect 11977 5219 12035 5225
rect 11977 5216 11989 5219
rect 11940 5188 11989 5216
rect 11940 5176 11946 5188
rect 11977 5185 11989 5188
rect 12023 5216 12035 5219
rect 14461 5219 14519 5225
rect 14461 5216 14473 5219
rect 12023 5188 12572 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 12544 5160 12572 5188
rect 13924 5188 14473 5216
rect 12434 5148 12440 5160
rect 11348 5120 12304 5148
rect 12395 5120 12440 5148
rect 4154 5080 4160 5092
rect 3252 5052 4160 5080
rect 3252 5024 3280 5052
rect 4154 5040 4160 5052
rect 4212 5040 4218 5092
rect 5068 5083 5126 5089
rect 5068 5049 5080 5083
rect 5114 5080 5126 5083
rect 5994 5080 6000 5092
rect 5114 5052 6000 5080
rect 5114 5049 5126 5052
rect 5068 5043 5126 5049
rect 5994 5040 6000 5052
rect 6052 5040 6058 5092
rect 6546 5040 6552 5092
rect 6604 5080 6610 5092
rect 7285 5083 7343 5089
rect 7285 5080 7297 5083
rect 6604 5052 7297 5080
rect 6604 5040 6610 5052
rect 7285 5049 7297 5052
rect 7331 5049 7343 5083
rect 11606 5080 11612 5092
rect 7285 5043 7343 5049
rect 8312 5052 11612 5080
rect 2317 5015 2375 5021
rect 2317 4981 2329 5015
rect 2363 5012 2375 5015
rect 2869 5015 2927 5021
rect 2869 5012 2881 5015
rect 2363 4984 2881 5012
rect 2363 4981 2375 4984
rect 2317 4975 2375 4981
rect 2869 4981 2881 4984
rect 2915 4981 2927 5015
rect 2869 4975 2927 4981
rect 3234 4972 3240 5024
rect 3292 4972 3298 5024
rect 3329 5015 3387 5021
rect 3329 4981 3341 5015
rect 3375 5012 3387 5015
rect 4062 5012 4068 5024
rect 3375 4984 4068 5012
rect 3375 4981 3387 4984
rect 3329 4975 3387 4981
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 8312 5021 8340 5052
rect 11606 5040 11612 5052
rect 11664 5040 11670 5092
rect 11701 5083 11759 5089
rect 11701 5049 11713 5083
rect 11747 5080 11759 5083
rect 12276 5080 12304 5120
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 12526 5108 12532 5160
rect 12584 5148 12590 5160
rect 13924 5157 13952 5188
rect 14461 5185 14473 5188
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 14734 5176 14740 5228
rect 14792 5216 14798 5228
rect 14792 5188 15424 5216
rect 14792 5176 14798 5188
rect 12693 5151 12751 5157
rect 12693 5148 12705 5151
rect 12584 5120 12705 5148
rect 12584 5108 12590 5120
rect 12693 5117 12705 5120
rect 12739 5117 12751 5151
rect 12693 5111 12751 5117
rect 13909 5151 13967 5157
rect 13909 5117 13921 5151
rect 13955 5117 13967 5151
rect 14274 5148 14280 5160
rect 14235 5120 14280 5148
rect 13909 5111 13967 5117
rect 14274 5108 14280 5120
rect 14332 5108 14338 5160
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5148 15255 5151
rect 15286 5148 15292 5160
rect 15243 5120 15292 5148
rect 15243 5117 15255 5120
rect 15197 5111 15255 5117
rect 15286 5108 15292 5120
rect 15344 5108 15350 5160
rect 15396 5148 15424 5188
rect 15470 5176 15476 5228
rect 15528 5216 15534 5228
rect 15528 5188 15573 5216
rect 15528 5176 15534 5188
rect 15746 5176 15752 5228
rect 15804 5216 15810 5228
rect 16114 5216 16120 5228
rect 15804 5188 16120 5216
rect 15804 5176 15810 5188
rect 16114 5176 16120 5188
rect 16172 5216 16178 5228
rect 16301 5219 16359 5225
rect 16301 5216 16313 5219
rect 16172 5188 16313 5216
rect 16172 5176 16178 5188
rect 16301 5185 16313 5188
rect 16347 5185 16359 5219
rect 16301 5179 16359 5185
rect 16393 5219 16451 5225
rect 16393 5185 16405 5219
rect 16439 5185 16451 5219
rect 16393 5179 16451 5185
rect 16408 5148 16436 5179
rect 17236 5157 17264 5256
rect 17402 5216 17408 5228
rect 17363 5188 17408 5216
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 15396 5120 16436 5148
rect 17221 5151 17279 5157
rect 17221 5117 17233 5151
rect 17267 5117 17279 5151
rect 19794 5148 19800 5160
rect 19755 5120 19800 5148
rect 17221 5111 17279 5117
rect 19794 5108 19800 5120
rect 19852 5108 19858 5160
rect 12986 5080 12992 5092
rect 11747 5052 12204 5080
rect 12276 5052 12992 5080
rect 11747 5049 11759 5052
rect 11701 5043 11759 5049
rect 8297 5015 8355 5021
rect 8297 4981 8309 5015
rect 8343 4981 8355 5015
rect 10042 5012 10048 5024
rect 10003 4984 10048 5012
rect 8297 4975 8355 4981
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 10134 4972 10140 5024
rect 10192 5012 10198 5024
rect 10413 5015 10471 5021
rect 10413 5012 10425 5015
rect 10192 4984 10425 5012
rect 10192 4972 10198 4984
rect 10413 4981 10425 4984
rect 10459 5012 10471 5015
rect 12066 5012 12072 5024
rect 10459 4984 12072 5012
rect 10459 4981 10471 4984
rect 10413 4975 10471 4981
rect 12066 4972 12072 4984
rect 12124 4972 12130 5024
rect 12176 5012 12204 5052
rect 12986 5040 12992 5052
rect 13044 5040 13050 5092
rect 13446 5040 13452 5092
rect 13504 5080 13510 5092
rect 17313 5083 17371 5089
rect 17313 5080 17325 5083
rect 13504 5052 17325 5080
rect 13504 5040 13510 5052
rect 17313 5049 17325 5052
rect 17359 5049 17371 5083
rect 17313 5043 17371 5049
rect 12434 5012 12440 5024
rect 12176 4984 12440 5012
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 13998 5012 14004 5024
rect 12584 4984 14004 5012
rect 12584 4972 12590 4984
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 14093 5015 14151 5021
rect 14093 4981 14105 5015
rect 14139 5012 14151 5015
rect 15010 5012 15016 5024
rect 14139 4984 15016 5012
rect 14139 4981 14151 4984
rect 14093 4975 14151 4981
rect 15010 4972 15016 4984
rect 15068 4972 15074 5024
rect 15286 4972 15292 5024
rect 15344 5012 15350 5024
rect 15344 4984 15389 5012
rect 15344 4972 15350 4984
rect 15746 4972 15752 5024
rect 15804 5012 15810 5024
rect 15841 5015 15899 5021
rect 15841 5012 15853 5015
rect 15804 4984 15853 5012
rect 15804 4972 15810 4984
rect 15841 4981 15853 4984
rect 15887 4981 15899 5015
rect 15841 4975 15899 4981
rect 16022 4972 16028 5024
rect 16080 5012 16086 5024
rect 16209 5015 16267 5021
rect 16209 5012 16221 5015
rect 16080 4984 16221 5012
rect 16080 4972 16086 4984
rect 16209 4981 16221 4984
rect 16255 4981 16267 5015
rect 16850 5012 16856 5024
rect 16811 4984 16856 5012
rect 16209 4975 16267 4981
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 19981 5015 20039 5021
rect 19981 4981 19993 5015
rect 20027 5012 20039 5015
rect 20622 5012 20628 5024
rect 20027 4984 20628 5012
rect 20027 4981 20039 4984
rect 19981 4975 20039 4981
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 4062 4808 4068 4820
rect 4023 4780 4068 4808
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 4798 4768 4804 4820
rect 4856 4808 4862 4820
rect 5258 4808 5264 4820
rect 4856 4780 5264 4808
rect 4856 4768 4862 4780
rect 5258 4768 5264 4780
rect 5316 4768 5322 4820
rect 5534 4808 5540 4820
rect 5495 4780 5540 4808
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 6546 4808 6552 4820
rect 6507 4780 6552 4808
rect 6546 4768 6552 4780
rect 6604 4768 6610 4820
rect 7009 4811 7067 4817
rect 7009 4777 7021 4811
rect 7055 4808 7067 4811
rect 7561 4811 7619 4817
rect 7561 4808 7573 4811
rect 7055 4780 7573 4808
rect 7055 4777 7067 4780
rect 7009 4771 7067 4777
rect 7561 4777 7573 4780
rect 7607 4777 7619 4811
rect 7561 4771 7619 4777
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 10134 4808 10140 4820
rect 7708 4780 10140 4808
rect 7708 4768 7714 4780
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 10229 4811 10287 4817
rect 10229 4777 10241 4811
rect 10275 4808 10287 4811
rect 11609 4811 11667 4817
rect 11609 4808 11621 4811
rect 10275 4780 11621 4808
rect 10275 4777 10287 4780
rect 10229 4771 10287 4777
rect 11609 4777 11621 4780
rect 11655 4777 11667 4811
rect 11609 4771 11667 4777
rect 11701 4811 11759 4817
rect 11701 4777 11713 4811
rect 11747 4808 11759 4811
rect 12526 4808 12532 4820
rect 11747 4780 12532 4808
rect 11747 4777 11759 4780
rect 11701 4771 11759 4777
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 13906 4808 13912 4820
rect 12676 4780 13912 4808
rect 12676 4768 12682 4780
rect 13906 4768 13912 4780
rect 13964 4768 13970 4820
rect 14366 4768 14372 4820
rect 14424 4808 14430 4820
rect 15286 4808 15292 4820
rect 14424 4780 15148 4808
rect 15247 4780 15292 4808
rect 14424 4768 14430 4780
rect 3970 4700 3976 4752
rect 4028 4740 4034 4752
rect 4028 4712 4844 4740
rect 4028 4700 4034 4712
rect 1581 4675 1639 4681
rect 1581 4641 1593 4675
rect 1627 4672 1639 4675
rect 1670 4672 1676 4684
rect 1627 4644 1676 4672
rect 1627 4641 1639 4644
rect 1581 4635 1639 4641
rect 1670 4632 1676 4644
rect 1728 4632 1734 4684
rect 1848 4675 1906 4681
rect 1848 4641 1860 4675
rect 1894 4672 1906 4675
rect 2774 4672 2780 4684
rect 1894 4644 2780 4672
rect 1894 4641 1906 4644
rect 1848 4635 1906 4641
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 3142 4632 3148 4684
rect 3200 4672 3206 4684
rect 4154 4672 4160 4684
rect 3200 4644 4160 4672
rect 3200 4632 3206 4644
rect 4154 4632 4160 4644
rect 4212 4672 4218 4684
rect 4433 4675 4491 4681
rect 4433 4672 4445 4675
rect 4212 4644 4445 4672
rect 4212 4632 4218 4644
rect 4433 4641 4445 4644
rect 4479 4641 4491 4675
rect 4816 4672 4844 4712
rect 4890 4700 4896 4752
rect 4948 4740 4954 4752
rect 5350 4740 5356 4752
rect 4948 4712 5356 4740
rect 4948 4700 4954 4712
rect 5350 4700 5356 4712
rect 5408 4740 5414 4752
rect 5905 4743 5963 4749
rect 5905 4740 5917 4743
rect 5408 4712 5917 4740
rect 5408 4700 5414 4712
rect 5905 4709 5917 4712
rect 5951 4709 5963 4743
rect 8941 4743 8999 4749
rect 8941 4740 8953 4743
rect 5905 4703 5963 4709
rect 6748 4712 8953 4740
rect 6748 4672 6776 4712
rect 8941 4709 8953 4712
rect 8987 4740 8999 4743
rect 9493 4743 9551 4749
rect 9493 4740 9505 4743
rect 8987 4712 9505 4740
rect 8987 4709 8999 4712
rect 8941 4703 8999 4709
rect 9493 4709 9505 4712
rect 9539 4709 9551 4743
rect 9766 4740 9772 4752
rect 9727 4712 9772 4740
rect 9493 4703 9551 4709
rect 9766 4700 9772 4712
rect 9824 4700 9830 4752
rect 10042 4700 10048 4752
rect 10100 4740 10106 4752
rect 15120 4740 15148 4780
rect 15286 4768 15292 4780
rect 15344 4768 15350 4820
rect 15746 4808 15752 4820
rect 15707 4780 15752 4808
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 16298 4808 16304 4820
rect 16259 4780 16304 4808
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 16758 4740 16764 4752
rect 10100 4712 13400 4740
rect 10100 4700 10106 4712
rect 6914 4672 6920 4684
rect 4816 4644 6776 4672
rect 6875 4644 6920 4672
rect 4433 4635 4491 4641
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 7929 4675 7987 4681
rect 7929 4641 7941 4675
rect 7975 4672 7987 4675
rect 8662 4672 8668 4684
rect 7975 4644 8668 4672
rect 7975 4641 7987 4644
rect 7929 4635 7987 4641
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 9033 4675 9091 4681
rect 9033 4641 9045 4675
rect 9079 4672 9091 4675
rect 9306 4672 9312 4684
rect 9079 4644 9312 4672
rect 9079 4641 9091 4644
rect 9033 4635 9091 4641
rect 9306 4632 9312 4644
rect 9364 4672 9370 4684
rect 10597 4675 10655 4681
rect 10597 4672 10609 4675
rect 9364 4644 10609 4672
rect 9364 4632 9370 4644
rect 10597 4641 10609 4644
rect 10643 4641 10655 4675
rect 10597 4635 10655 4641
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4672 10747 4675
rect 10962 4672 10968 4684
rect 10735 4644 10968 4672
rect 10735 4641 10747 4644
rect 10689 4635 10747 4641
rect 3329 4607 3387 4613
rect 3329 4573 3341 4607
rect 3375 4604 3387 4607
rect 3418 4604 3424 4616
rect 3375 4576 3424 4604
rect 3375 4573 3387 4576
rect 3329 4567 3387 4573
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 4525 4607 4583 4613
rect 4525 4573 4537 4607
rect 4571 4573 4583 4607
rect 4706 4604 4712 4616
rect 4667 4576 4712 4604
rect 4525 4567 4583 4573
rect 2958 4468 2964 4480
rect 2919 4440 2964 4468
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 4540 4468 4568 4567
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4604 6055 4607
rect 6086 4604 6092 4616
rect 6043 4576 6092 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 6086 4564 6092 4576
rect 6144 4564 6150 4616
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4604 6239 4607
rect 6730 4604 6736 4616
rect 6227 4576 6736 4604
rect 6227 4573 6239 4576
rect 6181 4567 6239 4573
rect 6730 4564 6736 4576
rect 6788 4604 6794 4616
rect 7101 4607 7159 4613
rect 7101 4604 7113 4607
rect 6788 4576 7113 4604
rect 6788 4564 6794 4576
rect 7101 4573 7113 4576
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 7558 4564 7564 4616
rect 7616 4604 7622 4616
rect 8021 4607 8079 4613
rect 8021 4604 8033 4607
rect 7616 4576 8033 4604
rect 7616 4564 7622 4576
rect 8021 4573 8033 4576
rect 8067 4573 8079 4607
rect 8202 4604 8208 4616
rect 8163 4576 8208 4604
rect 8021 4567 8079 4573
rect 8036 4536 8064 4567
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 9214 4604 9220 4616
rect 8352 4576 8708 4604
rect 9175 4576 9220 4604
rect 8352 4564 8358 4576
rect 8478 4536 8484 4548
rect 8036 4508 8484 4536
rect 8478 4496 8484 4508
rect 8536 4496 8542 4548
rect 8386 4468 8392 4480
rect 4540 4440 8392 4468
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 8570 4468 8576 4480
rect 8531 4440 8576 4468
rect 8570 4428 8576 4440
rect 8628 4428 8634 4480
rect 8680 4468 8708 4576
rect 9214 4564 9220 4576
rect 9272 4604 9278 4616
rect 9950 4604 9956 4616
rect 9272 4576 9956 4604
rect 9272 4564 9278 4576
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 10042 4564 10048 4616
rect 10100 4604 10106 4616
rect 10704 4604 10732 4635
rect 10962 4632 10968 4644
rect 11020 4632 11026 4684
rect 11716 4644 12204 4672
rect 10870 4604 10876 4616
rect 10100 4576 10732 4604
rect 10831 4576 10876 4604
rect 10100 4564 10106 4576
rect 10870 4564 10876 4576
rect 10928 4604 10934 4616
rect 11716 4604 11744 4644
rect 11882 4604 11888 4616
rect 10928 4576 11744 4604
rect 11843 4576 11888 4604
rect 10928 4564 10934 4576
rect 11882 4564 11888 4576
rect 11940 4564 11946 4616
rect 12176 4604 12204 4644
rect 12250 4632 12256 4684
rect 12308 4672 12314 4684
rect 12529 4675 12587 4681
rect 12529 4672 12541 4675
rect 12308 4644 12541 4672
rect 12308 4632 12314 4644
rect 12529 4641 12541 4644
rect 12575 4641 12587 4675
rect 12529 4635 12587 4641
rect 12618 4632 12624 4684
rect 12676 4632 12682 4684
rect 12796 4675 12854 4681
rect 12796 4641 12808 4675
rect 12842 4672 12854 4675
rect 13078 4672 13084 4684
rect 12842 4644 13084 4672
rect 12842 4641 12854 4644
rect 12796 4635 12854 4641
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13372 4672 13400 4712
rect 14476 4712 14688 4740
rect 15120 4712 16764 4740
rect 14476 4672 14504 4712
rect 13372 4644 14504 4672
rect 14660 4672 14688 4712
rect 16758 4700 16764 4712
rect 16816 4700 16822 4752
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 14660 4644 15669 4672
rect 15657 4641 15669 4644
rect 15703 4641 15715 4675
rect 15657 4635 15715 4641
rect 16022 4632 16028 4684
rect 16080 4672 16086 4684
rect 16669 4675 16727 4681
rect 16669 4672 16681 4675
rect 16080 4644 16681 4672
rect 16080 4632 16086 4644
rect 16669 4641 16681 4644
rect 16715 4641 16727 4675
rect 17954 4672 17960 4684
rect 17915 4644 17960 4672
rect 16669 4635 16727 4641
rect 17954 4632 17960 4644
rect 18012 4632 18018 4684
rect 12636 4604 12664 4632
rect 14458 4604 14464 4616
rect 12176 4576 12664 4604
rect 13832 4576 14228 4604
rect 14419 4576 14464 4604
rect 9493 4539 9551 4545
rect 9493 4505 9505 4539
rect 9539 4536 9551 4539
rect 11054 4536 11060 4548
rect 9539 4508 11060 4536
rect 9539 4505 9551 4508
rect 9493 4499 9551 4505
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 11790 4536 11796 4548
rect 11164 4508 11796 4536
rect 9582 4468 9588 4480
rect 8680 4440 9588 4468
rect 9582 4428 9588 4440
rect 9640 4468 9646 4480
rect 11164 4468 11192 4508
rect 11790 4496 11796 4508
rect 11848 4496 11854 4548
rect 9640 4440 11192 4468
rect 11241 4471 11299 4477
rect 9640 4428 9646 4440
rect 11241 4437 11253 4471
rect 11287 4468 11299 4471
rect 12526 4468 12532 4480
rect 11287 4440 12532 4468
rect 11287 4437 11299 4440
rect 11241 4431 11299 4437
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 12894 4428 12900 4480
rect 12952 4468 12958 4480
rect 13832 4468 13860 4576
rect 13998 4536 14004 4548
rect 13959 4508 14004 4536
rect 13998 4496 14004 4508
rect 14056 4496 14062 4548
rect 12952 4440 13860 4468
rect 14200 4468 14228 4576
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 14642 4604 14648 4616
rect 14603 4576 14648 4604
rect 14642 4564 14648 4576
rect 14700 4564 14706 4616
rect 15562 4564 15568 4616
rect 15620 4604 15626 4616
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 15620 4576 15853 4604
rect 15620 4564 15626 4576
rect 15841 4573 15853 4576
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 15930 4564 15936 4616
rect 15988 4604 15994 4616
rect 16853 4607 16911 4613
rect 16853 4604 16865 4607
rect 15988 4576 16865 4604
rect 15988 4564 15994 4576
rect 16853 4573 16865 4576
rect 16899 4604 16911 4607
rect 17402 4604 17408 4616
rect 16899 4576 17408 4604
rect 16899 4573 16911 4576
rect 16853 4567 16911 4573
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 14366 4468 14372 4480
rect 14200 4440 14372 4468
rect 12952 4428 12958 4440
rect 14366 4428 14372 4440
rect 14424 4428 14430 4480
rect 18141 4471 18199 4477
rect 18141 4437 18153 4471
rect 18187 4468 18199 4471
rect 18782 4468 18788 4480
rect 18187 4440 18788 4468
rect 18187 4437 18199 4440
rect 18141 4431 18199 4437
rect 18782 4428 18788 4440
rect 18840 4428 18846 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 6825 4267 6883 4273
rect 3804 4236 5672 4264
rect 1670 4088 1676 4140
rect 1728 4128 1734 4140
rect 1765 4131 1823 4137
rect 1765 4128 1777 4131
rect 1728 4100 1777 4128
rect 1728 4088 1734 4100
rect 1765 4097 1777 4100
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 2032 4063 2090 4069
rect 2032 4029 2044 4063
rect 2078 4060 2090 4063
rect 3326 4060 3332 4072
rect 2078 4032 3332 4060
rect 2078 4029 2090 4032
rect 2032 4023 2090 4029
rect 3326 4020 3332 4032
rect 3384 4060 3390 4072
rect 3804 4060 3832 4236
rect 4356 4196 4384 4236
rect 4264 4168 4384 4196
rect 5644 4196 5672 4236
rect 6825 4233 6837 4267
rect 6871 4264 6883 4267
rect 6914 4264 6920 4276
rect 6871 4236 6920 4264
rect 6871 4233 6883 4236
rect 6825 4227 6883 4233
rect 6914 4224 6920 4236
rect 6972 4224 6978 4276
rect 14642 4264 14648 4276
rect 7024 4236 14648 4264
rect 7024 4196 7052 4236
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 8202 4196 8208 4208
rect 5644 4168 7052 4196
rect 7484 4168 8208 4196
rect 4062 4128 4068 4140
rect 4023 4100 4068 4128
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4264 4137 4292 4168
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4097 4307 4131
rect 4249 4091 4307 4097
rect 4338 4088 4344 4140
rect 4396 4128 4402 4140
rect 7484 4137 7512 4168
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 10778 4196 10784 4208
rect 8496 4168 10784 4196
rect 7469 4131 7527 4137
rect 4396 4100 4660 4128
rect 4396 4088 4402 4100
rect 4632 4069 4660 4100
rect 7469 4097 7481 4131
rect 7515 4097 7527 4131
rect 8294 4128 8300 4140
rect 7469 4091 7527 4097
rect 7760 4100 8300 4128
rect 4617 4063 4675 4069
rect 3384 4032 3832 4060
rect 3896 4032 4568 4060
rect 3384 4020 3390 4032
rect 198 3952 204 4004
rect 256 3992 262 4004
rect 3896 3992 3924 4032
rect 256 3964 3924 3992
rect 3973 3995 4031 4001
rect 256 3952 262 3964
rect 3973 3961 3985 3995
rect 4019 3992 4031 3995
rect 4430 3992 4436 4004
rect 4019 3964 4436 3992
rect 4019 3961 4031 3964
rect 3973 3955 4031 3961
rect 4430 3952 4436 3964
rect 4488 3952 4494 4004
rect 4540 3992 4568 4032
rect 4617 4029 4629 4063
rect 4663 4060 4675 4063
rect 4706 4060 4712 4072
rect 4663 4032 4712 4060
rect 4663 4029 4675 4032
rect 4617 4023 4675 4029
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 7282 4060 7288 4072
rect 4816 4032 7288 4060
rect 4816 3992 4844 4032
rect 7282 4020 7288 4032
rect 7340 4020 7346 4072
rect 4540 3964 4844 3992
rect 4884 3995 4942 4001
rect 4884 3961 4896 3995
rect 4930 3992 4942 3995
rect 5442 3992 5448 4004
rect 4930 3964 5448 3992
rect 4930 3961 4942 3964
rect 4884 3955 4942 3961
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 6454 3952 6460 4004
rect 6512 3992 6518 4004
rect 7760 3992 7788 4100
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 8386 4088 8392 4140
rect 8444 4128 8450 4140
rect 8496 4137 8524 4168
rect 8481 4131 8539 4137
rect 8481 4128 8493 4131
rect 8444 4100 8493 4128
rect 8444 4088 8450 4100
rect 8481 4097 8493 4100
rect 8527 4097 8539 4131
rect 8481 4091 8539 4097
rect 8938 4088 8944 4140
rect 8996 4128 9002 4140
rect 10060 4137 10088 4168
rect 10778 4156 10784 4168
rect 10836 4156 10842 4208
rect 11054 4156 11060 4208
rect 11112 4196 11118 4208
rect 12342 4196 12348 4208
rect 11112 4168 12348 4196
rect 11112 4156 11118 4168
rect 12342 4156 12348 4168
rect 12400 4156 12406 4208
rect 12434 4156 12440 4208
rect 12492 4196 12498 4208
rect 12492 4168 12537 4196
rect 12492 4156 12498 4168
rect 12710 4156 12716 4208
rect 12768 4196 12774 4208
rect 12768 4168 13032 4196
rect 12768 4156 12774 4168
rect 10045 4131 10103 4137
rect 8996 4100 9904 4128
rect 8996 4088 9002 4100
rect 8205 4063 8263 4069
rect 8205 4029 8217 4063
rect 8251 4060 8263 4063
rect 8570 4060 8576 4072
rect 8251 4032 8576 4060
rect 8251 4029 8263 4032
rect 8205 4023 8263 4029
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 9766 4060 9772 4072
rect 9727 4032 9772 4060
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 9876 4060 9904 4100
rect 10045 4097 10057 4131
rect 10091 4097 10103 4131
rect 10962 4128 10968 4140
rect 10923 4100 10968 4128
rect 10045 4091 10103 4097
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 12894 4128 12900 4140
rect 11348 4100 12900 4128
rect 10781 4063 10839 4069
rect 10781 4060 10793 4063
rect 9876 4032 10793 4060
rect 10781 4029 10793 4032
rect 10827 4029 10839 4063
rect 10781 4023 10839 4029
rect 10873 4063 10931 4069
rect 10873 4029 10885 4063
rect 10919 4060 10931 4063
rect 11348 4060 11376 4100
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 13004 4137 13032 4168
rect 13354 4156 13360 4208
rect 13412 4196 13418 4208
rect 15930 4196 15936 4208
rect 13412 4168 15936 4196
rect 13412 4156 13418 4168
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 13906 4088 13912 4140
rect 13964 4128 13970 4140
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13964 4100 14013 4128
rect 13964 4088 13970 4100
rect 14001 4097 14013 4100
rect 14047 4128 14059 4131
rect 14047 4100 14596 4128
rect 14047 4097 14059 4100
rect 14001 4091 14059 4097
rect 10919 4032 11376 4060
rect 11609 4063 11667 4069
rect 10919 4029 10931 4032
rect 10873 4023 10931 4029
rect 11609 4029 11621 4063
rect 11655 4029 11667 4063
rect 11609 4023 11667 4029
rect 11885 4063 11943 4069
rect 11885 4029 11897 4063
rect 11931 4060 11943 4063
rect 13170 4060 13176 4072
rect 11931 4032 13176 4060
rect 11931 4029 11943 4032
rect 11885 4023 11943 4029
rect 10226 3992 10232 4004
rect 6512 3964 7788 3992
rect 7852 3964 10232 3992
rect 6512 3952 6518 3964
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 3145 3927 3203 3933
rect 3145 3924 3157 3927
rect 2832 3896 3157 3924
rect 2832 3884 2838 3896
rect 3145 3893 3157 3896
rect 3191 3893 3203 3927
rect 3602 3924 3608 3936
rect 3563 3896 3608 3924
rect 3145 3887 3203 3893
rect 3602 3884 3608 3896
rect 3660 3884 3666 3936
rect 5994 3924 6000 3936
rect 5955 3896 6000 3924
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 6270 3924 6276 3936
rect 6231 3896 6276 3924
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 7852 3933 7880 3964
rect 10226 3952 10232 3964
rect 10284 3952 10290 4004
rect 7193 3927 7251 3933
rect 7193 3924 7205 3927
rect 7156 3896 7205 3924
rect 7156 3884 7162 3896
rect 7193 3893 7205 3896
rect 7239 3893 7251 3927
rect 7193 3887 7251 3893
rect 7837 3927 7895 3933
rect 7837 3893 7849 3927
rect 7883 3893 7895 3927
rect 7837 3887 7895 3893
rect 8202 3884 8208 3936
rect 8260 3924 8266 3936
rect 8297 3927 8355 3933
rect 8297 3924 8309 3927
rect 8260 3896 8309 3924
rect 8260 3884 8266 3896
rect 8297 3893 8309 3896
rect 8343 3893 8355 3927
rect 8297 3887 8355 3893
rect 9401 3927 9459 3933
rect 9401 3893 9413 3927
rect 9447 3924 9459 3927
rect 9766 3924 9772 3936
rect 9447 3896 9772 3924
rect 9447 3893 9459 3896
rect 9401 3887 9459 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 9861 3927 9919 3933
rect 9861 3893 9873 3927
rect 9907 3924 9919 3927
rect 9950 3924 9956 3936
rect 9907 3896 9956 3924
rect 9907 3893 9919 3896
rect 9861 3887 9919 3893
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 10410 3924 10416 3936
rect 10371 3896 10416 3924
rect 10410 3884 10416 3896
rect 10468 3884 10474 3936
rect 10796 3924 10824 4023
rect 10962 3952 10968 4004
rect 11020 3992 11026 4004
rect 11020 3964 11284 3992
rect 11020 3952 11026 3964
rect 11146 3924 11152 3936
rect 10796 3896 11152 3924
rect 11146 3884 11152 3896
rect 11204 3884 11210 3936
rect 11256 3924 11284 3964
rect 11330 3952 11336 4004
rect 11388 3992 11394 4004
rect 11624 3992 11652 4023
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 14568 4069 14596 4100
rect 14642 4088 14648 4140
rect 14700 4128 14706 4140
rect 15764 4137 15792 4168
rect 15930 4156 15936 4168
rect 15988 4156 15994 4208
rect 16574 4156 16580 4208
rect 16632 4196 16638 4208
rect 16945 4199 17003 4205
rect 16945 4196 16957 4199
rect 16632 4168 16957 4196
rect 16632 4156 16638 4168
rect 16945 4165 16957 4168
rect 16991 4165 17003 4199
rect 16945 4159 17003 4165
rect 14737 4131 14795 4137
rect 14737 4128 14749 4131
rect 14700 4100 14749 4128
rect 14700 4088 14706 4100
rect 14737 4097 14749 4100
rect 14783 4097 14795 4131
rect 14737 4091 14795 4097
rect 15749 4131 15807 4137
rect 15749 4097 15761 4131
rect 15795 4097 15807 4131
rect 15749 4091 15807 4097
rect 14553 4063 14611 4069
rect 14553 4029 14565 4063
rect 14599 4029 14611 4063
rect 15657 4063 15715 4069
rect 15657 4060 15669 4063
rect 14553 4023 14611 4029
rect 14752 4032 15669 4060
rect 11388 3964 11652 3992
rect 12805 3995 12863 4001
rect 11388 3952 11394 3964
rect 12805 3961 12817 3995
rect 12851 3992 12863 3995
rect 12851 3964 13032 3992
rect 12851 3961 12863 3964
rect 12805 3955 12863 3961
rect 13004 3936 13032 3964
rect 13906 3952 13912 4004
rect 13964 3992 13970 4004
rect 14642 3992 14648 4004
rect 13964 3964 14228 3992
rect 14603 3964 14648 3992
rect 13964 3952 13970 3964
rect 12342 3924 12348 3936
rect 11256 3896 12348 3924
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 12618 3884 12624 3936
rect 12676 3924 12682 3936
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 12676 3896 12909 3924
rect 12676 3884 12682 3896
rect 12897 3893 12909 3896
rect 12943 3893 12955 3927
rect 12897 3887 12955 3893
rect 12986 3884 12992 3936
rect 13044 3884 13050 3936
rect 13354 3884 13360 3936
rect 13412 3924 13418 3936
rect 13814 3924 13820 3936
rect 13412 3896 13820 3924
rect 13412 3884 13418 3896
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 14200 3933 14228 3964
rect 14642 3952 14648 3964
rect 14700 3952 14706 4004
rect 14185 3927 14243 3933
rect 14185 3893 14197 3927
rect 14231 3893 14243 3927
rect 14185 3887 14243 3893
rect 14366 3884 14372 3936
rect 14424 3924 14430 3936
rect 14752 3924 14780 4032
rect 15657 4029 15669 4032
rect 15703 4060 15715 4063
rect 15930 4060 15936 4072
rect 15703 4032 15936 4060
rect 15703 4029 15715 4032
rect 15657 4023 15715 4029
rect 15930 4020 15936 4032
rect 15988 4020 15994 4072
rect 16206 4060 16212 4072
rect 16167 4032 16212 4060
rect 16206 4020 16212 4032
rect 16264 4020 16270 4072
rect 16761 4063 16819 4069
rect 16761 4029 16773 4063
rect 16807 4029 16819 4063
rect 16761 4023 16819 4029
rect 15102 3952 15108 4004
rect 15160 3992 15166 4004
rect 16776 3992 16804 4023
rect 15160 3964 16804 3992
rect 15160 3952 15166 3964
rect 15194 3924 15200 3936
rect 14424 3896 14780 3924
rect 15155 3896 15200 3924
rect 14424 3884 14430 3896
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 15562 3924 15568 3936
rect 15523 3896 15568 3924
rect 15562 3884 15568 3896
rect 15620 3884 15626 3936
rect 15746 3884 15752 3936
rect 15804 3924 15810 3936
rect 16393 3927 16451 3933
rect 16393 3924 16405 3927
rect 15804 3896 16405 3924
rect 15804 3884 15810 3896
rect 16393 3893 16405 3896
rect 16439 3893 16451 3927
rect 16393 3887 16451 3893
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 22462 3924 22468 3936
rect 16816 3896 22468 3924
rect 16816 3884 16822 3896
rect 22462 3884 22468 3896
rect 22520 3884 22526 3936
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 1578 3680 1584 3732
rect 1636 3720 1642 3732
rect 1949 3723 2007 3729
rect 1949 3720 1961 3723
rect 1636 3692 1961 3720
rect 1636 3680 1642 3692
rect 1949 3689 1961 3692
rect 1995 3689 2007 3723
rect 1949 3683 2007 3689
rect 3329 3723 3387 3729
rect 3329 3689 3341 3723
rect 3375 3720 3387 3723
rect 6270 3720 6276 3732
rect 3375 3692 6276 3720
rect 3375 3689 3387 3692
rect 3329 3683 3387 3689
rect 6270 3680 6276 3692
rect 6328 3680 6334 3732
rect 6825 3723 6883 3729
rect 6825 3689 6837 3723
rect 6871 3720 6883 3723
rect 7742 3720 7748 3732
rect 6871 3692 7748 3720
rect 6871 3689 6883 3692
rect 6825 3683 6883 3689
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 8386 3720 8392 3732
rect 8347 3692 8392 3720
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 8570 3680 8576 3732
rect 8628 3720 8634 3732
rect 9122 3720 9128 3732
rect 8628 3692 9128 3720
rect 8628 3680 8634 3692
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9490 3680 9496 3732
rect 9548 3720 9554 3732
rect 9950 3720 9956 3732
rect 9548 3692 9956 3720
rect 9548 3680 9554 3692
rect 9950 3680 9956 3692
rect 10008 3680 10014 3732
rect 10594 3680 10600 3732
rect 10652 3720 10658 3732
rect 10962 3720 10968 3732
rect 10652 3692 10968 3720
rect 10652 3680 10658 3692
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 11241 3723 11299 3729
rect 11241 3689 11253 3723
rect 11287 3689 11299 3723
rect 11241 3683 11299 3689
rect 11333 3723 11391 3729
rect 11333 3689 11345 3723
rect 11379 3720 11391 3723
rect 12802 3720 12808 3732
rect 11379 3692 12808 3720
rect 11379 3689 11391 3692
rect 11333 3683 11391 3689
rect 2148 3624 2452 3652
rect 1118 3476 1124 3528
rect 1176 3516 1182 3528
rect 2148 3516 2176 3624
rect 2314 3584 2320 3596
rect 2275 3556 2320 3584
rect 2314 3544 2320 3556
rect 2372 3544 2378 3596
rect 2424 3584 2452 3624
rect 4154 3612 4160 3664
rect 4212 3652 4218 3664
rect 6365 3655 6423 3661
rect 6365 3652 6377 3655
rect 4212 3624 6377 3652
rect 4212 3612 4218 3624
rect 6365 3621 6377 3624
rect 6411 3652 6423 3655
rect 7098 3652 7104 3664
rect 6411 3624 7104 3652
rect 6411 3621 6423 3624
rect 6365 3615 6423 3621
rect 7098 3612 7104 3624
rect 7156 3612 7162 3664
rect 7208 3624 7871 3652
rect 3142 3584 3148 3596
rect 2424 3556 3148 3584
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 3418 3584 3424 3596
rect 3379 3556 3424 3584
rect 3418 3544 3424 3556
rect 3476 3544 3482 3596
rect 4413 3587 4471 3593
rect 4413 3584 4425 3587
rect 3988 3556 4425 3584
rect 1176 3488 2176 3516
rect 2409 3519 2467 3525
rect 1176 3476 1182 3488
rect 2409 3485 2421 3519
rect 2455 3516 2467 3519
rect 2498 3516 2504 3528
rect 2455 3488 2504 3516
rect 2455 3485 2467 3488
rect 2409 3479 2467 3485
rect 2498 3476 2504 3488
rect 2556 3476 2562 3528
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3516 2651 3519
rect 2958 3516 2964 3528
rect 2639 3488 2964 3516
rect 2639 3485 2651 3488
rect 2593 3479 2651 3485
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 3510 3516 3516 3528
rect 3471 3488 3516 3516
rect 3510 3476 3516 3488
rect 3568 3516 3574 3528
rect 3988 3516 4016 3556
rect 4413 3553 4425 3556
rect 4459 3553 4471 3587
rect 4413 3547 4471 3553
rect 5994 3544 6000 3596
rect 6052 3584 6058 3596
rect 7208 3584 7236 3624
rect 6052 3556 7236 3584
rect 7276 3587 7334 3593
rect 6052 3544 6058 3556
rect 7276 3553 7288 3587
rect 7322 3584 7334 3587
rect 7742 3584 7748 3596
rect 7322 3556 7748 3584
rect 7322 3553 7334 3556
rect 7276 3547 7334 3553
rect 7742 3544 7748 3556
rect 7800 3544 7806 3596
rect 7843 3584 7871 3624
rect 8312 3624 10364 3652
rect 8312 3584 8340 3624
rect 9030 3584 9036 3596
rect 7843 3556 8340 3584
rect 8991 3556 9036 3584
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 9674 3544 9680 3596
rect 9732 3584 9738 3596
rect 10117 3587 10175 3593
rect 10117 3584 10129 3587
rect 9732 3556 10129 3584
rect 9732 3544 9738 3556
rect 10117 3553 10129 3556
rect 10163 3553 10175 3587
rect 10336 3584 10364 3624
rect 10410 3612 10416 3664
rect 10468 3652 10474 3664
rect 11054 3652 11060 3664
rect 10468 3624 11060 3652
rect 10468 3612 10474 3624
rect 11054 3612 11060 3624
rect 11112 3612 11118 3664
rect 11146 3612 11152 3664
rect 11204 3652 11210 3664
rect 11256 3652 11284 3683
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 12897 3723 12955 3729
rect 12897 3689 12909 3723
rect 12943 3720 12955 3723
rect 13078 3720 13084 3732
rect 12943 3692 13084 3720
rect 12943 3689 12955 3692
rect 12897 3683 12955 3689
rect 13078 3680 13084 3692
rect 13136 3720 13142 3732
rect 14185 3723 14243 3729
rect 13136 3692 13860 3720
rect 13136 3680 13142 3692
rect 11204 3624 11468 3652
rect 11204 3612 11210 3624
rect 11333 3587 11391 3593
rect 11333 3584 11345 3587
rect 10336 3556 11345 3584
rect 10117 3547 10175 3553
rect 11333 3553 11345 3556
rect 11379 3553 11391 3587
rect 11440 3584 11468 3624
rect 13262 3612 13268 3664
rect 13320 3652 13326 3664
rect 13446 3652 13452 3664
rect 13320 3624 13452 3652
rect 13320 3612 13326 3624
rect 13446 3612 13452 3624
rect 13504 3652 13510 3664
rect 13541 3655 13599 3661
rect 13541 3652 13553 3655
rect 13504 3624 13553 3652
rect 13504 3612 13510 3624
rect 13541 3621 13553 3624
rect 13587 3621 13599 3655
rect 13541 3615 13599 3621
rect 13633 3655 13691 3661
rect 13633 3621 13645 3655
rect 13679 3652 13691 3655
rect 13722 3652 13728 3664
rect 13679 3624 13728 3652
rect 13679 3621 13691 3624
rect 13633 3615 13691 3621
rect 13722 3612 13728 3624
rect 13780 3612 13786 3664
rect 11773 3587 11831 3593
rect 11773 3584 11785 3587
rect 11440 3556 11785 3584
rect 11333 3547 11391 3553
rect 11773 3553 11785 3556
rect 11819 3553 11831 3587
rect 13832 3584 13860 3692
rect 14185 3689 14197 3723
rect 14231 3689 14243 3723
rect 14185 3683 14243 3689
rect 14200 3596 14228 3683
rect 14366 3680 14372 3732
rect 14424 3720 14430 3732
rect 14645 3723 14703 3729
rect 14645 3720 14657 3723
rect 14424 3692 14657 3720
rect 14424 3680 14430 3692
rect 14645 3689 14657 3692
rect 14691 3720 14703 3723
rect 16298 3720 16304 3732
rect 14691 3692 16304 3720
rect 14691 3689 14703 3692
rect 14645 3683 14703 3689
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 15930 3612 15936 3664
rect 15988 3652 15994 3664
rect 15988 3624 17172 3652
rect 15988 3612 15994 3624
rect 11773 3547 11831 3553
rect 13740 3556 13860 3584
rect 4154 3516 4160 3528
rect 3568 3488 4016 3516
rect 4115 3488 4160 3516
rect 3568 3476 3574 3488
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 6454 3516 6460 3528
rect 5920 3488 6460 3516
rect 658 3408 664 3460
rect 716 3448 722 3460
rect 716 3420 4200 3448
rect 716 3408 722 3420
rect 2961 3383 3019 3389
rect 2961 3349 2973 3383
rect 3007 3380 3019 3383
rect 4062 3380 4068 3392
rect 3007 3352 4068 3380
rect 3007 3349 3019 3352
rect 2961 3343 3019 3349
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 4172 3380 4200 3420
rect 5442 3408 5448 3460
rect 5500 3448 5506 3460
rect 5537 3451 5595 3457
rect 5537 3448 5549 3451
rect 5500 3420 5549 3448
rect 5500 3408 5506 3420
rect 5537 3417 5549 3420
rect 5583 3417 5595 3451
rect 5537 3411 5595 3417
rect 5920 3380 5948 3488
rect 6454 3476 6460 3488
rect 6512 3476 6518 3528
rect 6546 3476 6552 3528
rect 6604 3516 6610 3528
rect 6641 3519 6699 3525
rect 6641 3516 6653 3519
rect 6604 3488 6653 3516
rect 6604 3476 6610 3488
rect 6641 3485 6653 3488
rect 6687 3516 6699 3519
rect 6825 3519 6883 3525
rect 6825 3516 6837 3519
rect 6687 3488 6837 3516
rect 6687 3485 6699 3488
rect 6641 3479 6699 3485
rect 6825 3485 6837 3488
rect 6871 3485 6883 3519
rect 7006 3516 7012 3528
rect 6967 3488 7012 3516
rect 6825 3479 6883 3485
rect 7006 3476 7012 3488
rect 7064 3476 7070 3528
rect 9858 3516 9864 3528
rect 9819 3488 9864 3516
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 11514 3516 11520 3528
rect 11475 3488 11520 3516
rect 11514 3476 11520 3488
rect 11572 3476 11578 3528
rect 13354 3516 13360 3528
rect 13096 3488 13360 3516
rect 13096 3448 13124 3488
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 13740 3525 13768 3556
rect 14182 3544 14188 3596
rect 14240 3544 14246 3596
rect 14274 3544 14280 3596
rect 14332 3584 14338 3596
rect 14553 3587 14611 3593
rect 14553 3584 14565 3587
rect 14332 3556 14565 3584
rect 14332 3544 14338 3556
rect 14553 3553 14565 3556
rect 14599 3553 14611 3587
rect 14553 3547 14611 3553
rect 15194 3544 15200 3596
rect 15252 3584 15258 3596
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 15252 3556 15301 3584
rect 15252 3544 15258 3556
rect 15289 3553 15301 3556
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 15565 3587 15623 3593
rect 15565 3553 15577 3587
rect 15611 3584 15623 3587
rect 16025 3587 16083 3593
rect 16025 3584 16037 3587
rect 15611 3556 16037 3584
rect 15611 3553 15623 3556
rect 15565 3547 15623 3553
rect 16025 3553 16037 3556
rect 16071 3553 16083 3587
rect 16025 3547 16083 3553
rect 16577 3587 16635 3593
rect 16577 3553 16589 3587
rect 16623 3584 16635 3587
rect 16666 3584 16672 3596
rect 16623 3556 16672 3584
rect 16623 3553 16635 3556
rect 16577 3547 16635 3553
rect 16666 3544 16672 3556
rect 16724 3544 16730 3596
rect 17144 3593 17172 3624
rect 17129 3587 17187 3593
rect 17129 3553 17141 3587
rect 17175 3553 17187 3587
rect 17129 3547 17187 3553
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3485 13783 3519
rect 14458 3516 14464 3528
rect 13725 3479 13783 3485
rect 13832 3488 14464 3516
rect 12452 3420 13124 3448
rect 13173 3451 13231 3457
rect 12452 3392 12480 3420
rect 13173 3417 13185 3451
rect 13219 3448 13231 3451
rect 13832 3448 13860 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 14737 3519 14795 3525
rect 14737 3485 14749 3519
rect 14783 3485 14795 3519
rect 20162 3516 20168 3528
rect 14737 3479 14795 3485
rect 14835 3488 20168 3516
rect 13219 3420 13860 3448
rect 14108 3420 14320 3448
rect 13219 3417 13231 3420
rect 13173 3411 13231 3417
rect 4172 3352 5948 3380
rect 5997 3383 6055 3389
rect 5997 3349 6009 3383
rect 6043 3380 6055 3383
rect 7742 3380 7748 3392
rect 6043 3352 7748 3380
rect 6043 3349 6055 3352
rect 5997 3343 6055 3349
rect 7742 3340 7748 3352
rect 7800 3340 7806 3392
rect 9217 3383 9275 3389
rect 9217 3349 9229 3383
rect 9263 3380 9275 3383
rect 12158 3380 12164 3392
rect 9263 3352 12164 3380
rect 9263 3349 9275 3352
rect 9217 3343 9275 3349
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 12434 3340 12440 3392
rect 12492 3340 12498 3392
rect 12618 3340 12624 3392
rect 12676 3380 12682 3392
rect 14108 3380 14136 3420
rect 12676 3352 14136 3380
rect 14292 3380 14320 3420
rect 14550 3408 14556 3460
rect 14608 3448 14614 3460
rect 14752 3448 14780 3479
rect 14608 3420 14780 3448
rect 14608 3408 14614 3420
rect 14835 3380 14863 3488
rect 20162 3476 20168 3488
rect 20220 3476 20226 3528
rect 16761 3451 16819 3457
rect 16761 3417 16773 3451
rect 16807 3448 16819 3451
rect 17402 3448 17408 3460
rect 16807 3420 17408 3448
rect 16807 3417 16819 3420
rect 16761 3411 16819 3417
rect 17402 3408 17408 3420
rect 17460 3408 17466 3460
rect 14292 3352 14863 3380
rect 16209 3383 16267 3389
rect 12676 3340 12682 3352
rect 16209 3349 16221 3383
rect 16255 3380 16267 3383
rect 16942 3380 16948 3392
rect 16255 3352 16948 3380
rect 16255 3349 16267 3352
rect 16209 3343 16267 3349
rect 16942 3340 16948 3352
rect 17000 3340 17006 3392
rect 17310 3380 17316 3392
rect 17271 3352 17316 3380
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 4709 3179 4767 3185
rect 2332 3148 4016 3176
rect 2332 2981 2360 3148
rect 3988 3108 4016 3148
rect 4709 3145 4721 3179
rect 4755 3176 4767 3179
rect 9674 3176 9680 3188
rect 4755 3148 9536 3176
rect 9635 3148 9680 3176
rect 4755 3145 4767 3148
rect 4709 3139 4767 3145
rect 5258 3108 5264 3120
rect 3988 3080 5264 3108
rect 5258 3068 5264 3080
rect 5316 3068 5322 3120
rect 7006 3068 7012 3120
rect 7064 3108 7070 3120
rect 8113 3111 8171 3117
rect 8113 3108 8125 3111
rect 7064 3080 8125 3108
rect 7064 3068 7070 3080
rect 8113 3077 8125 3080
rect 8159 3077 8171 3111
rect 8113 3071 8171 3077
rect 2406 3000 2412 3052
rect 2464 3040 2470 3052
rect 2593 3043 2651 3049
rect 2464 3012 2509 3040
rect 2464 3000 2470 3012
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 2639 3012 2912 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 2317 2975 2375 2981
rect 2317 2941 2329 2975
rect 2363 2941 2375 2975
rect 2317 2935 2375 2941
rect 2682 2904 2688 2916
rect 1964 2876 2688 2904
rect 1964 2845 1992 2876
rect 2682 2864 2688 2876
rect 2740 2864 2746 2916
rect 1949 2839 2007 2845
rect 1949 2805 1961 2839
rect 1995 2805 2007 2839
rect 2884 2836 2912 3012
rect 2958 3000 2964 3052
rect 3016 3040 3022 3052
rect 5353 3043 5411 3049
rect 3016 3012 3061 3040
rect 3016 3000 3022 3012
rect 5353 3009 5365 3043
rect 5399 3040 5411 3043
rect 5442 3040 5448 3052
rect 5399 3012 5448 3040
rect 5399 3009 5411 3012
rect 5353 3003 5411 3009
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3040 6423 3043
rect 6546 3040 6552 3052
rect 6411 3012 6552 3040
rect 6411 3009 6423 3012
rect 6365 3003 6423 3009
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 7742 3040 7748 3052
rect 7703 3012 7748 3040
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3040 7987 3043
rect 9508 3040 9536 3148
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 10137 3179 10195 3185
rect 10137 3145 10149 3179
rect 10183 3176 10195 3179
rect 12618 3176 12624 3188
rect 10183 3148 12624 3176
rect 10183 3145 10195 3148
rect 10137 3139 10195 3145
rect 12618 3136 12624 3148
rect 12676 3136 12682 3188
rect 12802 3136 12808 3188
rect 12860 3176 12866 3188
rect 15657 3179 15715 3185
rect 12860 3148 15056 3176
rect 12860 3136 12866 3148
rect 9858 3068 9864 3120
rect 9916 3108 9922 3120
rect 10042 3108 10048 3120
rect 9916 3080 10048 3108
rect 9916 3068 9922 3080
rect 10042 3068 10048 3080
rect 10100 3068 10106 3120
rect 10505 3111 10563 3117
rect 10505 3077 10517 3111
rect 10551 3108 10563 3111
rect 11790 3108 11796 3120
rect 10551 3080 11796 3108
rect 10551 3077 10563 3080
rect 10505 3071 10563 3077
rect 11790 3068 11796 3080
rect 11848 3068 11854 3120
rect 12437 3111 12495 3117
rect 12437 3077 12449 3111
rect 12483 3077 12495 3111
rect 12437 3071 12495 3077
rect 14461 3111 14519 3117
rect 14461 3077 14473 3111
rect 14507 3077 14519 3111
rect 14461 3071 14519 3077
rect 10318 3040 10324 3052
rect 7975 3012 8432 3040
rect 9508 3012 10324 3040
rect 7975 3009 7987 3012
rect 7929 3003 7987 3009
rect 8404 2984 8432 3012
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 10594 3000 10600 3052
rect 10652 3040 10658 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10652 3012 10977 3040
rect 10652 3000 10658 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 11204 3012 11249 3040
rect 11204 3000 11210 3012
rect 11330 3000 11336 3052
rect 11388 3040 11394 3052
rect 12452 3040 12480 3071
rect 11388 3012 12480 3040
rect 11388 3000 11394 3012
rect 12526 3000 12532 3052
rect 12584 3040 12590 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12584 3012 13001 3040
rect 12584 3000 12590 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 14093 3043 14151 3049
rect 14093 3009 14105 3043
rect 14139 3040 14151 3043
rect 14366 3040 14372 3052
rect 14139 3012 14372 3040
rect 14139 3009 14151 3012
rect 14093 3003 14151 3009
rect 14366 3000 14372 3012
rect 14424 3000 14430 3052
rect 14476 3040 14504 3071
rect 14642 3040 14648 3052
rect 14476 3012 14648 3040
rect 14642 3000 14648 3012
rect 14700 3000 14706 3052
rect 15028 3049 15056 3148
rect 15657 3145 15669 3179
rect 15703 3176 15715 3179
rect 22002 3176 22008 3188
rect 15703 3148 22008 3176
rect 15703 3145 15715 3148
rect 15657 3139 15715 3145
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 16577 3111 16635 3117
rect 16577 3077 16589 3111
rect 16623 3108 16635 3111
rect 19702 3108 19708 3120
rect 16623 3080 19708 3108
rect 16623 3077 16635 3080
rect 16577 3071 16635 3077
rect 19702 3068 19708 3080
rect 19760 3068 19766 3120
rect 15013 3043 15071 3049
rect 15013 3009 15025 3043
rect 15059 3009 15071 3043
rect 15013 3003 15071 3009
rect 15562 3000 15568 3052
rect 15620 3040 15626 3052
rect 15620 3012 18460 3040
rect 15620 3000 15626 3012
rect 3050 2932 3056 2984
rect 3108 2972 3114 2984
rect 3217 2975 3275 2981
rect 3217 2972 3229 2975
rect 3108 2944 3229 2972
rect 3108 2932 3114 2944
rect 3217 2941 3229 2944
rect 3263 2941 3275 2975
rect 3217 2935 3275 2941
rect 4062 2932 4068 2984
rect 4120 2972 4126 2984
rect 5077 2975 5135 2981
rect 5077 2972 5089 2975
rect 4120 2944 5089 2972
rect 4120 2932 4126 2944
rect 5077 2941 5089 2944
rect 5123 2941 5135 2975
rect 5077 2935 5135 2941
rect 5994 2932 6000 2984
rect 6052 2972 6058 2984
rect 6181 2975 6239 2981
rect 6181 2972 6193 2975
rect 6052 2944 6193 2972
rect 6052 2932 6058 2944
rect 6181 2941 6193 2944
rect 6227 2972 6239 2975
rect 8113 2975 8171 2981
rect 6227 2944 8064 2972
rect 6227 2941 6239 2944
rect 6181 2935 6239 2941
rect 3418 2864 3424 2916
rect 3476 2904 3482 2916
rect 5350 2904 5356 2916
rect 3476 2876 5356 2904
rect 3476 2864 3482 2876
rect 5350 2864 5356 2876
rect 5408 2864 5414 2916
rect 7653 2907 7711 2913
rect 7653 2904 7665 2907
rect 5736 2876 7665 2904
rect 3510 2836 3516 2848
rect 2884 2808 3516 2836
rect 1949 2799 2007 2805
rect 3510 2796 3516 2808
rect 3568 2836 3574 2848
rect 4341 2839 4399 2845
rect 4341 2836 4353 2839
rect 3568 2808 4353 2836
rect 3568 2796 3574 2808
rect 4341 2805 4353 2808
rect 4387 2836 4399 2839
rect 4614 2836 4620 2848
rect 4387 2808 4620 2836
rect 4387 2805 4399 2808
rect 4341 2799 4399 2805
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 5736 2845 5764 2876
rect 7653 2873 7665 2876
rect 7699 2873 7711 2907
rect 8036 2904 8064 2944
rect 8113 2941 8125 2975
rect 8159 2972 8171 2975
rect 8297 2975 8355 2981
rect 8297 2972 8309 2975
rect 8159 2944 8309 2972
rect 8159 2941 8171 2944
rect 8113 2935 8171 2941
rect 8297 2941 8309 2944
rect 8343 2941 8355 2975
rect 8297 2935 8355 2941
rect 8386 2932 8392 2984
rect 8444 2972 8450 2984
rect 8553 2975 8611 2981
rect 8553 2972 8565 2975
rect 8444 2944 8565 2972
rect 8444 2932 8450 2944
rect 8553 2941 8565 2944
rect 8599 2941 8611 2975
rect 9858 2972 9864 2984
rect 8553 2935 8611 2941
rect 8680 2944 9864 2972
rect 8680 2904 8708 2944
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 9953 2975 10011 2981
rect 9953 2941 9965 2975
rect 9999 2972 10011 2975
rect 10134 2972 10140 2984
rect 9999 2944 10140 2972
rect 9999 2941 10011 2944
rect 9953 2935 10011 2941
rect 10134 2932 10140 2944
rect 10192 2972 10198 2984
rect 10413 2975 10471 2981
rect 10413 2972 10425 2975
rect 10192 2944 10425 2972
rect 10192 2932 10198 2944
rect 10413 2941 10425 2944
rect 10459 2941 10471 2975
rect 10413 2935 10471 2941
rect 10870 2932 10876 2984
rect 10928 2972 10934 2984
rect 10928 2944 10973 2972
rect 10928 2932 10934 2944
rect 11606 2932 11612 2984
rect 11664 2972 11670 2984
rect 11664 2944 11709 2972
rect 11664 2932 11670 2944
rect 12066 2932 12072 2984
rect 12124 2972 12130 2984
rect 13817 2975 13875 2981
rect 13817 2972 13829 2975
rect 12124 2944 13829 2972
rect 12124 2932 12130 2944
rect 13817 2941 13829 2944
rect 13863 2941 13875 2975
rect 13817 2935 13875 2941
rect 13909 2975 13967 2981
rect 13909 2941 13921 2975
rect 13955 2972 13967 2975
rect 13998 2972 14004 2984
rect 13955 2944 14004 2972
rect 13955 2941 13967 2944
rect 13909 2935 13967 2941
rect 13998 2932 14004 2944
rect 14056 2932 14062 2984
rect 15470 2972 15476 2984
rect 15431 2944 15476 2972
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 16390 2972 16396 2984
rect 16351 2944 16396 2972
rect 16390 2932 16396 2944
rect 16448 2932 16454 2984
rect 18432 2981 18460 3012
rect 16945 2975 17003 2981
rect 16945 2941 16957 2975
rect 16991 2941 17003 2975
rect 16945 2935 17003 2941
rect 18417 2975 18475 2981
rect 18417 2941 18429 2975
rect 18463 2941 18475 2975
rect 18417 2935 18475 2941
rect 8036 2876 8708 2904
rect 7653 2867 7711 2873
rect 9030 2864 9036 2916
rect 9088 2904 9094 2916
rect 11885 2907 11943 2913
rect 11885 2904 11897 2907
rect 9088 2876 11897 2904
rect 9088 2864 9094 2876
rect 11885 2873 11897 2876
rect 11931 2873 11943 2907
rect 11885 2867 11943 2873
rect 12618 2864 12624 2916
rect 12676 2904 12682 2916
rect 12897 2907 12955 2913
rect 12897 2904 12909 2907
rect 12676 2876 12909 2904
rect 12676 2864 12682 2876
rect 12897 2873 12909 2876
rect 12943 2904 12955 2907
rect 12943 2876 14228 2904
rect 12943 2873 12955 2876
rect 12897 2867 12955 2873
rect 5721 2839 5779 2845
rect 5224 2808 5269 2836
rect 5224 2796 5230 2808
rect 5721 2805 5733 2839
rect 5767 2805 5779 2839
rect 6086 2836 6092 2848
rect 6047 2808 6092 2836
rect 5721 2799 5779 2805
rect 6086 2796 6092 2808
rect 6144 2796 6150 2848
rect 7285 2839 7343 2845
rect 7285 2805 7297 2839
rect 7331 2836 7343 2839
rect 8294 2836 8300 2848
rect 7331 2808 8300 2836
rect 7331 2805 7343 2808
rect 7285 2799 7343 2805
rect 8294 2796 8300 2808
rect 8352 2796 8358 2848
rect 8662 2796 8668 2848
rect 8720 2836 8726 2848
rect 10134 2836 10140 2848
rect 8720 2808 10140 2836
rect 8720 2796 8726 2808
rect 10134 2796 10140 2808
rect 10192 2796 10198 2848
rect 10413 2839 10471 2845
rect 10413 2805 10425 2839
rect 10459 2836 10471 2839
rect 12805 2839 12863 2845
rect 12805 2836 12817 2839
rect 10459 2808 12817 2836
rect 10459 2805 10471 2808
rect 10413 2799 10471 2805
rect 12805 2805 12817 2808
rect 12851 2805 12863 2839
rect 12805 2799 12863 2805
rect 13262 2796 13268 2848
rect 13320 2836 13326 2848
rect 13449 2839 13507 2845
rect 13449 2836 13461 2839
rect 13320 2808 13461 2836
rect 13320 2796 13326 2808
rect 13449 2805 13461 2808
rect 13495 2805 13507 2839
rect 14200 2836 14228 2876
rect 14366 2864 14372 2916
rect 14424 2904 14430 2916
rect 14921 2907 14979 2913
rect 14921 2904 14933 2907
rect 14424 2876 14933 2904
rect 14424 2864 14430 2876
rect 14921 2873 14933 2876
rect 14967 2873 14979 2907
rect 14921 2867 14979 2873
rect 14458 2836 14464 2848
rect 14200 2808 14464 2836
rect 13449 2799 13507 2805
rect 14458 2796 14464 2808
rect 14516 2796 14522 2848
rect 14829 2839 14887 2845
rect 14829 2805 14841 2839
rect 14875 2836 14887 2839
rect 15194 2836 15200 2848
rect 14875 2808 15200 2836
rect 14875 2805 14887 2808
rect 14829 2799 14887 2805
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 16114 2796 16120 2848
rect 16172 2836 16178 2848
rect 16960 2836 16988 2935
rect 17770 2864 17776 2916
rect 17828 2904 17834 2916
rect 21542 2904 21548 2916
rect 17828 2876 21548 2904
rect 17828 2864 17834 2876
rect 21542 2864 21548 2876
rect 21600 2864 21606 2916
rect 16172 2808 16988 2836
rect 17129 2839 17187 2845
rect 16172 2796 16178 2808
rect 17129 2805 17141 2839
rect 17175 2836 17187 2839
rect 17862 2836 17868 2848
rect 17175 2808 17868 2836
rect 17175 2805 17187 2808
rect 17129 2799 17187 2805
rect 17862 2796 17868 2808
rect 17920 2796 17926 2848
rect 18601 2839 18659 2845
rect 18601 2805 18613 2839
rect 18647 2836 18659 2839
rect 19242 2836 19248 2848
rect 18647 2808 19248 2836
rect 18647 2805 18659 2808
rect 18601 2799 18659 2805
rect 19242 2796 19248 2808
rect 19300 2796 19306 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 2314 2632 2320 2644
rect 1995 2604 2320 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 2314 2592 2320 2604
rect 2372 2592 2378 2644
rect 2682 2592 2688 2644
rect 2740 2632 2746 2644
rect 3326 2632 3332 2644
rect 2740 2604 3332 2632
rect 2740 2592 2746 2604
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 3421 2635 3479 2641
rect 3421 2601 3433 2635
rect 3467 2632 3479 2635
rect 3789 2635 3847 2641
rect 3789 2632 3801 2635
rect 3467 2604 3801 2632
rect 3467 2601 3479 2604
rect 3421 2595 3479 2601
rect 3789 2601 3801 2604
rect 3835 2601 3847 2635
rect 3789 2595 3847 2601
rect 4065 2635 4123 2641
rect 4065 2601 4077 2635
rect 4111 2632 4123 2635
rect 5166 2632 5172 2644
rect 4111 2604 5172 2632
rect 4111 2601 4123 2604
rect 4065 2595 4123 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5350 2592 5356 2644
rect 5408 2632 5414 2644
rect 5537 2635 5595 2641
rect 5537 2632 5549 2635
rect 5408 2604 5549 2632
rect 5408 2592 5414 2604
rect 5537 2601 5549 2604
rect 5583 2601 5595 2635
rect 5537 2595 5595 2601
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 8662 2632 8668 2644
rect 5868 2604 8668 2632
rect 5868 2592 5874 2604
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 10226 2632 10232 2644
rect 10187 2604 10232 2632
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 10597 2635 10655 2641
rect 10597 2601 10609 2635
rect 10643 2632 10655 2635
rect 10870 2632 10876 2644
rect 10643 2604 10876 2632
rect 10643 2601 10655 2604
rect 10597 2595 10655 2601
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11149 2635 11207 2641
rect 11149 2632 11161 2635
rect 11112 2604 11161 2632
rect 11112 2592 11118 2604
rect 11149 2601 11161 2604
rect 11195 2601 11207 2635
rect 11149 2595 11207 2601
rect 11241 2635 11299 2641
rect 11241 2601 11253 2635
rect 11287 2632 11299 2635
rect 11330 2632 11336 2644
rect 11287 2604 11336 2632
rect 11287 2601 11299 2604
rect 11241 2595 11299 2601
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 12989 2635 13047 2641
rect 12989 2601 13001 2635
rect 13035 2632 13047 2635
rect 14182 2632 14188 2644
rect 13035 2604 14188 2632
rect 13035 2601 13047 2604
rect 12989 2595 13047 2601
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 14458 2592 14464 2644
rect 14516 2632 14522 2644
rect 14829 2635 14887 2641
rect 14516 2604 14780 2632
rect 14516 2592 14522 2604
rect 3694 2524 3700 2576
rect 3752 2564 3758 2576
rect 4433 2567 4491 2573
rect 4433 2564 4445 2567
rect 3752 2536 4445 2564
rect 3752 2524 3758 2536
rect 4433 2533 4445 2536
rect 4479 2533 4491 2567
rect 4433 2527 4491 2533
rect 5074 2524 5080 2576
rect 5132 2564 5138 2576
rect 7469 2567 7527 2573
rect 7469 2564 7481 2567
rect 5132 2536 7481 2564
rect 5132 2524 5138 2536
rect 7469 2533 7481 2536
rect 7515 2533 7527 2567
rect 7469 2527 7527 2533
rect 8294 2524 8300 2576
rect 8352 2564 8358 2576
rect 9033 2567 9091 2573
rect 9033 2564 9045 2567
rect 8352 2536 9045 2564
rect 8352 2524 8358 2536
rect 9033 2533 9045 2536
rect 9079 2533 9091 2567
rect 9033 2527 9091 2533
rect 9766 2524 9772 2576
rect 9824 2564 9830 2576
rect 10137 2567 10195 2573
rect 10137 2564 10149 2567
rect 9824 2536 10149 2564
rect 9824 2524 9830 2536
rect 10137 2533 10149 2536
rect 10183 2533 10195 2567
rect 10137 2527 10195 2533
rect 11606 2524 11612 2576
rect 11664 2564 11670 2576
rect 13081 2567 13139 2573
rect 13081 2564 13093 2567
rect 11664 2536 13093 2564
rect 11664 2524 11670 2536
rect 13081 2533 13093 2536
rect 13127 2533 13139 2567
rect 13081 2527 13139 2533
rect 13446 2524 13452 2576
rect 13504 2564 13510 2576
rect 14752 2564 14780 2604
rect 14829 2601 14841 2635
rect 14875 2632 14887 2635
rect 15470 2632 15476 2644
rect 14875 2604 15476 2632
rect 14875 2601 14887 2604
rect 14829 2595 14887 2601
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 15657 2635 15715 2641
rect 15657 2601 15669 2635
rect 15703 2632 15715 2635
rect 17770 2632 17776 2644
rect 15703 2604 17776 2632
rect 15703 2601 15715 2604
rect 15657 2595 15715 2601
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 13504 2536 14688 2564
rect 14752 2536 16620 2564
rect 13504 2524 13510 2536
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2496 2375 2499
rect 2682 2496 2688 2508
rect 2363 2468 2688 2496
rect 2363 2465 2375 2468
rect 2317 2459 2375 2465
rect 2682 2456 2688 2468
rect 2740 2456 2746 2508
rect 3326 2496 3332 2508
rect 3287 2468 3332 2496
rect 3326 2456 3332 2468
rect 3384 2456 3390 2508
rect 5445 2499 5503 2505
rect 5445 2496 5457 2499
rect 3528 2468 5457 2496
rect 2406 2428 2412 2440
rect 2367 2400 2412 2428
rect 2406 2388 2412 2400
rect 2464 2388 2470 2440
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2774 2428 2780 2440
rect 2639 2400 2780 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2774 2388 2780 2400
rect 2832 2428 2838 2440
rect 3418 2428 3424 2440
rect 2832 2400 3424 2428
rect 2832 2388 2838 2400
rect 3418 2388 3424 2400
rect 3476 2388 3482 2440
rect 2961 2363 3019 2369
rect 2961 2329 2973 2363
rect 3007 2360 3019 2363
rect 3528 2360 3556 2468
rect 5445 2465 5457 2468
rect 5491 2465 5503 2499
rect 10594 2496 10600 2508
rect 5445 2459 5503 2465
rect 8680 2468 10600 2496
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2397 3663 2431
rect 3605 2391 3663 2397
rect 3007 2332 3556 2360
rect 3620 2360 3648 2391
rect 4154 2388 4160 2440
rect 4212 2428 4218 2440
rect 4525 2431 4583 2437
rect 4525 2428 4537 2431
rect 4212 2400 4537 2428
rect 4212 2388 4218 2400
rect 4525 2397 4537 2400
rect 4571 2397 4583 2431
rect 4525 2391 4583 2397
rect 4614 2388 4620 2440
rect 4672 2428 4678 2440
rect 5629 2431 5687 2437
rect 5629 2428 5641 2431
rect 4672 2400 4717 2428
rect 5460 2400 5641 2428
rect 4672 2388 4678 2400
rect 4632 2360 4660 2388
rect 5460 2372 5488 2400
rect 5629 2397 5641 2400
rect 5675 2397 5687 2431
rect 7558 2428 7564 2440
rect 7519 2400 7564 2428
rect 5629 2391 5687 2397
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 7742 2428 7748 2440
rect 7703 2400 7748 2428
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 3620 2332 4660 2360
rect 4724 2332 5212 2360
rect 3007 2329 3019 2332
rect 2961 2323 3019 2329
rect 3789 2295 3847 2301
rect 3789 2261 3801 2295
rect 3835 2292 3847 2295
rect 4724 2292 4752 2332
rect 5074 2292 5080 2304
rect 3835 2264 4752 2292
rect 5035 2264 5080 2292
rect 3835 2261 3847 2264
rect 3789 2255 3847 2261
rect 5074 2252 5080 2264
rect 5132 2252 5138 2304
rect 5184 2292 5212 2332
rect 5442 2320 5448 2372
rect 5500 2320 5506 2372
rect 7101 2363 7159 2369
rect 7101 2329 7113 2363
rect 7147 2360 7159 2363
rect 8110 2360 8116 2372
rect 7147 2332 8116 2360
rect 7147 2329 7159 2332
rect 7101 2323 7159 2329
rect 8110 2320 8116 2332
rect 8168 2320 8174 2372
rect 8680 2369 8708 2468
rect 10594 2456 10600 2468
rect 10652 2456 10658 2508
rect 10778 2456 10784 2508
rect 10836 2496 10842 2508
rect 11790 2496 11796 2508
rect 10836 2468 11376 2496
rect 11751 2468 11796 2496
rect 10836 2456 10842 2468
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9674 2428 9680 2440
rect 9355 2400 9680 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 8665 2363 8723 2369
rect 8665 2329 8677 2363
rect 8711 2329 8723 2363
rect 9140 2360 9168 2391
rect 9674 2388 9680 2400
rect 9732 2428 9738 2440
rect 11348 2437 11376 2468
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 11974 2456 11980 2508
rect 12032 2496 12038 2508
rect 12032 2468 13308 2496
rect 12032 2456 12038 2468
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 9732 2400 10333 2428
rect 9732 2388 9738 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 11333 2431 11391 2437
rect 11333 2397 11345 2431
rect 11379 2397 11391 2431
rect 11333 2391 11391 2397
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2397 12127 2431
rect 13170 2428 13176 2440
rect 13131 2400 13176 2428
rect 12069 2391 12127 2397
rect 10781 2363 10839 2369
rect 10781 2360 10793 2363
rect 9140 2332 10793 2360
rect 8665 2323 8723 2329
rect 10781 2329 10793 2332
rect 10827 2329 10839 2363
rect 12084 2360 12112 2391
rect 13170 2388 13176 2400
rect 13228 2388 13234 2440
rect 13280 2360 13308 2468
rect 13354 2456 13360 2508
rect 13412 2496 13418 2508
rect 14660 2505 14688 2536
rect 14001 2499 14059 2505
rect 14001 2496 14013 2499
rect 13412 2468 14013 2496
rect 13412 2456 13418 2468
rect 14001 2465 14013 2468
rect 14047 2465 14059 2499
rect 14001 2459 14059 2465
rect 14093 2499 14151 2505
rect 14093 2465 14105 2499
rect 14139 2496 14151 2499
rect 14645 2499 14703 2505
rect 14139 2468 14596 2496
rect 14139 2465 14151 2468
rect 14093 2459 14151 2465
rect 14182 2428 14188 2440
rect 14143 2400 14188 2428
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 14568 2428 14596 2468
rect 14645 2465 14657 2499
rect 14691 2465 14703 2499
rect 14645 2459 14703 2465
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2496 15531 2499
rect 15838 2496 15844 2508
rect 15519 2468 15844 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 15838 2456 15844 2468
rect 15896 2456 15902 2508
rect 16025 2499 16083 2505
rect 16025 2465 16037 2499
rect 16071 2496 16083 2499
rect 16114 2496 16120 2508
rect 16071 2468 16120 2496
rect 16071 2465 16083 2468
rect 16025 2459 16083 2465
rect 16114 2456 16120 2468
rect 16172 2456 16178 2508
rect 16592 2505 16620 2536
rect 16577 2499 16635 2505
rect 16577 2465 16589 2499
rect 16623 2465 16635 2499
rect 17494 2496 17500 2508
rect 17455 2468 17500 2496
rect 16577 2459 16635 2465
rect 17494 2456 17500 2468
rect 17552 2456 17558 2508
rect 16850 2428 16856 2440
rect 14568 2400 16856 2428
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 13633 2363 13691 2369
rect 13633 2360 13645 2363
rect 12084 2332 12848 2360
rect 13280 2332 13645 2360
rect 10781 2323 10839 2329
rect 5626 2292 5632 2304
rect 5184 2264 5632 2292
rect 5626 2252 5632 2264
rect 5684 2252 5690 2304
rect 9769 2295 9827 2301
rect 9769 2261 9781 2295
rect 9815 2292 9827 2295
rect 10597 2295 10655 2301
rect 10597 2292 10609 2295
rect 9815 2264 10609 2292
rect 9815 2261 9827 2264
rect 9769 2255 9827 2261
rect 10597 2261 10609 2264
rect 10643 2261 10655 2295
rect 12618 2292 12624 2304
rect 12579 2264 12624 2292
rect 10597 2255 10655 2261
rect 12618 2252 12624 2264
rect 12676 2252 12682 2304
rect 12820 2292 12848 2332
rect 13633 2329 13645 2332
rect 13679 2329 13691 2363
rect 15102 2360 15108 2372
rect 13633 2323 13691 2329
rect 14752 2332 15108 2360
rect 14752 2292 14780 2332
rect 15102 2320 15108 2332
rect 15160 2320 15166 2372
rect 16022 2320 16028 2372
rect 16080 2360 16086 2372
rect 16761 2363 16819 2369
rect 16761 2360 16773 2363
rect 16080 2332 16773 2360
rect 16080 2320 16086 2332
rect 16761 2329 16773 2332
rect 16807 2329 16819 2363
rect 16761 2323 16819 2329
rect 12820 2264 14780 2292
rect 16209 2295 16267 2301
rect 16209 2261 16221 2295
rect 16255 2292 16267 2295
rect 16482 2292 16488 2304
rect 16255 2264 16488 2292
rect 16255 2261 16267 2264
rect 16209 2255 16267 2261
rect 16482 2252 16488 2264
rect 16540 2252 16546 2304
rect 17681 2295 17739 2301
rect 17681 2261 17693 2295
rect 17727 2292 17739 2295
rect 17954 2292 17960 2304
rect 17727 2264 17960 2292
rect 17727 2261 17739 2264
rect 17681 2255 17739 2261
rect 17954 2252 17960 2264
rect 18012 2252 18018 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 2406 2048 2412 2100
rect 2464 2088 2470 2100
rect 13262 2088 13268 2100
rect 2464 2060 13268 2088
rect 2464 2048 2470 2060
rect 13262 2048 13268 2060
rect 13320 2048 13326 2100
rect 15470 2048 15476 2100
rect 15528 2088 15534 2100
rect 21082 2088 21088 2100
rect 15528 2060 21088 2088
rect 15528 2048 15534 2060
rect 21082 2048 21088 2060
rect 21140 2048 21146 2100
rect 2682 1980 2688 2032
rect 2740 2020 2746 2032
rect 2740 1992 5028 2020
rect 2740 1980 2746 1992
rect 5000 1952 5028 1992
rect 5074 1980 5080 2032
rect 5132 2020 5138 2032
rect 14366 2020 14372 2032
rect 5132 1992 14372 2020
rect 5132 1980 5138 1992
rect 14366 1980 14372 1992
rect 14424 1980 14430 2032
rect 13906 1952 13912 1964
rect 5000 1924 13912 1952
rect 13906 1912 13912 1924
rect 13964 1912 13970 1964
rect 14090 1912 14096 1964
rect 14148 1952 14154 1964
rect 16574 1952 16580 1964
rect 14148 1924 16580 1952
rect 14148 1912 14154 1924
rect 16574 1912 16580 1924
rect 16632 1912 16638 1964
rect 2498 1844 2504 1896
rect 2556 1884 2562 1896
rect 12618 1884 12624 1896
rect 2556 1856 12624 1884
rect 2556 1844 2562 1856
rect 12618 1844 12624 1856
rect 12676 1844 12682 1896
rect 2958 1776 2964 1828
rect 3016 1816 3022 1828
rect 4890 1816 4896 1828
rect 3016 1788 4896 1816
rect 3016 1776 3022 1788
rect 4890 1776 4896 1788
rect 4948 1776 4954 1828
rect 11606 1816 11612 1828
rect 5000 1788 11612 1816
rect 3510 1708 3516 1760
rect 3568 1748 3574 1760
rect 5000 1748 5028 1788
rect 11606 1776 11612 1788
rect 11664 1776 11670 1828
rect 3568 1720 5028 1748
rect 3568 1708 3574 1720
rect 5626 1708 5632 1760
rect 5684 1748 5690 1760
rect 6638 1748 6644 1760
rect 5684 1720 6644 1748
rect 5684 1708 5690 1720
rect 6638 1708 6644 1720
rect 6696 1708 6702 1760
rect 13170 1748 13176 1760
rect 6748 1720 13176 1748
rect 3418 1640 3424 1692
rect 3476 1680 3482 1692
rect 6748 1680 6776 1720
rect 13170 1708 13176 1720
rect 13228 1708 13234 1760
rect 14550 1708 14556 1760
rect 14608 1748 14614 1760
rect 17310 1748 17316 1760
rect 14608 1720 17316 1748
rect 14608 1708 14614 1720
rect 17310 1708 17316 1720
rect 17368 1708 17374 1760
rect 3476 1652 6776 1680
rect 3476 1640 3482 1652
rect 8110 1640 8116 1692
rect 8168 1680 8174 1692
rect 8754 1680 8760 1692
rect 8168 1652 8760 1680
rect 8168 1640 8174 1652
rect 8754 1640 8760 1652
rect 8812 1640 8818 1692
rect 9306 1640 9312 1692
rect 9364 1680 9370 1692
rect 13354 1680 13360 1692
rect 9364 1652 13360 1680
rect 9364 1640 9370 1652
rect 13354 1640 13360 1652
rect 13412 1640 13418 1692
rect 2498 1572 2504 1624
rect 2556 1612 2562 1624
rect 7558 1612 7564 1624
rect 2556 1584 7564 1612
rect 2556 1572 2562 1584
rect 7558 1572 7564 1584
rect 7616 1572 7622 1624
rect 12158 1572 12164 1624
rect 12216 1612 12222 1624
rect 13170 1612 13176 1624
rect 12216 1584 13176 1612
rect 12216 1572 12222 1584
rect 13170 1572 13176 1584
rect 13228 1572 13234 1624
rect 3418 1504 3424 1556
rect 3476 1544 3482 1556
rect 9306 1544 9312 1556
rect 3476 1516 9312 1544
rect 3476 1504 3482 1516
rect 9306 1504 9312 1516
rect 9364 1504 9370 1556
rect 1578 1436 1584 1488
rect 1636 1476 1642 1488
rect 5994 1476 6000 1488
rect 1636 1448 6000 1476
rect 1636 1436 1642 1448
rect 5994 1436 6000 1448
rect 6052 1436 6058 1488
rect 2038 1368 2044 1420
rect 2096 1408 2102 1420
rect 6086 1408 6092 1420
rect 2096 1380 6092 1408
rect 2096 1368 2102 1380
rect 6086 1368 6092 1380
rect 6144 1368 6150 1420
rect 11330 1368 11336 1420
rect 11388 1408 11394 1420
rect 12342 1408 12348 1420
rect 11388 1380 12348 1408
rect 11388 1368 11394 1380
rect 12342 1368 12348 1380
rect 12400 1368 12406 1420
rect 4062 1300 4068 1352
rect 4120 1340 4126 1352
rect 14274 1340 14280 1352
rect 4120 1312 14280 1340
rect 4120 1300 4126 1312
rect 14274 1300 14280 1312
rect 14332 1300 14338 1352
rect 3970 1164 3976 1216
rect 4028 1204 4034 1216
rect 13998 1204 14004 1216
rect 4028 1176 14004 1204
rect 4028 1164 4034 1176
rect 13998 1164 14004 1176
rect 14056 1164 14062 1216
<< via1 >>
rect 4068 21088 4120 21140
rect 6276 21088 6328 21140
rect 3976 20952 4028 21004
rect 8208 20952 8260 21004
rect 3516 20816 3568 20868
rect 7380 20816 7432 20868
rect 8668 20816 8720 20868
rect 9036 20816 9088 20868
rect 3332 20680 3384 20732
rect 6460 20680 6512 20732
rect 3332 20408 3384 20460
rect 4988 20408 5040 20460
rect 5724 20408 5776 20460
rect 6828 20408 6880 20460
rect 2228 20340 2280 20392
rect 6920 20340 6972 20392
rect 2872 20272 2924 20324
rect 9772 20272 9824 20324
rect 4068 20204 4120 20256
rect 8852 20204 8904 20256
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 5172 20000 5224 20052
rect 5264 20000 5316 20052
rect 8944 20000 8996 20052
rect 2872 19932 2924 19984
rect 11796 19932 11848 19984
rect 1676 19907 1728 19916
rect 1676 19873 1685 19907
rect 1685 19873 1719 19907
rect 1719 19873 1728 19907
rect 1676 19864 1728 19873
rect 2228 19907 2280 19916
rect 2228 19873 2237 19907
rect 2237 19873 2271 19907
rect 2271 19873 2280 19907
rect 2228 19864 2280 19873
rect 3608 19864 3660 19916
rect 5632 19864 5684 19916
rect 4712 19839 4764 19848
rect 1860 19703 1912 19712
rect 1860 19669 1869 19703
rect 1869 19669 1903 19703
rect 1903 19669 1912 19703
rect 1860 19660 1912 19669
rect 2964 19703 3016 19712
rect 2964 19669 2973 19703
rect 2973 19669 3007 19703
rect 3007 19669 3016 19703
rect 2964 19660 3016 19669
rect 4160 19660 4212 19712
rect 4712 19805 4721 19839
rect 4721 19805 4755 19839
rect 4755 19805 4764 19839
rect 4712 19796 4764 19805
rect 4896 19839 4948 19848
rect 4896 19805 4905 19839
rect 4905 19805 4939 19839
rect 4939 19805 4948 19839
rect 4896 19796 4948 19805
rect 6000 19839 6052 19848
rect 6000 19805 6009 19839
rect 6009 19805 6043 19839
rect 6043 19805 6052 19839
rect 6000 19796 6052 19805
rect 5172 19728 5224 19780
rect 7012 19864 7064 19916
rect 9680 19864 9732 19916
rect 10508 19907 10560 19916
rect 9220 19839 9272 19848
rect 9220 19805 9229 19839
rect 9229 19805 9263 19839
rect 9263 19805 9272 19839
rect 9220 19796 9272 19805
rect 10508 19873 10517 19907
rect 10517 19873 10551 19907
rect 10551 19873 10560 19907
rect 10508 19864 10560 19873
rect 13176 20000 13228 20052
rect 13636 20000 13688 20052
rect 17408 20000 17460 20052
rect 12164 19932 12216 19984
rect 7288 19660 7340 19712
rect 7656 19660 7708 19712
rect 8392 19660 8444 19712
rect 10048 19796 10100 19848
rect 12348 19864 12400 19916
rect 12624 19907 12676 19916
rect 12624 19873 12633 19907
rect 12633 19873 12667 19907
rect 12667 19873 12676 19907
rect 12624 19864 12676 19873
rect 13360 19864 13412 19916
rect 19340 19932 19392 19984
rect 20168 19932 20220 19984
rect 16396 19864 16448 19916
rect 19708 19796 19760 19848
rect 18696 19660 18748 19712
rect 19340 19660 19392 19712
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 4068 19456 4120 19508
rect 5724 19456 5776 19508
rect 6920 19499 6972 19508
rect 6920 19465 6929 19499
rect 6929 19465 6963 19499
rect 6963 19465 6972 19499
rect 6920 19456 6972 19465
rect 5632 19388 5684 19440
rect 6736 19388 6788 19440
rect 7748 19388 7800 19440
rect 8300 19320 8352 19372
rect 1584 19295 1636 19304
rect 1584 19261 1593 19295
rect 1593 19261 1627 19295
rect 1627 19261 1636 19295
rect 1584 19252 1636 19261
rect 3976 19252 4028 19304
rect 2412 19227 2464 19236
rect 2412 19193 2421 19227
rect 2421 19193 2455 19227
rect 2455 19193 2464 19227
rect 2412 19184 2464 19193
rect 3056 19184 3108 19236
rect 4252 19252 4304 19304
rect 5816 19295 5868 19304
rect 1768 19159 1820 19168
rect 1768 19125 1777 19159
rect 1777 19125 1811 19159
rect 1811 19125 1820 19159
rect 1768 19116 1820 19125
rect 2136 19116 2188 19168
rect 3332 19159 3384 19168
rect 3332 19125 3341 19159
rect 3341 19125 3375 19159
rect 3375 19125 3384 19159
rect 3332 19116 3384 19125
rect 4068 19116 4120 19168
rect 4160 19116 4212 19168
rect 5448 19184 5500 19236
rect 5816 19261 5825 19295
rect 5825 19261 5859 19295
rect 5859 19261 5868 19295
rect 5816 19252 5868 19261
rect 6920 19252 6972 19304
rect 7472 19252 7524 19304
rect 4896 19116 4948 19168
rect 11060 19252 11112 19304
rect 11704 19295 11756 19304
rect 11704 19261 11713 19295
rect 11713 19261 11747 19295
rect 11747 19261 11756 19295
rect 11704 19252 11756 19261
rect 12532 19252 12584 19304
rect 14188 19252 14240 19304
rect 14280 19252 14332 19304
rect 15200 19295 15252 19304
rect 15200 19261 15209 19295
rect 15209 19261 15243 19295
rect 15243 19261 15252 19295
rect 15200 19252 15252 19261
rect 15752 19295 15804 19304
rect 15752 19261 15761 19295
rect 15761 19261 15795 19295
rect 15795 19261 15804 19295
rect 15752 19252 15804 19261
rect 16304 19295 16356 19304
rect 16304 19261 16313 19295
rect 16313 19261 16347 19295
rect 16347 19261 16356 19295
rect 16304 19252 16356 19261
rect 16856 19295 16908 19304
rect 16856 19261 16865 19295
rect 16865 19261 16899 19295
rect 16899 19261 16908 19295
rect 16856 19252 16908 19261
rect 10140 19184 10192 19236
rect 10232 19184 10284 19236
rect 12716 19227 12768 19236
rect 12716 19193 12750 19227
rect 12750 19193 12768 19227
rect 12716 19184 12768 19193
rect 13636 19184 13688 19236
rect 17500 19252 17552 19304
rect 19156 19295 19208 19304
rect 17316 19184 17368 19236
rect 19156 19261 19165 19295
rect 19165 19261 19199 19295
rect 19199 19261 19208 19295
rect 19156 19252 19208 19261
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 18696 19184 18748 19236
rect 21548 19184 21600 19236
rect 6276 19116 6328 19168
rect 8484 19116 8536 19168
rect 8576 19116 8628 19168
rect 8760 19116 8812 19168
rect 9220 19116 9272 19168
rect 12072 19116 12124 19168
rect 13820 19159 13872 19168
rect 13820 19125 13829 19159
rect 13829 19125 13863 19159
rect 13863 19125 13872 19159
rect 13820 19116 13872 19125
rect 14556 19116 14608 19168
rect 15016 19116 15068 19168
rect 15568 19116 15620 19168
rect 16028 19116 16080 19168
rect 16488 19159 16540 19168
rect 16488 19125 16497 19159
rect 16497 19125 16531 19159
rect 16531 19125 16540 19159
rect 16488 19116 16540 19125
rect 16948 19116 17000 19168
rect 17868 19116 17920 19168
rect 18512 19116 18564 19168
rect 18788 19159 18840 19168
rect 18788 19125 18797 19159
rect 18797 19125 18831 19159
rect 18831 19125 18840 19159
rect 18788 19116 18840 19125
rect 19248 19116 19300 19168
rect 20628 19116 20680 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 3332 18912 3384 18964
rect 2136 18776 2188 18828
rect 2964 18776 3016 18828
rect 2504 18751 2556 18760
rect 2504 18717 2513 18751
rect 2513 18717 2547 18751
rect 2547 18717 2556 18751
rect 2504 18708 2556 18717
rect 4252 18844 4304 18896
rect 4436 18844 4488 18896
rect 5816 18844 5868 18896
rect 6000 18887 6052 18896
rect 6000 18853 6034 18887
rect 6034 18853 6052 18887
rect 6000 18844 6052 18853
rect 7012 18912 7064 18964
rect 7656 18887 7708 18896
rect 7656 18853 7668 18887
rect 7668 18853 7708 18887
rect 7656 18844 7708 18853
rect 8300 18912 8352 18964
rect 8668 18844 8720 18896
rect 8852 18912 8904 18964
rect 9680 18912 9732 18964
rect 10876 18912 10928 18964
rect 11060 18912 11112 18964
rect 12808 18912 12860 18964
rect 8760 18776 8812 18828
rect 3424 18708 3476 18760
rect 3516 18708 3568 18760
rect 4068 18751 4120 18760
rect 4068 18717 4077 18751
rect 4077 18717 4111 18751
rect 4111 18717 4120 18751
rect 4068 18708 4120 18717
rect 5356 18708 5408 18760
rect 7288 18708 7340 18760
rect 12992 18844 13044 18896
rect 14280 18844 14332 18896
rect 16856 18844 16908 18896
rect 19708 18844 19760 18896
rect 10048 18776 10100 18828
rect 10692 18776 10744 18828
rect 11980 18776 12032 18828
rect 13268 18776 13320 18828
rect 13820 18819 13872 18828
rect 13820 18785 13829 18819
rect 13829 18785 13863 18819
rect 13863 18785 13872 18819
rect 13820 18776 13872 18785
rect 15384 18776 15436 18828
rect 18788 18819 18840 18828
rect 18788 18785 18797 18819
rect 18797 18785 18831 18819
rect 18831 18785 18840 18819
rect 18788 18776 18840 18785
rect 19340 18776 19392 18828
rect 21088 18776 21140 18828
rect 9864 18708 9916 18760
rect 10140 18708 10192 18760
rect 10600 18708 10652 18760
rect 5448 18683 5500 18692
rect 5448 18649 5457 18683
rect 5457 18649 5491 18683
rect 5491 18649 5500 18683
rect 5448 18640 5500 18649
rect 7012 18640 7064 18692
rect 8484 18640 8536 18692
rect 10324 18640 10376 18692
rect 12716 18640 12768 18692
rect 6368 18572 6420 18624
rect 6460 18572 6512 18624
rect 12072 18572 12124 18624
rect 12808 18615 12860 18624
rect 12808 18581 12817 18615
rect 12817 18581 12851 18615
rect 12851 18581 12860 18615
rect 12808 18572 12860 18581
rect 12992 18572 13044 18624
rect 15108 18572 15160 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 3056 18368 3108 18420
rect 4252 18368 4304 18420
rect 6000 18368 6052 18420
rect 6368 18368 6420 18420
rect 10324 18411 10376 18420
rect 10324 18377 10333 18411
rect 10333 18377 10367 18411
rect 10367 18377 10376 18411
rect 10324 18368 10376 18377
rect 10508 18368 10560 18420
rect 5724 18300 5776 18352
rect 7196 18300 7248 18352
rect 7748 18300 7800 18352
rect 7840 18232 7892 18284
rect 8116 18275 8168 18284
rect 8116 18241 8125 18275
rect 8125 18241 8159 18275
rect 8159 18241 8168 18275
rect 8116 18232 8168 18241
rect 9496 18300 9548 18352
rect 13728 18368 13780 18420
rect 12808 18300 12860 18352
rect 11612 18232 11664 18284
rect 11796 18275 11848 18284
rect 11796 18241 11805 18275
rect 11805 18241 11839 18275
rect 11839 18241 11848 18275
rect 11796 18232 11848 18241
rect 12624 18275 12676 18284
rect 12624 18241 12633 18275
rect 12633 18241 12667 18275
rect 12667 18241 12676 18275
rect 12624 18232 12676 18241
rect 13360 18275 13412 18284
rect 13360 18241 13369 18275
rect 13369 18241 13403 18275
rect 13403 18241 13412 18275
rect 13360 18232 13412 18241
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 2688 18164 2740 18216
rect 3516 18164 3568 18216
rect 4068 18096 4120 18148
rect 5356 18164 5408 18216
rect 6644 18164 6696 18216
rect 4896 18096 4948 18148
rect 5540 18096 5592 18148
rect 7104 18096 7156 18148
rect 9220 18164 9272 18216
rect 10416 18164 10468 18216
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 2044 18028 2096 18080
rect 7472 18071 7524 18080
rect 7472 18037 7481 18071
rect 7481 18037 7515 18071
rect 7515 18037 7524 18071
rect 7472 18028 7524 18037
rect 8024 18096 8076 18148
rect 11704 18096 11756 18148
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12440 18164 12492 18173
rect 7748 18028 7800 18080
rect 8300 18028 8352 18080
rect 11152 18071 11204 18080
rect 11152 18037 11161 18071
rect 11161 18037 11195 18071
rect 11195 18037 11204 18071
rect 11152 18028 11204 18037
rect 12072 18028 12124 18080
rect 12348 18028 12400 18080
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1676 17824 1728 17876
rect 2964 17824 3016 17876
rect 3516 17824 3568 17876
rect 4712 17824 4764 17876
rect 5540 17824 5592 17876
rect 6920 17824 6972 17876
rect 11704 17824 11756 17876
rect 11980 17867 12032 17876
rect 11980 17833 11989 17867
rect 11989 17833 12023 17867
rect 12023 17833 12032 17867
rect 11980 17824 12032 17833
rect 2320 17731 2372 17740
rect 2320 17697 2329 17731
rect 2329 17697 2363 17731
rect 2363 17697 2372 17731
rect 2320 17688 2372 17697
rect 3240 17688 3292 17740
rect 5172 17731 5224 17740
rect 5172 17697 5181 17731
rect 5181 17697 5215 17731
rect 5215 17697 5224 17731
rect 5172 17688 5224 17697
rect 5816 17756 5868 17808
rect 7840 17756 7892 17808
rect 6368 17688 6420 17740
rect 7196 17688 7248 17740
rect 8208 17688 8260 17740
rect 8760 17731 8812 17740
rect 8760 17697 8769 17731
rect 8769 17697 8803 17731
rect 8803 17697 8812 17731
rect 8760 17688 8812 17697
rect 9772 17756 9824 17808
rect 11060 17756 11112 17808
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 3608 17620 3660 17672
rect 5448 17663 5500 17672
rect 5448 17629 5457 17663
rect 5457 17629 5491 17663
rect 5491 17629 5500 17663
rect 5448 17620 5500 17629
rect 6920 17620 6972 17672
rect 1676 17527 1728 17536
rect 1676 17493 1685 17527
rect 1685 17493 1719 17527
rect 1719 17493 1728 17527
rect 1676 17484 1728 17493
rect 3056 17552 3108 17604
rect 10140 17620 10192 17672
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 9772 17552 9824 17604
rect 8300 17484 8352 17536
rect 10876 17484 10928 17536
rect 11888 17620 11940 17672
rect 19340 17824 19392 17876
rect 12348 17552 12400 17604
rect 14464 17688 14516 17740
rect 22008 17552 22060 17604
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 8208 17323 8260 17332
rect 1584 17144 1636 17196
rect 1768 17144 1820 17196
rect 3240 17187 3292 17196
rect 3240 17153 3249 17187
rect 3249 17153 3283 17187
rect 3283 17153 3292 17187
rect 3240 17144 3292 17153
rect 4252 17187 4304 17196
rect 4252 17153 4261 17187
rect 4261 17153 4295 17187
rect 4295 17153 4304 17187
rect 4252 17144 4304 17153
rect 5908 17144 5960 17196
rect 2228 17119 2280 17128
rect 2228 17085 2237 17119
rect 2237 17085 2271 17119
rect 2271 17085 2280 17119
rect 2228 17076 2280 17085
rect 4068 17076 4120 17128
rect 8208 17289 8217 17323
rect 8217 17289 8251 17323
rect 8251 17289 8260 17323
rect 8208 17280 8260 17289
rect 6920 17076 6972 17128
rect 9680 17212 9732 17264
rect 14096 17280 14148 17332
rect 3516 16940 3568 16992
rect 7104 17051 7156 17060
rect 7104 17017 7138 17051
rect 7138 17017 7156 17051
rect 7104 17008 7156 17017
rect 7288 17008 7340 17060
rect 9772 17008 9824 17060
rect 12440 17212 12492 17264
rect 10140 17187 10192 17196
rect 10140 17153 10149 17187
rect 10149 17153 10183 17187
rect 10183 17153 10192 17187
rect 10140 17144 10192 17153
rect 11152 17144 11204 17196
rect 10232 17076 10284 17128
rect 14464 17144 14516 17196
rect 13176 17076 13228 17128
rect 11060 17008 11112 17060
rect 5080 16983 5132 16992
rect 5080 16949 5089 16983
rect 5089 16949 5123 16983
rect 5123 16949 5132 16983
rect 5080 16940 5132 16949
rect 5632 16940 5684 16992
rect 6092 16983 6144 16992
rect 6092 16949 6101 16983
rect 6101 16949 6135 16983
rect 6135 16949 6144 16983
rect 6092 16940 6144 16949
rect 7380 16940 7432 16992
rect 7656 16940 7708 16992
rect 11428 16940 11480 16992
rect 11612 16940 11664 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 2228 16736 2280 16788
rect 7104 16779 7156 16788
rect 2780 16668 2832 16720
rect 3056 16668 3108 16720
rect 2320 16600 2372 16652
rect 2964 16600 3016 16652
rect 2228 16575 2280 16584
rect 2228 16541 2237 16575
rect 2237 16541 2271 16575
rect 2271 16541 2280 16575
rect 2228 16532 2280 16541
rect 4160 16600 4212 16652
rect 5908 16668 5960 16720
rect 7104 16745 7113 16779
rect 7113 16745 7147 16779
rect 7147 16745 7156 16779
rect 7104 16736 7156 16745
rect 7380 16779 7432 16788
rect 7380 16745 7389 16779
rect 7389 16745 7423 16779
rect 7423 16745 7432 16779
rect 7380 16736 7432 16745
rect 8852 16779 8904 16788
rect 8852 16745 8861 16779
rect 8861 16745 8895 16779
rect 8895 16745 8904 16779
rect 8852 16736 8904 16745
rect 9956 16736 10008 16788
rect 10048 16779 10100 16788
rect 10048 16745 10057 16779
rect 10057 16745 10091 16779
rect 10091 16745 10100 16779
rect 10876 16779 10928 16788
rect 10048 16736 10100 16745
rect 10876 16745 10885 16779
rect 10885 16745 10919 16779
rect 10919 16745 10928 16779
rect 10876 16736 10928 16745
rect 11612 16736 11664 16788
rect 11888 16779 11940 16788
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 12256 16736 12308 16788
rect 7380 16600 7432 16652
rect 3976 16464 4028 16516
rect 5540 16532 5592 16584
rect 10232 16668 10284 16720
rect 8760 16643 8812 16652
rect 8760 16609 8769 16643
rect 8769 16609 8803 16643
rect 8803 16609 8812 16643
rect 8760 16600 8812 16609
rect 9036 16600 9088 16652
rect 11520 16668 11572 16720
rect 13176 16711 13228 16720
rect 13176 16677 13185 16711
rect 13185 16677 13219 16711
rect 13219 16677 13228 16711
rect 13176 16668 13228 16677
rect 11152 16600 11204 16652
rect 11796 16600 11848 16652
rect 12348 16600 12400 16652
rect 12624 16600 12676 16652
rect 7840 16575 7892 16584
rect 7840 16541 7849 16575
rect 7849 16541 7883 16575
rect 7883 16541 7892 16575
rect 7840 16532 7892 16541
rect 7104 16464 7156 16516
rect 8760 16464 8812 16516
rect 10324 16575 10376 16584
rect 10324 16541 10333 16575
rect 10333 16541 10367 16575
rect 10367 16541 10376 16575
rect 10324 16532 10376 16541
rect 11060 16532 11112 16584
rect 1676 16439 1728 16448
rect 1676 16405 1685 16439
rect 1685 16405 1719 16439
rect 1719 16405 1728 16439
rect 1676 16396 1728 16405
rect 5448 16439 5500 16448
rect 5448 16405 5457 16439
rect 5457 16405 5491 16439
rect 5491 16405 5500 16439
rect 5448 16396 5500 16405
rect 6368 16396 6420 16448
rect 9772 16464 9824 16516
rect 9680 16439 9732 16448
rect 9680 16405 9689 16439
rect 9689 16405 9723 16439
rect 9723 16405 9732 16439
rect 9680 16396 9732 16405
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 4160 16192 4212 16244
rect 5908 16192 5960 16244
rect 6092 16192 6144 16244
rect 7380 16192 7432 16244
rect 9220 16192 9272 16244
rect 1860 16031 1912 16040
rect 1860 15997 1869 16031
rect 1869 15997 1903 16031
rect 1903 15997 1912 16031
rect 1860 15988 1912 15997
rect 2688 15988 2740 16040
rect 3976 15988 4028 16040
rect 4160 15988 4212 16040
rect 5540 15988 5592 16040
rect 8392 16124 8444 16176
rect 6092 16056 6144 16108
rect 6184 15988 6236 16040
rect 7104 16056 7156 16108
rect 8760 16056 8812 16108
rect 9220 16056 9272 16108
rect 9496 16056 9548 16108
rect 9588 15988 9640 16040
rect 9772 16124 9824 16176
rect 10692 16124 10744 16176
rect 10324 16056 10376 16108
rect 11704 16056 11756 16108
rect 10232 15988 10284 16040
rect 10508 15988 10560 16040
rect 11336 15988 11388 16040
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 14004 15988 14056 16040
rect 1492 15920 1544 15972
rect 3608 15920 3660 15972
rect 5448 15920 5500 15972
rect 3332 15852 3384 15904
rect 4988 15852 5040 15904
rect 6920 15920 6972 15972
rect 10048 15920 10100 15972
rect 11704 15920 11756 15972
rect 12164 15920 12216 15972
rect 12716 15963 12768 15972
rect 12716 15929 12750 15963
rect 12750 15929 12768 15963
rect 12716 15920 12768 15929
rect 6552 15852 6604 15904
rect 6736 15852 6788 15904
rect 11980 15852 12032 15904
rect 13360 15852 13412 15904
rect 14372 15852 14424 15904
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1584 15691 1636 15700
rect 1584 15657 1593 15691
rect 1593 15657 1627 15691
rect 1627 15657 1636 15691
rect 1584 15648 1636 15657
rect 2044 15648 2096 15700
rect 2964 15691 3016 15700
rect 2964 15657 2973 15691
rect 2973 15657 3007 15691
rect 3007 15657 3016 15691
rect 2964 15648 3016 15657
rect 3332 15691 3384 15700
rect 3332 15657 3341 15691
rect 3341 15657 3375 15691
rect 3375 15657 3384 15691
rect 3332 15648 3384 15657
rect 5080 15648 5132 15700
rect 5632 15648 5684 15700
rect 6092 15648 6144 15700
rect 9404 15648 9456 15700
rect 11336 15691 11388 15700
rect 11336 15657 11345 15691
rect 11345 15657 11379 15691
rect 11379 15657 11388 15691
rect 11336 15648 11388 15657
rect 12532 15648 12584 15700
rect 14372 15691 14424 15700
rect 10692 15580 10744 15632
rect 11888 15580 11940 15632
rect 2872 15512 2924 15564
rect 4988 15512 5040 15564
rect 6092 15512 6144 15564
rect 7288 15555 7340 15564
rect 7288 15521 7297 15555
rect 7297 15521 7331 15555
rect 7331 15521 7340 15555
rect 7288 15512 7340 15521
rect 8208 15555 8260 15564
rect 8208 15521 8242 15555
rect 8242 15521 8260 15555
rect 8208 15512 8260 15521
rect 9036 15512 9088 15564
rect 2044 15444 2096 15496
rect 3424 15487 3476 15496
rect 3424 15453 3433 15487
rect 3433 15453 3467 15487
rect 3467 15453 3476 15487
rect 3424 15444 3476 15453
rect 3608 15487 3660 15496
rect 3608 15453 3617 15487
rect 3617 15453 3651 15487
rect 3651 15453 3660 15487
rect 3608 15444 3660 15453
rect 5448 15487 5500 15496
rect 4896 15376 4948 15428
rect 5172 15376 5224 15428
rect 5448 15453 5457 15487
rect 5457 15453 5491 15487
rect 5491 15453 5500 15487
rect 5448 15444 5500 15453
rect 7012 15444 7064 15496
rect 3056 15308 3108 15360
rect 3700 15308 3752 15360
rect 5080 15308 5132 15360
rect 5448 15308 5500 15360
rect 7840 15444 7892 15496
rect 9128 15308 9180 15360
rect 11060 15351 11112 15360
rect 11060 15317 11069 15351
rect 11069 15317 11103 15351
rect 11103 15317 11112 15351
rect 11060 15308 11112 15317
rect 12716 15580 12768 15632
rect 14372 15657 14381 15691
rect 14381 15657 14415 15691
rect 14415 15657 14424 15691
rect 14372 15648 14424 15657
rect 14004 15580 14056 15632
rect 12440 15512 12492 15564
rect 14280 15512 14332 15564
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 1584 15147 1636 15156
rect 1584 15113 1593 15147
rect 1593 15113 1627 15147
rect 1627 15113 1636 15147
rect 1584 15104 1636 15113
rect 2872 15104 2924 15156
rect 204 14968 256 15020
rect 1676 14968 1728 15020
rect 2596 15011 2648 15020
rect 2596 14977 2605 15011
rect 2605 14977 2639 15011
rect 2639 14977 2648 15011
rect 2596 14968 2648 14977
rect 4252 15104 4304 15156
rect 7012 15104 7064 15156
rect 7748 15104 7800 15156
rect 8208 15147 8260 15156
rect 8208 15113 8217 15147
rect 8217 15113 8251 15147
rect 8251 15113 8260 15147
rect 8208 15104 8260 15113
rect 9496 15104 9548 15156
rect 12624 15104 12676 15156
rect 5540 15036 5592 15088
rect 10508 15036 10560 15088
rect 1492 14900 1544 14952
rect 2136 14900 2188 14952
rect 2964 14943 3016 14952
rect 2964 14909 2973 14943
rect 2973 14909 3007 14943
rect 3007 14909 3016 14943
rect 2964 14900 3016 14909
rect 5356 15011 5408 15020
rect 5356 14977 5365 15011
rect 5365 14977 5399 15011
rect 5399 14977 5408 15011
rect 5356 14968 5408 14977
rect 9128 15011 9180 15020
rect 9128 14977 9137 15011
rect 9137 14977 9171 15011
rect 9171 14977 9180 15011
rect 9128 14968 9180 14977
rect 9404 14968 9456 15020
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 6920 14900 6972 14952
rect 664 14832 716 14884
rect 2964 14764 3016 14816
rect 3332 14832 3384 14884
rect 7656 14900 7708 14952
rect 9496 14900 9548 14952
rect 10140 14900 10192 14952
rect 10600 14943 10652 14952
rect 10600 14909 10609 14943
rect 10609 14909 10643 14943
rect 10643 14909 10652 14943
rect 10600 14900 10652 14909
rect 3792 14764 3844 14816
rect 4160 14764 4212 14816
rect 4344 14764 4396 14816
rect 4712 14807 4764 14816
rect 4712 14773 4721 14807
rect 4721 14773 4755 14807
rect 4755 14773 4764 14807
rect 4712 14764 4764 14773
rect 5080 14807 5132 14816
rect 5080 14773 5089 14807
rect 5089 14773 5123 14807
rect 5123 14773 5132 14807
rect 5080 14764 5132 14773
rect 8484 14832 8536 14884
rect 12072 14968 12124 15020
rect 11060 14832 11112 14884
rect 8944 14807 8996 14816
rect 8944 14773 8953 14807
rect 8953 14773 8987 14807
rect 8987 14773 8996 14807
rect 8944 14764 8996 14773
rect 9036 14807 9088 14816
rect 9036 14773 9045 14807
rect 9045 14773 9079 14807
rect 9079 14773 9088 14807
rect 9036 14764 9088 14773
rect 10600 14764 10652 14816
rect 14004 14968 14056 15020
rect 15016 14900 15068 14952
rect 13176 14832 13228 14884
rect 15292 14832 15344 14884
rect 11980 14807 12032 14816
rect 11980 14773 11989 14807
rect 11989 14773 12023 14807
rect 12023 14773 12032 14807
rect 11980 14764 12032 14773
rect 13912 14764 13964 14816
rect 14096 14807 14148 14816
rect 14096 14773 14105 14807
rect 14105 14773 14139 14807
rect 14139 14773 14148 14807
rect 14096 14764 14148 14773
rect 14556 14807 14608 14816
rect 14556 14773 14565 14807
rect 14565 14773 14599 14807
rect 14599 14773 14608 14807
rect 14556 14764 14608 14773
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 3148 14560 3200 14612
rect 1768 14492 1820 14544
rect 3976 14560 4028 14612
rect 4712 14560 4764 14612
rect 7472 14560 7524 14612
rect 7656 14560 7708 14612
rect 8944 14560 8996 14612
rect 10600 14560 10652 14612
rect 10876 14560 10928 14612
rect 14556 14560 14608 14612
rect 2504 14424 2556 14476
rect 2412 14399 2464 14408
rect 2412 14365 2421 14399
rect 2421 14365 2455 14399
rect 2455 14365 2464 14399
rect 2412 14356 2464 14365
rect 2688 14356 2740 14408
rect 5632 14492 5684 14544
rect 6092 14492 6144 14544
rect 9496 14492 9548 14544
rect 11060 14492 11112 14544
rect 3700 14424 3752 14476
rect 6552 14424 6604 14476
rect 8024 14467 8076 14476
rect 8024 14433 8033 14467
rect 8033 14433 8067 14467
rect 8067 14433 8076 14467
rect 8024 14424 8076 14433
rect 10784 14424 10836 14476
rect 12624 14492 12676 14544
rect 15752 14492 15804 14544
rect 16212 14492 16264 14544
rect 3608 14399 3660 14408
rect 3608 14365 3617 14399
rect 3617 14365 3651 14399
rect 3651 14365 3660 14399
rect 3608 14356 3660 14365
rect 4344 14356 4396 14408
rect 6920 14356 6972 14408
rect 8116 14356 8168 14408
rect 8208 14356 8260 14408
rect 9312 14356 9364 14408
rect 9588 14356 9640 14408
rect 10508 14399 10560 14408
rect 10508 14365 10517 14399
rect 10517 14365 10551 14399
rect 10551 14365 10560 14399
rect 10508 14356 10560 14365
rect 10600 14356 10652 14408
rect 11980 14399 12032 14408
rect 4160 14288 4212 14340
rect 7288 14288 7340 14340
rect 11980 14365 11989 14399
rect 11989 14365 12023 14399
rect 12023 14365 12032 14399
rect 11980 14356 12032 14365
rect 1124 14220 1176 14272
rect 3608 14220 3660 14272
rect 6000 14220 6052 14272
rect 12440 14288 12492 14340
rect 12992 14424 13044 14476
rect 13452 14424 13504 14476
rect 13912 14356 13964 14408
rect 19156 14424 19208 14476
rect 15292 14356 15344 14408
rect 14280 14331 14332 14340
rect 14280 14297 14289 14331
rect 14289 14297 14323 14331
rect 14323 14297 14332 14331
rect 14280 14288 14332 14297
rect 7656 14263 7708 14272
rect 7656 14229 7665 14263
rect 7665 14229 7699 14263
rect 7699 14229 7708 14263
rect 7656 14220 7708 14229
rect 9496 14220 9548 14272
rect 12808 14220 12860 14272
rect 12900 14220 12952 14272
rect 15200 14288 15252 14340
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 22468 14288 22520 14340
rect 15292 14263 15344 14272
rect 15292 14229 15301 14263
rect 15301 14229 15335 14263
rect 15335 14229 15344 14263
rect 15292 14220 15344 14229
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 3424 14016 3476 14068
rect 1676 13880 1728 13932
rect 2044 13923 2096 13932
rect 1124 13812 1176 13864
rect 2044 13889 2053 13923
rect 2053 13889 2087 13923
rect 2087 13889 2096 13923
rect 2044 13880 2096 13889
rect 2136 13880 2188 13932
rect 6000 14016 6052 14068
rect 8944 14016 8996 14068
rect 9036 14016 9088 14068
rect 10784 14016 10836 14068
rect 12532 14059 12584 14068
rect 12532 14025 12541 14059
rect 12541 14025 12575 14059
rect 12575 14025 12584 14059
rect 12532 14016 12584 14025
rect 14280 14016 14332 14068
rect 4252 13880 4304 13932
rect 2688 13787 2740 13796
rect 2688 13753 2711 13787
rect 2711 13753 2740 13787
rect 2688 13744 2740 13753
rect 3608 13744 3660 13796
rect 4252 13744 4304 13796
rect 6184 13812 6236 13864
rect 6920 13948 6972 14000
rect 8024 13948 8076 14000
rect 8300 13948 8352 14000
rect 7288 13855 7340 13864
rect 7288 13821 7297 13855
rect 7297 13821 7331 13855
rect 7331 13821 7340 13855
rect 7288 13812 7340 13821
rect 7656 13812 7708 13864
rect 8484 13880 8536 13932
rect 9312 13923 9364 13932
rect 9312 13889 9321 13923
rect 9321 13889 9355 13923
rect 9355 13889 9364 13923
rect 9312 13880 9364 13889
rect 15292 13948 15344 14000
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 10968 13812 11020 13864
rect 11520 13923 11572 13932
rect 11520 13889 11529 13923
rect 11529 13889 11563 13923
rect 11563 13889 11572 13923
rect 11520 13880 11572 13889
rect 12808 13880 12860 13932
rect 12900 13812 12952 13864
rect 13452 13880 13504 13932
rect 15016 13923 15068 13932
rect 15016 13889 15025 13923
rect 15025 13889 15059 13923
rect 15059 13889 15068 13923
rect 15016 13880 15068 13889
rect 15200 13923 15252 13932
rect 15200 13889 15209 13923
rect 15209 13889 15243 13923
rect 15243 13889 15252 13923
rect 15200 13880 15252 13889
rect 15844 13880 15896 13932
rect 13912 13855 13964 13864
rect 13912 13821 13921 13855
rect 13921 13821 13955 13855
rect 13955 13821 13964 13855
rect 13912 13812 13964 13821
rect 8300 13744 8352 13796
rect 2964 13676 3016 13728
rect 3700 13676 3752 13728
rect 3792 13719 3844 13728
rect 3792 13685 3801 13719
rect 3801 13685 3835 13719
rect 3835 13685 3844 13719
rect 5816 13719 5868 13728
rect 3792 13676 3844 13685
rect 5816 13685 5825 13719
rect 5825 13685 5859 13719
rect 5859 13685 5868 13719
rect 5816 13676 5868 13685
rect 6000 13676 6052 13728
rect 6552 13676 6604 13728
rect 10140 13744 10192 13796
rect 8760 13676 8812 13728
rect 9128 13719 9180 13728
rect 9128 13685 9137 13719
rect 9137 13685 9171 13719
rect 9171 13685 9180 13719
rect 9128 13676 9180 13685
rect 9220 13719 9272 13728
rect 9220 13685 9229 13719
rect 9229 13685 9263 13719
rect 9263 13685 9272 13719
rect 9220 13676 9272 13685
rect 9680 13676 9732 13728
rect 10876 13676 10928 13728
rect 11244 13719 11296 13728
rect 11244 13685 11253 13719
rect 11253 13685 11287 13719
rect 11287 13685 11296 13719
rect 11244 13676 11296 13685
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 12900 13676 12952 13685
rect 13728 13676 13780 13728
rect 14372 13676 14424 13728
rect 14648 13744 14700 13796
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 4712 13472 4764 13524
rect 9220 13472 9272 13524
rect 2228 13404 2280 13456
rect 3424 13447 3476 13456
rect 3424 13413 3433 13447
rect 3433 13413 3467 13447
rect 3467 13413 3476 13447
rect 3424 13404 3476 13413
rect 4160 13404 4212 13456
rect 5632 13447 5684 13456
rect 5632 13413 5641 13447
rect 5641 13413 5675 13447
rect 5675 13413 5684 13447
rect 5632 13404 5684 13413
rect 5816 13404 5868 13456
rect 1584 13336 1636 13388
rect 3056 13336 3108 13388
rect 5540 13379 5592 13388
rect 2504 13268 2556 13320
rect 3424 13268 3476 13320
rect 3608 13311 3660 13320
rect 3608 13277 3617 13311
rect 3617 13277 3651 13311
rect 3651 13277 3660 13311
rect 3608 13268 3660 13277
rect 3792 13268 3844 13320
rect 5540 13345 5549 13379
rect 5549 13345 5583 13379
rect 5583 13345 5592 13379
rect 5540 13336 5592 13345
rect 8484 13336 8536 13388
rect 8760 13336 8812 13388
rect 9588 13404 9640 13456
rect 13176 13472 13228 13524
rect 13452 13515 13504 13524
rect 13452 13481 13461 13515
rect 13461 13481 13495 13515
rect 13495 13481 13504 13515
rect 13452 13472 13504 13481
rect 14096 13472 14148 13524
rect 14372 13472 14424 13524
rect 15660 13472 15712 13524
rect 10140 13404 10192 13456
rect 11060 13336 11112 13388
rect 4068 13243 4120 13252
rect 4068 13209 4077 13243
rect 4077 13209 4111 13243
rect 4111 13209 4120 13243
rect 4068 13200 4120 13209
rect 5264 13200 5316 13252
rect 6000 13268 6052 13320
rect 7380 13268 7432 13320
rect 7748 13268 7800 13320
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 10876 13268 10928 13320
rect 12164 13336 12216 13388
rect 15292 13336 15344 13388
rect 19432 13379 19484 13388
rect 19432 13345 19466 13379
rect 19466 13345 19484 13379
rect 19432 13336 19484 13345
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 14372 13311 14424 13320
rect 14372 13277 14381 13311
rect 14381 13277 14415 13311
rect 14415 13277 14424 13311
rect 14372 13268 14424 13277
rect 19156 13311 19208 13320
rect 19156 13277 19165 13311
rect 19165 13277 19199 13311
rect 19199 13277 19208 13311
rect 19156 13268 19208 13277
rect 3516 13132 3568 13184
rect 3976 13132 4028 13184
rect 5080 13132 5132 13184
rect 6092 13132 6144 13184
rect 7104 13132 7156 13184
rect 7656 13132 7708 13184
rect 8208 13132 8260 13184
rect 8300 13132 8352 13184
rect 11244 13200 11296 13252
rect 12072 13200 12124 13252
rect 14096 13200 14148 13252
rect 14464 13200 14516 13252
rect 11612 13132 11664 13184
rect 14280 13132 14332 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 2412 12971 2464 12980
rect 2412 12937 2421 12971
rect 2421 12937 2455 12971
rect 2455 12937 2464 12971
rect 2412 12928 2464 12937
rect 3700 12928 3752 12980
rect 3976 12928 4028 12980
rect 10876 12928 10928 12980
rect 12164 12928 12216 12980
rect 12624 12928 12676 12980
rect 12992 12928 13044 12980
rect 2688 12860 2740 12912
rect 3516 12860 3568 12912
rect 8760 12903 8812 12912
rect 2964 12835 3016 12844
rect 2964 12801 2973 12835
rect 2973 12801 3007 12835
rect 3007 12801 3016 12835
rect 2964 12792 3016 12801
rect 3240 12792 3292 12844
rect 2688 12724 2740 12776
rect 4068 12792 4120 12844
rect 5172 12792 5224 12844
rect 5816 12792 5868 12844
rect 6184 12835 6236 12844
rect 6184 12801 6193 12835
rect 6193 12801 6227 12835
rect 6227 12801 6236 12835
rect 6184 12792 6236 12801
rect 6092 12767 6144 12776
rect 3240 12656 3292 12708
rect 3884 12656 3936 12708
rect 2044 12631 2096 12640
rect 2044 12597 2053 12631
rect 2053 12597 2087 12631
rect 2087 12597 2096 12631
rect 2044 12588 2096 12597
rect 3424 12588 3476 12640
rect 4804 12656 4856 12708
rect 5080 12656 5132 12708
rect 4712 12588 4764 12640
rect 5632 12631 5684 12640
rect 5632 12597 5641 12631
rect 5641 12597 5675 12631
rect 5675 12597 5684 12631
rect 5632 12588 5684 12597
rect 6092 12733 6101 12767
rect 6101 12733 6135 12767
rect 6135 12733 6144 12767
rect 6092 12724 6144 12733
rect 8760 12869 8769 12903
rect 8769 12869 8803 12903
rect 8803 12869 8812 12903
rect 8760 12860 8812 12869
rect 9128 12860 9180 12912
rect 7380 12835 7432 12844
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 10416 12860 10468 12912
rect 9588 12835 9640 12844
rect 9588 12801 9597 12835
rect 9597 12801 9631 12835
rect 9631 12801 9640 12835
rect 9588 12792 9640 12801
rect 13544 12928 13596 12980
rect 19156 12928 19208 12980
rect 17316 12835 17368 12844
rect 17316 12801 17325 12835
rect 17325 12801 17359 12835
rect 17359 12801 17368 12835
rect 17316 12792 17368 12801
rect 7656 12767 7708 12776
rect 7656 12733 7690 12767
rect 7690 12733 7708 12767
rect 7656 12724 7708 12733
rect 8944 12724 8996 12776
rect 10416 12724 10468 12776
rect 10784 12724 10836 12776
rect 12992 12724 13044 12776
rect 14372 12724 14424 12776
rect 17040 12767 17092 12776
rect 17040 12733 17049 12767
rect 17049 12733 17083 12767
rect 17083 12733 17092 12767
rect 17040 12724 17092 12733
rect 11888 12656 11940 12708
rect 8392 12588 8444 12640
rect 9404 12631 9456 12640
rect 9404 12597 9413 12631
rect 9413 12597 9447 12631
rect 9447 12597 9456 12631
rect 9404 12588 9456 12597
rect 9588 12588 9640 12640
rect 12532 12588 12584 12640
rect 14188 12656 14240 12708
rect 13912 12588 13964 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 1860 12384 1912 12436
rect 2504 12427 2556 12436
rect 2504 12393 2513 12427
rect 2513 12393 2547 12427
rect 2547 12393 2556 12427
rect 2504 12384 2556 12393
rect 2688 12384 2740 12436
rect 5632 12384 5684 12436
rect 7564 12427 7616 12436
rect 7564 12393 7573 12427
rect 7573 12393 7607 12427
rect 7607 12393 7616 12427
rect 7564 12384 7616 12393
rect 7656 12427 7708 12436
rect 7656 12393 7665 12427
rect 7665 12393 7699 12427
rect 7699 12393 7708 12427
rect 7656 12384 7708 12393
rect 9404 12384 9456 12436
rect 2964 12316 3016 12368
rect 4252 12316 4304 12368
rect 1860 12291 1912 12300
rect 1860 12257 1869 12291
rect 1869 12257 1903 12291
rect 1903 12257 1912 12291
rect 1860 12248 1912 12257
rect 6000 12316 6052 12368
rect 6644 12316 6696 12368
rect 7380 12316 7432 12368
rect 8392 12316 8444 12368
rect 11060 12384 11112 12436
rect 12532 12384 12584 12436
rect 12624 12384 12676 12436
rect 12992 12384 13044 12436
rect 15292 12427 15344 12436
rect 15292 12393 15301 12427
rect 15301 12393 15335 12427
rect 15335 12393 15344 12427
rect 15292 12384 15344 12393
rect 15476 12384 15528 12436
rect 16304 12384 16356 12436
rect 11796 12316 11848 12368
rect 12440 12359 12492 12368
rect 12440 12325 12449 12359
rect 12449 12325 12483 12359
rect 12483 12325 12492 12359
rect 12440 12316 12492 12325
rect 13268 12316 13320 12368
rect 13912 12316 13964 12368
rect 14004 12316 14056 12368
rect 5264 12248 5316 12300
rect 5632 12248 5684 12300
rect 8944 12291 8996 12300
rect 8944 12257 8953 12291
rect 8953 12257 8987 12291
rect 8987 12257 8996 12291
rect 8944 12248 8996 12257
rect 11704 12248 11756 12300
rect 11888 12248 11940 12300
rect 13544 12291 13596 12300
rect 1952 12223 2004 12232
rect 1952 12189 1961 12223
rect 1961 12189 1995 12223
rect 1995 12189 2004 12223
rect 1952 12180 2004 12189
rect 3056 12180 3108 12232
rect 3608 12180 3660 12232
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 7472 12180 7524 12232
rect 8576 12180 8628 12232
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 10600 12223 10652 12232
rect 9864 12112 9916 12164
rect 9956 12112 10008 12164
rect 10600 12189 10609 12223
rect 10609 12189 10643 12223
rect 10643 12189 10652 12223
rect 10600 12180 10652 12189
rect 12164 12180 12216 12232
rect 13544 12257 13553 12291
rect 13553 12257 13587 12291
rect 13587 12257 13596 12291
rect 13544 12248 13596 12257
rect 12992 12180 13044 12232
rect 14924 12180 14976 12232
rect 15844 12223 15896 12232
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 15844 12180 15896 12189
rect 13544 12112 13596 12164
rect 5724 12044 5776 12096
rect 6184 12044 6236 12096
rect 7748 12044 7800 12096
rect 12900 12044 12952 12096
rect 13176 12044 13228 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 2780 11840 2832 11892
rect 3976 11840 4028 11892
rect 6644 11840 6696 11892
rect 8760 11840 8812 11892
rect 8944 11883 8996 11892
rect 8944 11849 8953 11883
rect 8953 11849 8987 11883
rect 8987 11849 8996 11883
rect 8944 11840 8996 11849
rect 9220 11840 9272 11892
rect 2412 11704 2464 11756
rect 3608 11747 3660 11756
rect 3608 11713 3617 11747
rect 3617 11713 3651 11747
rect 3651 11713 3660 11747
rect 3608 11704 3660 11713
rect 6000 11704 6052 11756
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 3700 11636 3752 11688
rect 3792 11636 3844 11688
rect 4804 11679 4856 11688
rect 3056 11568 3108 11620
rect 3884 11568 3936 11620
rect 4252 11611 4304 11620
rect 4252 11577 4261 11611
rect 4261 11577 4295 11611
rect 4295 11577 4304 11611
rect 4252 11568 4304 11577
rect 4804 11645 4813 11679
rect 4813 11645 4847 11679
rect 4847 11645 4856 11679
rect 4804 11636 4856 11645
rect 5540 11636 5592 11688
rect 6184 11636 6236 11688
rect 6644 11704 6696 11756
rect 10600 11772 10652 11824
rect 11888 11840 11940 11892
rect 14372 11883 14424 11892
rect 14372 11849 14381 11883
rect 14381 11849 14415 11883
rect 14415 11849 14424 11883
rect 14372 11840 14424 11849
rect 12900 11772 12952 11824
rect 7932 11704 7984 11756
rect 8668 11679 8720 11688
rect 8668 11645 8677 11679
rect 8677 11645 8711 11679
rect 8711 11645 8720 11679
rect 8668 11636 8720 11645
rect 9312 11704 9364 11756
rect 12992 11747 13044 11756
rect 9680 11636 9732 11688
rect 10416 11636 10468 11688
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 12164 11636 12216 11688
rect 13728 11636 13780 11688
rect 14188 11636 14240 11688
rect 14924 11636 14976 11688
rect 6920 11568 6972 11620
rect 7196 11568 7248 11620
rect 7288 11568 7340 11620
rect 1492 11500 1544 11552
rect 3332 11543 3384 11552
rect 3332 11509 3341 11543
rect 3341 11509 3375 11543
rect 3375 11509 3384 11543
rect 3332 11500 3384 11509
rect 7472 11500 7524 11552
rect 11060 11568 11112 11620
rect 11520 11568 11572 11620
rect 12532 11568 12584 11620
rect 13360 11568 13412 11620
rect 14096 11568 14148 11620
rect 15844 11568 15896 11620
rect 9220 11500 9272 11552
rect 10600 11500 10652 11552
rect 14372 11500 14424 11552
rect 14556 11500 14608 11552
rect 15016 11543 15068 11552
rect 15016 11509 15025 11543
rect 15025 11509 15059 11543
rect 15059 11509 15068 11543
rect 15016 11500 15068 11509
rect 15108 11543 15160 11552
rect 15108 11509 15117 11543
rect 15117 11509 15151 11543
rect 15151 11509 15160 11543
rect 15108 11500 15160 11509
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 3332 11296 3384 11348
rect 7656 11296 7708 11348
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 8668 11296 8720 11348
rect 1400 11228 1452 11280
rect 4620 11228 4672 11280
rect 5264 11228 5316 11280
rect 5908 11228 5960 11280
rect 11428 11228 11480 11280
rect 11704 11296 11756 11348
rect 12256 11296 12308 11348
rect 13820 11339 13872 11348
rect 13820 11305 13829 11339
rect 13829 11305 13863 11339
rect 13863 11305 13872 11339
rect 13820 11296 13872 11305
rect 14280 11339 14332 11348
rect 14280 11305 14289 11339
rect 14289 11305 14323 11339
rect 14323 11305 14332 11339
rect 14280 11296 14332 11305
rect 12716 11228 12768 11280
rect 12808 11228 12860 11280
rect 12900 11228 12952 11280
rect 14556 11228 14608 11280
rect 1584 11203 1636 11212
rect 1584 11169 1593 11203
rect 1593 11169 1627 11203
rect 1627 11169 1636 11203
rect 1584 11160 1636 11169
rect 4896 11160 4948 11212
rect 6460 11203 6512 11212
rect 6460 11169 6469 11203
rect 6469 11169 6503 11203
rect 6503 11169 6512 11203
rect 6460 11160 6512 11169
rect 6920 11160 6972 11212
rect 7288 11203 7340 11212
rect 7288 11169 7297 11203
rect 7297 11169 7331 11203
rect 7331 11169 7340 11203
rect 7288 11160 7340 11169
rect 8576 11160 8628 11212
rect 8944 11203 8996 11212
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 9036 11203 9088 11212
rect 9036 11169 9045 11203
rect 9045 11169 9079 11203
rect 9079 11169 9088 11203
rect 9036 11160 9088 11169
rect 9496 11160 9548 11212
rect 10324 11203 10376 11212
rect 10324 11169 10333 11203
rect 10333 11169 10367 11203
rect 10367 11169 10376 11203
rect 10324 11160 10376 11169
rect 1676 11092 1728 11144
rect 4068 11092 4120 11144
rect 4712 11024 4764 11076
rect 7196 11092 7248 11144
rect 7380 11092 7432 11144
rect 8116 11092 8168 11144
rect 9312 11092 9364 11144
rect 9588 11092 9640 11144
rect 11336 11092 11388 11144
rect 12256 11092 12308 11144
rect 14004 11160 14056 11212
rect 5724 11024 5776 11076
rect 3700 10999 3752 11008
rect 3700 10965 3709 10999
rect 3709 10965 3743 10999
rect 3743 10965 3752 10999
rect 3700 10956 3752 10965
rect 4068 10999 4120 11008
rect 4068 10965 4077 10999
rect 4077 10965 4111 10999
rect 4111 10965 4120 10999
rect 4068 10956 4120 10965
rect 5908 10956 5960 11008
rect 6644 10956 6696 11008
rect 7656 11024 7708 11076
rect 11152 11024 11204 11076
rect 7380 10999 7432 11008
rect 7380 10965 7389 10999
rect 7389 10965 7423 10999
rect 7423 10965 7432 10999
rect 7380 10956 7432 10965
rect 11888 11024 11940 11076
rect 12900 11092 12952 11144
rect 13176 11092 13228 11144
rect 13268 11092 13320 11144
rect 13820 11092 13872 11144
rect 13912 11092 13964 11144
rect 14648 11135 14700 11144
rect 14648 11101 14657 11135
rect 14657 11101 14691 11135
rect 14691 11101 14700 11135
rect 14648 11092 14700 11101
rect 13360 11024 13412 11076
rect 14556 11024 14608 11076
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 2412 10752 2464 10804
rect 3056 10795 3108 10804
rect 3056 10761 3065 10795
rect 3065 10761 3099 10795
rect 3099 10761 3108 10795
rect 3056 10752 3108 10761
rect 5632 10752 5684 10804
rect 4988 10684 5040 10736
rect 3700 10616 3752 10668
rect 4712 10659 4764 10668
rect 4712 10625 4721 10659
rect 4721 10625 4755 10659
rect 4755 10625 4764 10659
rect 4712 10616 4764 10625
rect 5080 10616 5132 10668
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 6460 10616 6512 10668
rect 11060 10795 11112 10804
rect 11060 10761 11069 10795
rect 11069 10761 11103 10795
rect 11103 10761 11112 10795
rect 11060 10752 11112 10761
rect 12808 10752 12860 10804
rect 15016 10752 15068 10804
rect 4068 10548 4120 10600
rect 4344 10548 4396 10600
rect 6552 10548 6604 10600
rect 7380 10548 7432 10600
rect 7656 10548 7708 10600
rect 8116 10591 8168 10600
rect 8116 10557 8150 10591
rect 8150 10557 8168 10591
rect 8116 10548 8168 10557
rect 8576 10548 8628 10600
rect 9680 10591 9732 10600
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 9680 10548 9732 10557
rect 11060 10548 11112 10600
rect 17500 10684 17552 10736
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 13820 10616 13872 10668
rect 12716 10548 12768 10600
rect 14648 10548 14700 10600
rect 1676 10412 1728 10464
rect 11704 10480 11756 10532
rect 4436 10455 4488 10464
rect 4436 10421 4445 10455
rect 4445 10421 4479 10455
rect 4479 10421 4488 10455
rect 4436 10412 4488 10421
rect 5908 10412 5960 10464
rect 7288 10455 7340 10464
rect 7288 10421 7297 10455
rect 7297 10421 7331 10455
rect 7331 10421 7340 10455
rect 7288 10412 7340 10421
rect 8484 10412 8536 10464
rect 9588 10412 9640 10464
rect 12624 10455 12676 10464
rect 12624 10421 12633 10455
rect 12633 10421 12667 10455
rect 12667 10421 12676 10455
rect 12624 10412 12676 10421
rect 13636 10455 13688 10464
rect 13636 10421 13645 10455
rect 13645 10421 13679 10455
rect 13679 10421 13688 10455
rect 13636 10412 13688 10421
rect 13912 10412 13964 10464
rect 14188 10455 14240 10464
rect 14188 10421 14197 10455
rect 14197 10421 14231 10455
rect 14231 10421 14240 10455
rect 14188 10412 14240 10421
rect 14280 10412 14332 10464
rect 16396 10412 16448 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 2872 10208 2924 10260
rect 4436 10208 4488 10260
rect 4988 10208 5040 10260
rect 8208 10208 8260 10260
rect 4252 10140 4304 10192
rect 5172 10140 5224 10192
rect 5816 10140 5868 10192
rect 10968 10208 11020 10260
rect 11152 10208 11204 10260
rect 11888 10208 11940 10260
rect 14372 10251 14424 10260
rect 14372 10217 14381 10251
rect 14381 10217 14415 10251
rect 14415 10217 14424 10251
rect 14372 10208 14424 10217
rect 2412 10072 2464 10124
rect 4988 10115 5040 10124
rect 4988 10081 4997 10115
rect 4997 10081 5031 10115
rect 5031 10081 5040 10115
rect 4988 10072 5040 10081
rect 12440 10140 12492 10192
rect 1676 10004 1728 10056
rect 4068 10004 4120 10056
rect 5356 10004 5408 10056
rect 4804 9936 4856 9988
rect 8484 10072 8536 10124
rect 11888 10072 11940 10124
rect 9680 10047 9732 10056
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 3240 9868 3292 9920
rect 5080 9868 5132 9920
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 7656 9868 7708 9920
rect 9680 9868 9732 9920
rect 11980 9868 12032 9920
rect 13544 10072 13596 10124
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 4712 9664 4764 9716
rect 5816 9664 5868 9716
rect 7288 9664 7340 9716
rect 8300 9664 8352 9716
rect 2780 9596 2832 9648
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 1676 9460 1728 9512
rect 4804 9596 4856 9648
rect 6644 9596 6696 9648
rect 6828 9639 6880 9648
rect 6828 9605 6837 9639
rect 6837 9605 6871 9639
rect 6871 9605 6880 9639
rect 6828 9596 6880 9605
rect 7104 9596 7156 9648
rect 9772 9596 9824 9648
rect 2504 9392 2556 9444
rect 3240 9392 3292 9444
rect 5724 9460 5776 9512
rect 6460 9392 6512 9444
rect 1860 9324 1912 9376
rect 5356 9324 5408 9376
rect 6736 9528 6788 9580
rect 8208 9528 8260 9580
rect 8760 9528 8812 9580
rect 9956 9528 10008 9580
rect 11152 9664 11204 9716
rect 11888 9596 11940 9648
rect 10048 9460 10100 9512
rect 11520 9528 11572 9580
rect 11980 9571 12032 9580
rect 11980 9537 11989 9571
rect 11989 9537 12023 9571
rect 12023 9537 12032 9571
rect 11980 9528 12032 9537
rect 12532 9528 12584 9580
rect 12164 9460 12216 9512
rect 13728 9528 13780 9580
rect 14096 9528 14148 9580
rect 14556 9528 14608 9580
rect 15016 9571 15068 9580
rect 15016 9537 15025 9571
rect 15025 9537 15059 9571
rect 15059 9537 15068 9571
rect 15016 9528 15068 9537
rect 15108 9460 15160 9512
rect 7564 9392 7616 9444
rect 8852 9392 8904 9444
rect 8944 9392 8996 9444
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 8300 9367 8352 9376
rect 7288 9324 7340 9333
rect 8300 9333 8309 9367
rect 8309 9333 8343 9367
rect 8343 9333 8352 9367
rect 8300 9324 8352 9333
rect 9864 9324 9916 9376
rect 9956 9324 10008 9376
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10508 9367 10560 9376
rect 10140 9324 10192 9333
rect 10508 9333 10517 9367
rect 10517 9333 10551 9367
rect 10551 9333 10560 9367
rect 10508 9324 10560 9333
rect 11336 9367 11388 9376
rect 11336 9333 11345 9367
rect 11345 9333 11379 9367
rect 11379 9333 11388 9367
rect 11336 9324 11388 9333
rect 14188 9392 14240 9444
rect 14648 9392 14700 9444
rect 12716 9324 12768 9376
rect 13728 9324 13780 9376
rect 14004 9324 14056 9376
rect 14464 9367 14516 9376
rect 14464 9333 14473 9367
rect 14473 9333 14507 9367
rect 14507 9333 14516 9367
rect 14464 9324 14516 9333
rect 14556 9324 14608 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 1860 9163 1912 9172
rect 1860 9129 1869 9163
rect 1869 9129 1903 9163
rect 1903 9129 1912 9163
rect 1860 9120 1912 9129
rect 2504 9120 2556 9172
rect 7380 9120 7432 9172
rect 8300 9120 8352 9172
rect 10876 9120 10928 9172
rect 10968 9163 11020 9172
rect 10968 9129 10977 9163
rect 10977 9129 11011 9163
rect 11011 9129 11020 9163
rect 12164 9163 12216 9172
rect 10968 9120 11020 9129
rect 12164 9129 12173 9163
rect 12173 9129 12207 9163
rect 12207 9129 12216 9163
rect 12164 9120 12216 9129
rect 12716 9163 12768 9172
rect 12716 9129 12725 9163
rect 12725 9129 12759 9163
rect 12759 9129 12768 9163
rect 12716 9120 12768 9129
rect 12992 9120 13044 9172
rect 14280 9120 14332 9172
rect 2136 9052 2188 9104
rect 4252 9052 4304 9104
rect 4988 9052 5040 9104
rect 3884 8984 3936 9036
rect 4160 8984 4212 9036
rect 1952 8916 2004 8968
rect 2872 8916 2924 8968
rect 3148 8916 3200 8968
rect 3332 8959 3384 8968
rect 3332 8925 3341 8959
rect 3341 8925 3375 8959
rect 3375 8925 3384 8959
rect 3332 8916 3384 8925
rect 2412 8848 2464 8900
rect 3608 8916 3660 8968
rect 6368 8984 6420 9036
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 4804 8916 4856 8968
rect 5172 8916 5224 8968
rect 6736 8916 6788 8968
rect 7472 8916 7524 8968
rect 7656 8984 7708 9036
rect 7840 8984 7892 9036
rect 8760 8984 8812 9036
rect 13360 9052 13412 9104
rect 8392 8916 8444 8968
rect 8484 8959 8536 8968
rect 8484 8925 8493 8959
rect 8493 8925 8527 8959
rect 8527 8925 8536 8959
rect 10600 8984 10652 9036
rect 10784 8984 10836 9036
rect 12072 9027 12124 9036
rect 8484 8916 8536 8925
rect 10416 8916 10468 8968
rect 11152 8959 11204 8968
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 12072 8993 12081 9027
rect 12081 8993 12115 9027
rect 12115 8993 12124 9027
rect 12072 8984 12124 8993
rect 14372 8984 14424 9036
rect 11152 8916 11204 8925
rect 12440 8916 12492 8968
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 14188 8959 14240 8968
rect 14188 8925 14197 8959
rect 14197 8925 14231 8959
rect 14231 8925 14240 8959
rect 14188 8916 14240 8925
rect 4068 8848 4120 8900
rect 10140 8848 10192 8900
rect 10508 8848 10560 8900
rect 12900 8848 12952 8900
rect 12992 8848 13044 8900
rect 15016 8916 15068 8968
rect 3976 8780 4028 8832
rect 6644 8780 6696 8832
rect 7656 8780 7708 8832
rect 7840 8823 7892 8832
rect 7840 8789 7849 8823
rect 7849 8789 7883 8823
rect 7883 8789 7892 8823
rect 7840 8780 7892 8789
rect 9680 8780 9732 8832
rect 9772 8780 9824 8832
rect 10784 8780 10836 8832
rect 12624 8780 12676 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2412 8576 2464 8628
rect 3884 8619 3936 8628
rect 3884 8585 3893 8619
rect 3893 8585 3927 8619
rect 3927 8585 3936 8619
rect 3884 8576 3936 8585
rect 1492 8415 1544 8424
rect 1492 8381 1501 8415
rect 1501 8381 1535 8415
rect 1535 8381 1544 8415
rect 1492 8372 1544 8381
rect 1676 8372 1728 8424
rect 2872 8372 2924 8424
rect 4712 8440 4764 8492
rect 5448 8576 5500 8628
rect 6460 8619 6512 8628
rect 6460 8585 6469 8619
rect 6469 8585 6503 8619
rect 6503 8585 6512 8619
rect 10048 8619 10100 8628
rect 6460 8576 6512 8585
rect 10048 8585 10057 8619
rect 10057 8585 10091 8619
rect 10091 8585 10100 8619
rect 10048 8576 10100 8585
rect 12992 8576 13044 8628
rect 10416 8551 10468 8560
rect 10416 8517 10425 8551
rect 10425 8517 10459 8551
rect 10459 8517 10468 8551
rect 10416 8508 10468 8517
rect 13820 8576 13872 8628
rect 14188 8576 14240 8628
rect 16488 8508 16540 8560
rect 12716 8440 12768 8492
rect 12900 8483 12952 8492
rect 12900 8449 12909 8483
rect 12909 8449 12943 8483
rect 12943 8449 12952 8483
rect 12900 8440 12952 8449
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 13176 8440 13228 8492
rect 15016 8483 15068 8492
rect 5632 8372 5684 8424
rect 9680 8372 9732 8424
rect 3516 8304 3568 8356
rect 7104 8304 7156 8356
rect 7472 8304 7524 8356
rect 4068 8236 4120 8288
rect 5356 8236 5408 8288
rect 5632 8236 5684 8288
rect 6276 8236 6328 8288
rect 6552 8236 6604 8288
rect 8300 8236 8352 8288
rect 12532 8372 12584 8424
rect 12624 8372 12676 8424
rect 15016 8449 15025 8483
rect 15025 8449 15059 8483
rect 15059 8449 15068 8483
rect 15016 8440 15068 8449
rect 11152 8304 11204 8356
rect 11612 8304 11664 8356
rect 12440 8304 12492 8356
rect 12900 8304 12952 8356
rect 8576 8236 8628 8288
rect 14096 8236 14148 8288
rect 15016 8304 15068 8356
rect 15200 8236 15252 8288
rect 16672 8236 16724 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 3332 8032 3384 8084
rect 4160 8032 4212 8084
rect 6644 8075 6696 8084
rect 6644 8041 6653 8075
rect 6653 8041 6687 8075
rect 6687 8041 6696 8075
rect 6644 8032 6696 8041
rect 7288 8032 7340 8084
rect 10784 8032 10836 8084
rect 11888 8032 11940 8084
rect 12624 8032 12676 8084
rect 14004 8032 14056 8084
rect 2412 7964 2464 8016
rect 7564 7964 7616 8016
rect 7656 7964 7708 8016
rect 10048 7964 10100 8016
rect 12716 7964 12768 8016
rect 12992 7964 13044 8016
rect 3884 7896 3936 7948
rect 6276 7896 6328 7948
rect 6828 7896 6880 7948
rect 7748 7896 7800 7948
rect 12164 7896 12216 7948
rect 13544 7964 13596 8016
rect 13360 7939 13412 7948
rect 13360 7905 13394 7939
rect 13394 7905 13412 7939
rect 13360 7896 13412 7905
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 5908 7828 5960 7880
rect 8300 7871 8352 7880
rect 8300 7837 8309 7871
rect 8309 7837 8343 7871
rect 8343 7837 8352 7871
rect 8300 7828 8352 7837
rect 8392 7828 8444 7880
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 1676 7692 1728 7744
rect 2872 7692 2924 7744
rect 10600 7692 10652 7744
rect 10876 7692 10928 7744
rect 13360 7692 13412 7744
rect 14556 7692 14608 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 3792 7488 3844 7540
rect 5448 7488 5500 7540
rect 5816 7488 5868 7540
rect 6828 7531 6880 7540
rect 6828 7497 6837 7531
rect 6837 7497 6871 7531
rect 6871 7497 6880 7531
rect 6828 7488 6880 7497
rect 10784 7531 10836 7540
rect 10784 7497 10793 7531
rect 10793 7497 10827 7531
rect 10827 7497 10836 7531
rect 10784 7488 10836 7497
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 1676 7284 1728 7336
rect 2872 7284 2924 7336
rect 6000 7352 6052 7404
rect 8484 7420 8536 7472
rect 6736 7352 6788 7404
rect 7472 7352 7524 7404
rect 10968 7352 11020 7404
rect 13268 7488 13320 7540
rect 11520 7420 11572 7472
rect 12072 7352 12124 7404
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 13360 7352 13412 7404
rect 15016 7395 15068 7404
rect 15016 7361 15025 7395
rect 15025 7361 15059 7395
rect 15059 7361 15068 7395
rect 15016 7352 15068 7361
rect 5448 7284 5500 7336
rect 5724 7284 5776 7336
rect 6920 7284 6972 7336
rect 2780 7216 2832 7268
rect 5908 7216 5960 7268
rect 3332 7148 3384 7200
rect 4068 7148 4120 7200
rect 8576 7216 8628 7268
rect 9220 7284 9272 7336
rect 11152 7284 11204 7336
rect 13820 7327 13872 7336
rect 13820 7293 13829 7327
rect 13829 7293 13863 7327
rect 13863 7293 13872 7327
rect 13820 7284 13872 7293
rect 16304 7284 16356 7336
rect 10048 7216 10100 7268
rect 12256 7216 12308 7268
rect 6460 7148 6512 7200
rect 9036 7148 9088 7200
rect 10508 7148 10560 7200
rect 11244 7191 11296 7200
rect 11244 7157 11253 7191
rect 11253 7157 11287 7191
rect 11287 7157 11296 7191
rect 14004 7216 14056 7268
rect 15936 7259 15988 7268
rect 15936 7225 15945 7259
rect 15945 7225 15979 7259
rect 15979 7225 15988 7259
rect 15936 7216 15988 7225
rect 11244 7148 11296 7157
rect 12532 7148 12584 7200
rect 14188 7148 14240 7200
rect 14464 7191 14516 7200
rect 14464 7157 14473 7191
rect 14473 7157 14507 7191
rect 14507 7157 14516 7191
rect 14464 7148 14516 7157
rect 15200 7148 15252 7200
rect 16580 7148 16632 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 3240 6944 3292 6996
rect 5080 6944 5132 6996
rect 8208 6944 8260 6996
rect 8392 6987 8444 6996
rect 8392 6953 8401 6987
rect 8401 6953 8435 6987
rect 8435 6953 8444 6987
rect 8392 6944 8444 6953
rect 10048 6944 10100 6996
rect 11520 6944 11572 6996
rect 11980 6944 12032 6996
rect 12532 6944 12584 6996
rect 13452 6944 13504 6996
rect 15844 6944 15896 6996
rect 5816 6876 5868 6928
rect 9220 6876 9272 6928
rect 10876 6876 10928 6928
rect 3148 6808 3200 6860
rect 6460 6808 6512 6860
rect 8484 6851 8536 6860
rect 8484 6817 8493 6851
rect 8493 6817 8527 6851
rect 8527 6817 8536 6851
rect 8484 6808 8536 6817
rect 2964 6740 3016 6792
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 5448 6740 5500 6792
rect 3792 6672 3844 6724
rect 3700 6604 3752 6656
rect 4068 6647 4120 6656
rect 4068 6613 4077 6647
rect 4077 6613 4111 6647
rect 4111 6613 4120 6647
rect 4068 6604 4120 6613
rect 7196 6672 7248 6724
rect 8300 6740 8352 6792
rect 9772 6808 9824 6860
rect 12624 6876 12676 6928
rect 9680 6783 9732 6792
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 9680 6740 9732 6749
rect 10784 6740 10836 6792
rect 12072 6783 12124 6792
rect 12072 6749 12081 6783
rect 12081 6749 12115 6783
rect 12115 6749 12124 6783
rect 13820 6851 13872 6860
rect 13820 6817 13829 6851
rect 13829 6817 13863 6851
rect 13863 6817 13872 6851
rect 13820 6808 13872 6817
rect 13912 6851 13964 6860
rect 13912 6817 13921 6851
rect 13921 6817 13955 6851
rect 13955 6817 13964 6851
rect 13912 6808 13964 6817
rect 12072 6740 12124 6749
rect 12992 6740 13044 6792
rect 13360 6740 13412 6792
rect 14004 6783 14056 6792
rect 14004 6749 14013 6783
rect 14013 6749 14047 6783
rect 14047 6749 14056 6783
rect 14004 6740 14056 6749
rect 11060 6672 11112 6724
rect 11244 6672 11296 6724
rect 12256 6672 12308 6724
rect 9956 6604 10008 6656
rect 11796 6604 11848 6656
rect 13176 6604 13228 6656
rect 15292 6647 15344 6656
rect 15292 6613 15301 6647
rect 15301 6613 15335 6647
rect 15335 6613 15344 6647
rect 15292 6604 15344 6613
rect 15568 6604 15620 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 3148 6443 3200 6452
rect 3148 6409 3157 6443
rect 3157 6409 3191 6443
rect 3191 6409 3200 6443
rect 3148 6400 3200 6409
rect 3976 6400 4028 6452
rect 10784 6400 10836 6452
rect 11152 6400 11204 6452
rect 11612 6400 11664 6452
rect 13360 6400 13412 6452
rect 10416 6332 10468 6384
rect 11152 6264 11204 6316
rect 11612 6264 11664 6316
rect 1676 6196 1728 6248
rect 3700 6196 3752 6248
rect 4252 6196 4304 6248
rect 6736 6196 6788 6248
rect 7104 6196 7156 6248
rect 4712 6128 4764 6180
rect 9036 6196 9088 6248
rect 10048 6196 10100 6248
rect 13820 6264 13872 6316
rect 16764 6307 16816 6316
rect 16764 6273 16773 6307
rect 16773 6273 16807 6307
rect 16807 6273 16816 6307
rect 16764 6264 16816 6273
rect 3424 6103 3476 6112
rect 3424 6069 3433 6103
rect 3433 6069 3467 6103
rect 3467 6069 3476 6103
rect 3424 6060 3476 6069
rect 3608 6060 3660 6112
rect 5816 6060 5868 6112
rect 8944 6103 8996 6112
rect 8944 6069 8953 6103
rect 8953 6069 8987 6103
rect 8987 6069 8996 6103
rect 8944 6060 8996 6069
rect 9772 6060 9824 6112
rect 10416 6060 10468 6112
rect 11428 6128 11480 6180
rect 14464 6196 14516 6248
rect 16488 6196 16540 6248
rect 12716 6171 12768 6180
rect 12716 6137 12750 6171
rect 12750 6137 12768 6171
rect 12716 6128 12768 6137
rect 15568 6128 15620 6180
rect 16580 6171 16632 6180
rect 10784 6060 10836 6112
rect 11336 6060 11388 6112
rect 12164 6060 12216 6112
rect 12440 6060 12492 6112
rect 12624 6060 12676 6112
rect 15936 6103 15988 6112
rect 15936 6069 15945 6103
rect 15945 6069 15979 6103
rect 15979 6069 15988 6103
rect 15936 6060 15988 6069
rect 16580 6137 16589 6171
rect 16589 6137 16623 6171
rect 16623 6137 16632 6171
rect 16580 6128 16632 6137
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 3424 5856 3476 5908
rect 4068 5788 4120 5840
rect 1860 5720 1912 5772
rect 4712 5788 4764 5840
rect 9680 5788 9732 5840
rect 10048 5831 10100 5840
rect 10048 5797 10057 5831
rect 10057 5797 10091 5831
rect 10091 5797 10100 5831
rect 10048 5788 10100 5797
rect 10508 5788 10560 5840
rect 10876 5788 10928 5840
rect 3148 5652 3200 5704
rect 5356 5720 5408 5772
rect 4712 5695 4764 5704
rect 3056 5584 3108 5636
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 5448 5695 5500 5704
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 2320 5559 2372 5568
rect 2320 5525 2329 5559
rect 2329 5525 2363 5559
rect 2363 5525 2372 5559
rect 2320 5516 2372 5525
rect 4068 5559 4120 5568
rect 4068 5525 4077 5559
rect 4077 5525 4111 5559
rect 4111 5525 4120 5559
rect 4068 5516 4120 5525
rect 6736 5584 6788 5636
rect 6920 5516 6972 5568
rect 8944 5720 8996 5772
rect 9036 5720 9088 5772
rect 10784 5720 10836 5772
rect 11244 5763 11296 5772
rect 11244 5729 11253 5763
rect 11253 5729 11287 5763
rect 11287 5729 11296 5763
rect 11244 5720 11296 5729
rect 7104 5695 7156 5704
rect 7104 5661 7113 5695
rect 7113 5661 7147 5695
rect 7147 5661 7156 5695
rect 7104 5652 7156 5661
rect 10416 5652 10468 5704
rect 10876 5652 10928 5704
rect 12072 5720 12124 5772
rect 12440 5788 12492 5840
rect 13176 5720 13228 5772
rect 14464 5788 14516 5840
rect 13820 5763 13872 5772
rect 13820 5729 13854 5763
rect 13854 5729 13872 5763
rect 13820 5720 13872 5729
rect 15476 5788 15528 5840
rect 16028 5788 16080 5840
rect 15936 5720 15988 5772
rect 13360 5652 13412 5704
rect 17960 5652 18012 5704
rect 19800 5652 19852 5704
rect 16396 5584 16448 5636
rect 8208 5516 8260 5568
rect 9680 5559 9732 5568
rect 9680 5525 9689 5559
rect 9689 5525 9723 5559
rect 9723 5525 9732 5559
rect 9680 5516 9732 5525
rect 10048 5516 10100 5568
rect 11980 5516 12032 5568
rect 12532 5516 12584 5568
rect 13544 5516 13596 5568
rect 15568 5516 15620 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 1860 5355 1912 5364
rect 1860 5321 1869 5355
rect 1869 5321 1903 5355
rect 1903 5321 1912 5355
rect 1860 5312 1912 5321
rect 3240 5312 3292 5364
rect 3792 5312 3844 5364
rect 6184 5355 6236 5364
rect 6184 5321 6193 5355
rect 6193 5321 6227 5355
rect 6227 5321 6236 5355
rect 6184 5312 6236 5321
rect 6276 5312 6328 5364
rect 7380 5312 7432 5364
rect 3148 5176 3200 5228
rect 5816 5176 5868 5228
rect 2320 5108 2372 5160
rect 4068 5108 4120 5160
rect 4252 5108 4304 5160
rect 4620 5108 4672 5160
rect 5448 5108 5500 5160
rect 5540 5108 5592 5160
rect 12624 5312 12676 5364
rect 12716 5312 12768 5364
rect 13912 5312 13964 5364
rect 14556 5312 14608 5364
rect 14740 5312 14792 5364
rect 16028 5312 16080 5364
rect 8944 5219 8996 5228
rect 8944 5185 8953 5219
rect 8953 5185 8987 5219
rect 8987 5185 8996 5219
rect 8944 5176 8996 5185
rect 9588 5176 9640 5228
rect 10968 5176 11020 5228
rect 9680 5108 9732 5160
rect 12256 5244 12308 5296
rect 12440 5244 12492 5296
rect 13452 5244 13504 5296
rect 11796 5219 11848 5228
rect 11796 5185 11805 5219
rect 11805 5185 11839 5219
rect 11839 5185 11848 5219
rect 11796 5176 11848 5185
rect 11888 5176 11940 5228
rect 12440 5151 12492 5160
rect 4160 5040 4212 5092
rect 6000 5040 6052 5092
rect 6552 5040 6604 5092
rect 3240 4972 3292 5024
rect 4068 4972 4120 5024
rect 11612 5040 11664 5092
rect 12440 5117 12449 5151
rect 12449 5117 12483 5151
rect 12483 5117 12492 5151
rect 12440 5108 12492 5117
rect 12532 5108 12584 5160
rect 14740 5176 14792 5228
rect 14280 5151 14332 5160
rect 14280 5117 14289 5151
rect 14289 5117 14323 5151
rect 14323 5117 14332 5151
rect 14280 5108 14332 5117
rect 15292 5108 15344 5160
rect 15476 5219 15528 5228
rect 15476 5185 15485 5219
rect 15485 5185 15519 5219
rect 15519 5185 15528 5219
rect 15476 5176 15528 5185
rect 15752 5176 15804 5228
rect 16120 5176 16172 5228
rect 17408 5219 17460 5228
rect 17408 5185 17417 5219
rect 17417 5185 17451 5219
rect 17451 5185 17460 5219
rect 17408 5176 17460 5185
rect 19800 5151 19852 5160
rect 19800 5117 19809 5151
rect 19809 5117 19843 5151
rect 19843 5117 19852 5151
rect 19800 5108 19852 5117
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 10140 4972 10192 5024
rect 12072 4972 12124 5024
rect 12992 5040 13044 5092
rect 13452 5040 13504 5092
rect 12440 4972 12492 5024
rect 12532 4972 12584 5024
rect 14004 4972 14056 5024
rect 15016 4972 15068 5024
rect 15292 5015 15344 5024
rect 15292 4981 15301 5015
rect 15301 4981 15335 5015
rect 15335 4981 15344 5015
rect 15292 4972 15344 4981
rect 15752 4972 15804 5024
rect 16028 4972 16080 5024
rect 16856 5015 16908 5024
rect 16856 4981 16865 5015
rect 16865 4981 16899 5015
rect 16899 4981 16908 5015
rect 16856 4972 16908 4981
rect 20628 4972 20680 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 4068 4811 4120 4820
rect 4068 4777 4077 4811
rect 4077 4777 4111 4811
rect 4111 4777 4120 4811
rect 4068 4768 4120 4777
rect 4804 4768 4856 4820
rect 5264 4768 5316 4820
rect 5540 4811 5592 4820
rect 5540 4777 5549 4811
rect 5549 4777 5583 4811
rect 5583 4777 5592 4811
rect 5540 4768 5592 4777
rect 6552 4811 6604 4820
rect 6552 4777 6561 4811
rect 6561 4777 6595 4811
rect 6595 4777 6604 4811
rect 6552 4768 6604 4777
rect 7656 4768 7708 4820
rect 10140 4768 10192 4820
rect 12532 4768 12584 4820
rect 12624 4768 12676 4820
rect 13912 4811 13964 4820
rect 13912 4777 13921 4811
rect 13921 4777 13955 4811
rect 13955 4777 13964 4811
rect 13912 4768 13964 4777
rect 14372 4811 14424 4820
rect 14372 4777 14381 4811
rect 14381 4777 14415 4811
rect 14415 4777 14424 4811
rect 15292 4811 15344 4820
rect 14372 4768 14424 4777
rect 3976 4700 4028 4752
rect 1676 4632 1728 4684
rect 2780 4632 2832 4684
rect 3148 4632 3200 4684
rect 4160 4632 4212 4684
rect 4896 4700 4948 4752
rect 5356 4700 5408 4752
rect 9772 4743 9824 4752
rect 9772 4709 9781 4743
rect 9781 4709 9815 4743
rect 9815 4709 9824 4743
rect 9772 4700 9824 4709
rect 10048 4700 10100 4752
rect 15292 4777 15301 4811
rect 15301 4777 15335 4811
rect 15335 4777 15344 4811
rect 15292 4768 15344 4777
rect 15752 4811 15804 4820
rect 15752 4777 15761 4811
rect 15761 4777 15795 4811
rect 15795 4777 15804 4811
rect 15752 4768 15804 4777
rect 16304 4811 16356 4820
rect 16304 4777 16313 4811
rect 16313 4777 16347 4811
rect 16347 4777 16356 4811
rect 16304 4768 16356 4777
rect 16764 4743 16816 4752
rect 6920 4675 6972 4684
rect 6920 4641 6929 4675
rect 6929 4641 6963 4675
rect 6963 4641 6972 4675
rect 6920 4632 6972 4641
rect 8668 4632 8720 4684
rect 9312 4632 9364 4684
rect 3424 4607 3476 4616
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 4712 4607 4764 4616
rect 2964 4471 3016 4480
rect 2964 4437 2973 4471
rect 2973 4437 3007 4471
rect 3007 4437 3016 4471
rect 2964 4428 3016 4437
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 6092 4564 6144 4616
rect 6736 4564 6788 4616
rect 7564 4564 7616 4616
rect 8208 4607 8260 4616
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 8300 4564 8352 4616
rect 9220 4607 9272 4616
rect 8484 4496 8536 4548
rect 8392 4428 8444 4480
rect 8576 4471 8628 4480
rect 8576 4437 8585 4471
rect 8585 4437 8619 4471
rect 8619 4437 8628 4471
rect 8576 4428 8628 4437
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 9956 4564 10008 4616
rect 10048 4564 10100 4616
rect 10968 4632 11020 4684
rect 10876 4607 10928 4616
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 11888 4607 11940 4616
rect 10876 4564 10928 4573
rect 11888 4573 11897 4607
rect 11897 4573 11931 4607
rect 11931 4573 11940 4607
rect 11888 4564 11940 4573
rect 12256 4632 12308 4684
rect 12624 4632 12676 4684
rect 13084 4632 13136 4684
rect 16764 4709 16773 4743
rect 16773 4709 16807 4743
rect 16807 4709 16816 4743
rect 16764 4700 16816 4709
rect 16028 4632 16080 4684
rect 17960 4675 18012 4684
rect 17960 4641 17969 4675
rect 17969 4641 18003 4675
rect 18003 4641 18012 4675
rect 17960 4632 18012 4641
rect 14464 4607 14516 4616
rect 11060 4496 11112 4548
rect 9588 4428 9640 4480
rect 11796 4496 11848 4548
rect 12532 4428 12584 4480
rect 12900 4428 12952 4480
rect 14004 4539 14056 4548
rect 14004 4505 14013 4539
rect 14013 4505 14047 4539
rect 14047 4505 14056 4539
rect 14004 4496 14056 4505
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 14648 4607 14700 4616
rect 14648 4573 14657 4607
rect 14657 4573 14691 4607
rect 14691 4573 14700 4607
rect 14648 4564 14700 4573
rect 15568 4564 15620 4616
rect 15936 4564 15988 4616
rect 17408 4564 17460 4616
rect 14372 4428 14424 4480
rect 18788 4428 18840 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 1676 4088 1728 4140
rect 3332 4020 3384 4072
rect 6920 4224 6972 4276
rect 14648 4224 14700 4276
rect 4068 4131 4120 4140
rect 4068 4097 4077 4131
rect 4077 4097 4111 4131
rect 4111 4097 4120 4131
rect 4068 4088 4120 4097
rect 4344 4088 4396 4140
rect 8208 4156 8260 4208
rect 204 3952 256 4004
rect 4436 3952 4488 4004
rect 4712 4020 4764 4072
rect 7288 4063 7340 4072
rect 7288 4029 7297 4063
rect 7297 4029 7331 4063
rect 7331 4029 7340 4063
rect 7288 4020 7340 4029
rect 5448 3952 5500 4004
rect 6460 3952 6512 4004
rect 8300 4088 8352 4140
rect 8392 4088 8444 4140
rect 8944 4088 8996 4140
rect 10784 4156 10836 4208
rect 11060 4156 11112 4208
rect 12348 4156 12400 4208
rect 12440 4199 12492 4208
rect 12440 4165 12449 4199
rect 12449 4165 12483 4199
rect 12483 4165 12492 4199
rect 12440 4156 12492 4165
rect 12716 4156 12768 4208
rect 8576 4020 8628 4072
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 10968 4131 11020 4140
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 12900 4088 12952 4140
rect 13360 4156 13412 4208
rect 13912 4088 13964 4140
rect 2780 3884 2832 3936
rect 3608 3927 3660 3936
rect 3608 3893 3617 3927
rect 3617 3893 3651 3927
rect 3651 3893 3660 3927
rect 3608 3884 3660 3893
rect 6000 3927 6052 3936
rect 6000 3893 6009 3927
rect 6009 3893 6043 3927
rect 6043 3893 6052 3927
rect 6000 3884 6052 3893
rect 6276 3927 6328 3936
rect 6276 3893 6285 3927
rect 6285 3893 6319 3927
rect 6319 3893 6328 3927
rect 6276 3884 6328 3893
rect 7104 3884 7156 3936
rect 10232 3952 10284 4004
rect 8208 3884 8260 3936
rect 9772 3884 9824 3936
rect 9956 3884 10008 3936
rect 10416 3927 10468 3936
rect 10416 3893 10425 3927
rect 10425 3893 10459 3927
rect 10459 3893 10468 3927
rect 10416 3884 10468 3893
rect 10968 3952 11020 4004
rect 11152 3884 11204 3936
rect 11336 3952 11388 4004
rect 13176 4020 13228 4072
rect 14648 4088 14700 4140
rect 15936 4156 15988 4208
rect 16580 4156 16632 4208
rect 13912 3952 13964 4004
rect 14648 3995 14700 4004
rect 12348 3884 12400 3936
rect 12624 3884 12676 3936
rect 12992 3884 13044 3936
rect 13360 3884 13412 3936
rect 13820 3884 13872 3936
rect 14648 3961 14657 3995
rect 14657 3961 14691 3995
rect 14691 3961 14700 3995
rect 14648 3952 14700 3961
rect 14372 3884 14424 3936
rect 15936 4020 15988 4072
rect 16212 4063 16264 4072
rect 16212 4029 16221 4063
rect 16221 4029 16255 4063
rect 16255 4029 16264 4063
rect 16212 4020 16264 4029
rect 15108 3952 15160 4004
rect 15200 3927 15252 3936
rect 15200 3893 15209 3927
rect 15209 3893 15243 3927
rect 15243 3893 15252 3927
rect 15200 3884 15252 3893
rect 15568 3927 15620 3936
rect 15568 3893 15577 3927
rect 15577 3893 15611 3927
rect 15611 3893 15620 3927
rect 15568 3884 15620 3893
rect 15752 3884 15804 3936
rect 16764 3884 16816 3936
rect 22468 3884 22520 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 1584 3680 1636 3732
rect 6276 3680 6328 3732
rect 7748 3680 7800 3732
rect 8392 3723 8444 3732
rect 8392 3689 8401 3723
rect 8401 3689 8435 3723
rect 8435 3689 8444 3723
rect 8392 3680 8444 3689
rect 8576 3680 8628 3732
rect 9128 3680 9180 3732
rect 9496 3680 9548 3732
rect 9956 3680 10008 3732
rect 10600 3680 10652 3732
rect 10968 3680 11020 3732
rect 1124 3476 1176 3528
rect 2320 3587 2372 3596
rect 2320 3553 2329 3587
rect 2329 3553 2363 3587
rect 2363 3553 2372 3587
rect 2320 3544 2372 3553
rect 4160 3612 4212 3664
rect 7104 3612 7156 3664
rect 3148 3544 3200 3596
rect 3424 3587 3476 3596
rect 3424 3553 3433 3587
rect 3433 3553 3467 3587
rect 3467 3553 3476 3587
rect 3424 3544 3476 3553
rect 2504 3476 2556 3528
rect 2964 3476 3016 3528
rect 3516 3519 3568 3528
rect 3516 3485 3525 3519
rect 3525 3485 3559 3519
rect 3559 3485 3568 3519
rect 6000 3544 6052 3596
rect 7748 3544 7800 3596
rect 9036 3587 9088 3596
rect 9036 3553 9045 3587
rect 9045 3553 9079 3587
rect 9079 3553 9088 3587
rect 9036 3544 9088 3553
rect 9680 3544 9732 3596
rect 10416 3612 10468 3664
rect 11060 3612 11112 3664
rect 11152 3612 11204 3664
rect 12808 3680 12860 3732
rect 13084 3680 13136 3732
rect 13268 3612 13320 3664
rect 13452 3612 13504 3664
rect 13728 3612 13780 3664
rect 14372 3680 14424 3732
rect 16304 3680 16356 3732
rect 15936 3612 15988 3664
rect 4160 3519 4212 3528
rect 3516 3476 3568 3485
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 6460 3519 6512 3528
rect 664 3408 716 3460
rect 4068 3340 4120 3392
rect 5448 3408 5500 3460
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 6552 3476 6604 3528
rect 7012 3519 7064 3528
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 7012 3476 7064 3485
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 11520 3519 11572 3528
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11520 3476 11572 3485
rect 13360 3476 13412 3528
rect 14188 3544 14240 3596
rect 14280 3544 14332 3596
rect 15200 3544 15252 3596
rect 16672 3544 16724 3596
rect 14464 3476 14516 3528
rect 7748 3340 7800 3392
rect 12164 3340 12216 3392
rect 12440 3340 12492 3392
rect 12624 3340 12676 3392
rect 14556 3408 14608 3460
rect 20168 3476 20220 3528
rect 17408 3408 17460 3460
rect 16948 3340 17000 3392
rect 17316 3383 17368 3392
rect 17316 3349 17325 3383
rect 17325 3349 17359 3383
rect 17359 3349 17368 3383
rect 17316 3340 17368 3349
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 9680 3179 9732 3188
rect 5264 3068 5316 3120
rect 7012 3068 7064 3120
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 2688 2864 2740 2916
rect 2964 3043 3016 3052
rect 2964 3009 2973 3043
rect 2973 3009 3007 3043
rect 3007 3009 3016 3043
rect 2964 3000 3016 3009
rect 5448 3000 5500 3052
rect 6552 3000 6604 3052
rect 7748 3043 7800 3052
rect 7748 3009 7757 3043
rect 7757 3009 7791 3043
rect 7791 3009 7800 3043
rect 7748 3000 7800 3009
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 12624 3136 12676 3188
rect 12808 3136 12860 3188
rect 9864 3068 9916 3120
rect 10048 3068 10100 3120
rect 11796 3068 11848 3120
rect 10324 3000 10376 3052
rect 10600 3000 10652 3052
rect 11152 3043 11204 3052
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 11336 3000 11388 3052
rect 12532 3000 12584 3052
rect 14372 3000 14424 3052
rect 14648 3000 14700 3052
rect 22008 3136 22060 3188
rect 19708 3068 19760 3120
rect 15568 3000 15620 3052
rect 3056 2932 3108 2984
rect 4068 2932 4120 2984
rect 6000 2932 6052 2984
rect 3424 2864 3476 2916
rect 5356 2864 5408 2916
rect 3516 2796 3568 2848
rect 4620 2796 4672 2848
rect 5172 2839 5224 2848
rect 5172 2805 5181 2839
rect 5181 2805 5215 2839
rect 5215 2805 5224 2839
rect 8392 2932 8444 2984
rect 9864 2932 9916 2984
rect 10140 2932 10192 2984
rect 10876 2975 10928 2984
rect 10876 2941 10885 2975
rect 10885 2941 10919 2975
rect 10919 2941 10928 2975
rect 10876 2932 10928 2941
rect 11612 2975 11664 2984
rect 11612 2941 11621 2975
rect 11621 2941 11655 2975
rect 11655 2941 11664 2975
rect 11612 2932 11664 2941
rect 12072 2932 12124 2984
rect 14004 2932 14056 2984
rect 15476 2975 15528 2984
rect 15476 2941 15485 2975
rect 15485 2941 15519 2975
rect 15519 2941 15528 2975
rect 15476 2932 15528 2941
rect 16396 2975 16448 2984
rect 16396 2941 16405 2975
rect 16405 2941 16439 2975
rect 16439 2941 16448 2975
rect 16396 2932 16448 2941
rect 9036 2864 9088 2916
rect 12624 2864 12676 2916
rect 5172 2796 5224 2805
rect 6092 2839 6144 2848
rect 6092 2805 6101 2839
rect 6101 2805 6135 2839
rect 6135 2805 6144 2839
rect 6092 2796 6144 2805
rect 8300 2796 8352 2848
rect 8668 2796 8720 2848
rect 10140 2796 10192 2848
rect 13268 2796 13320 2848
rect 14372 2864 14424 2916
rect 14464 2796 14516 2848
rect 15200 2796 15252 2848
rect 16120 2796 16172 2848
rect 17776 2864 17828 2916
rect 21548 2864 21600 2916
rect 17868 2796 17920 2848
rect 19248 2796 19300 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 2320 2592 2372 2644
rect 2688 2592 2740 2644
rect 3332 2592 3384 2644
rect 5172 2592 5224 2644
rect 5356 2592 5408 2644
rect 5816 2592 5868 2644
rect 8668 2592 8720 2644
rect 10232 2635 10284 2644
rect 10232 2601 10241 2635
rect 10241 2601 10275 2635
rect 10275 2601 10284 2635
rect 10232 2592 10284 2601
rect 10876 2592 10928 2644
rect 11060 2592 11112 2644
rect 11336 2592 11388 2644
rect 14188 2592 14240 2644
rect 14464 2592 14516 2644
rect 3700 2524 3752 2576
rect 5080 2524 5132 2576
rect 8300 2524 8352 2576
rect 9772 2524 9824 2576
rect 11612 2524 11664 2576
rect 13452 2524 13504 2576
rect 15476 2592 15528 2644
rect 17776 2592 17828 2644
rect 2688 2456 2740 2508
rect 3332 2499 3384 2508
rect 3332 2465 3341 2499
rect 3341 2465 3375 2499
rect 3375 2465 3384 2499
rect 3332 2456 3384 2465
rect 2412 2431 2464 2440
rect 2412 2397 2421 2431
rect 2421 2397 2455 2431
rect 2455 2397 2464 2431
rect 2412 2388 2464 2397
rect 2780 2388 2832 2440
rect 3424 2388 3476 2440
rect 4160 2388 4212 2440
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 7564 2431 7616 2440
rect 7564 2397 7573 2431
rect 7573 2397 7607 2431
rect 7607 2397 7616 2431
rect 7564 2388 7616 2397
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 5080 2295 5132 2304
rect 5080 2261 5089 2295
rect 5089 2261 5123 2295
rect 5123 2261 5132 2295
rect 5080 2252 5132 2261
rect 5448 2320 5500 2372
rect 8116 2320 8168 2372
rect 10600 2456 10652 2508
rect 10784 2456 10836 2508
rect 11796 2499 11848 2508
rect 9680 2388 9732 2440
rect 11796 2465 11805 2499
rect 11805 2465 11839 2499
rect 11839 2465 11848 2499
rect 11796 2456 11848 2465
rect 11980 2456 12032 2508
rect 13176 2431 13228 2440
rect 13176 2397 13185 2431
rect 13185 2397 13219 2431
rect 13219 2397 13228 2431
rect 13176 2388 13228 2397
rect 13360 2456 13412 2508
rect 14188 2431 14240 2440
rect 14188 2397 14197 2431
rect 14197 2397 14231 2431
rect 14231 2397 14240 2431
rect 14188 2388 14240 2397
rect 15844 2456 15896 2508
rect 16120 2456 16172 2508
rect 17500 2499 17552 2508
rect 17500 2465 17509 2499
rect 17509 2465 17543 2499
rect 17543 2465 17552 2499
rect 17500 2456 17552 2465
rect 16856 2388 16908 2440
rect 5632 2252 5684 2304
rect 12624 2295 12676 2304
rect 12624 2261 12633 2295
rect 12633 2261 12667 2295
rect 12667 2261 12676 2295
rect 12624 2252 12676 2261
rect 15108 2320 15160 2372
rect 16028 2320 16080 2372
rect 16488 2252 16540 2304
rect 17960 2252 18012 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 2412 2048 2464 2100
rect 13268 2048 13320 2100
rect 15476 2048 15528 2100
rect 21088 2048 21140 2100
rect 2688 1980 2740 2032
rect 5080 1980 5132 2032
rect 14372 1980 14424 2032
rect 13912 1912 13964 1964
rect 14096 1912 14148 1964
rect 16580 1912 16632 1964
rect 2504 1844 2556 1896
rect 12624 1844 12676 1896
rect 2964 1776 3016 1828
rect 4896 1776 4948 1828
rect 3516 1708 3568 1760
rect 11612 1776 11664 1828
rect 5632 1708 5684 1760
rect 6644 1708 6696 1760
rect 3424 1640 3476 1692
rect 13176 1708 13228 1760
rect 14556 1708 14608 1760
rect 17316 1708 17368 1760
rect 8116 1640 8168 1692
rect 8760 1640 8812 1692
rect 9312 1640 9364 1692
rect 13360 1640 13412 1692
rect 2504 1572 2556 1624
rect 7564 1572 7616 1624
rect 12164 1572 12216 1624
rect 13176 1572 13228 1624
rect 3424 1504 3476 1556
rect 9312 1504 9364 1556
rect 1584 1436 1636 1488
rect 6000 1436 6052 1488
rect 2044 1368 2096 1420
rect 6092 1368 6144 1420
rect 11336 1368 11388 1420
rect 12348 1368 12400 1420
rect 4068 1300 4120 1352
rect 14280 1300 14332 1352
rect 3976 1164 4028 1216
rect 14004 1164 14056 1216
<< metal2 >>
rect 202 22320 258 22800
rect 662 22320 718 22800
rect 1122 22320 1178 22800
rect 1582 22320 1638 22800
rect 2042 22320 2098 22800
rect 2502 22320 2558 22800
rect 2962 22320 3018 22800
rect 3422 22320 3478 22800
rect 3514 22536 3570 22545
rect 3514 22471 3570 22480
rect 216 15026 244 22320
rect 204 15020 256 15026
rect 204 14962 256 14968
rect 676 14890 704 22320
rect 664 14884 716 14890
rect 664 14826 716 14832
rect 1136 14278 1164 22320
rect 1596 19394 1624 22320
rect 1676 19916 1728 19922
rect 1676 19858 1728 19864
rect 1504 19366 1624 19394
rect 1504 16096 1532 19366
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1596 17202 1624 19246
rect 1688 17882 1716 19858
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1768 19168 1820 19174
rect 1768 19110 1820 19116
rect 1780 18329 1808 19110
rect 1872 18737 1900 19654
rect 1858 18728 1914 18737
rect 1858 18663 1914 18672
rect 1766 18320 1822 18329
rect 1766 18255 1822 18264
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 1688 16833 1716 17478
rect 1780 17202 1808 18158
rect 2056 18086 2084 22320
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2516 20346 2544 22320
rect 2240 19922 2268 20334
rect 2516 20318 2636 20346
rect 2228 19916 2280 19922
rect 2228 19858 2280 19864
rect 2412 19236 2464 19242
rect 2412 19178 2464 19184
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2148 18834 2176 19110
rect 2318 19000 2374 19009
rect 2318 18935 2374 18944
rect 2136 18828 2188 18834
rect 2136 18770 2188 18776
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 2044 18080 2096 18086
rect 2044 18022 2096 18028
rect 1964 17377 1992 18022
rect 1950 17368 2006 17377
rect 1950 17303 2006 17312
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1674 16824 1730 16833
rect 1674 16759 1730 16768
rect 1676 16448 1728 16454
rect 1674 16416 1676 16425
rect 1728 16416 1730 16425
rect 1674 16351 1730 16360
rect 1504 16068 1808 16096
rect 1492 15972 1544 15978
rect 1492 15914 1544 15920
rect 1504 14958 1532 15914
rect 1582 15872 1638 15881
rect 1582 15807 1638 15816
rect 1596 15706 1624 15807
rect 1584 15700 1636 15706
rect 1584 15642 1636 15648
rect 1582 15464 1638 15473
rect 1582 15399 1638 15408
rect 1596 15162 1624 15399
rect 1584 15156 1636 15162
rect 1584 15098 1636 15104
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1492 14952 1544 14958
rect 1492 14894 1544 14900
rect 1582 14920 1638 14929
rect 1582 14855 1638 14864
rect 1124 14272 1176 14278
rect 1124 14214 1176 14220
rect 1136 13870 1164 14214
rect 1124 13864 1176 13870
rect 1124 13806 1176 13812
rect 1596 13530 1624 14855
rect 1688 13938 1716 14962
rect 1780 14550 1808 16068
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 1768 14544 1820 14550
rect 1768 14486 1820 14492
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1596 12986 1624 13330
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1872 12442 1900 15982
rect 2056 15706 2084 18022
rect 2332 17746 2360 18935
rect 2424 18873 2452 19178
rect 2410 18864 2466 18873
rect 2410 18799 2466 18808
rect 2504 18760 2556 18766
rect 2502 18728 2504 18737
rect 2556 18728 2558 18737
rect 2502 18663 2558 18672
rect 2608 18329 2636 20318
rect 2872 20324 2924 20330
rect 2872 20266 2924 20272
rect 2884 19990 2912 20266
rect 2872 19984 2924 19990
rect 2872 19926 2924 19932
rect 2976 19802 3004 22320
rect 3330 22128 3386 22137
rect 3330 22063 3386 22072
rect 3344 20738 3372 22063
rect 3332 20732 3384 20738
rect 3332 20674 3384 20680
rect 3330 20632 3386 20641
rect 3330 20567 3386 20576
rect 3344 20466 3372 20567
rect 3332 20460 3384 20466
rect 3332 20402 3384 20408
rect 3436 20074 3464 22320
rect 3528 20874 3556 22471
rect 3882 22320 3938 22800
rect 4342 22320 4398 22800
rect 4802 22320 4858 22800
rect 5262 22320 5318 22800
rect 5722 22320 5778 22800
rect 6182 22320 6238 22800
rect 6642 22320 6698 22800
rect 7102 22320 7158 22800
rect 7562 22320 7618 22800
rect 8114 22320 8170 22800
rect 8574 22320 8630 22800
rect 9034 22320 9090 22800
rect 9494 22320 9550 22800
rect 9954 22320 10010 22800
rect 10414 22320 10470 22800
rect 10874 22320 10930 22800
rect 11334 22320 11390 22800
rect 11794 22320 11850 22800
rect 12254 22320 12310 22800
rect 12714 22320 12770 22800
rect 13174 22320 13230 22800
rect 13634 22320 13690 22800
rect 14094 22320 14150 22800
rect 14554 22320 14610 22800
rect 15014 22320 15070 22800
rect 15566 22320 15622 22800
rect 16026 22320 16082 22800
rect 16486 22320 16542 22800
rect 16946 22320 17002 22800
rect 17406 22320 17462 22800
rect 17866 22320 17922 22800
rect 18326 22320 18382 22800
rect 18786 22320 18842 22800
rect 19246 22320 19302 22800
rect 19706 22320 19762 22800
rect 20166 22320 20222 22800
rect 20626 22320 20682 22800
rect 21086 22320 21142 22800
rect 21546 22320 21602 22800
rect 22006 22320 22062 22800
rect 22466 22320 22522 22800
rect 3516 20868 3568 20874
rect 3516 20810 3568 20816
rect 3436 20046 3740 20074
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 2884 19774 3004 19802
rect 2594 18320 2650 18329
rect 2594 18255 2650 18264
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 2228 17128 2280 17134
rect 2228 17070 2280 17076
rect 2240 16794 2268 17070
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2320 16652 2372 16658
rect 2320 16594 2372 16600
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 2056 13938 2084 15438
rect 2136 14952 2188 14958
rect 2136 14894 2188 14900
rect 2148 13938 2176 14894
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2056 13705 2084 13874
rect 2042 13696 2098 13705
rect 2042 13631 2098 13640
rect 2240 13462 2268 16526
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1412 11286 1440 11630
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1400 11280 1452 11286
rect 1400 11222 1452 11228
rect 1504 8430 1532 11494
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 204 4004 256 4010
rect 204 3946 256 3952
rect 216 480 244 3946
rect 1596 3738 1624 11154
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1688 10470 1716 11086
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 10062 1716 10406
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1688 9518 1716 9998
rect 1676 9512 1728 9518
rect 1872 9489 1900 12242
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1964 11801 1992 12174
rect 1950 11792 2006 11801
rect 1950 11727 2006 11736
rect 2056 10713 2084 12582
rect 2042 10704 2098 10713
rect 2042 10639 2098 10648
rect 2332 9738 2360 16594
rect 2700 16046 2728 18158
rect 2778 16824 2834 16833
rect 2778 16759 2834 16768
rect 2792 16726 2820 16759
rect 2780 16720 2832 16726
rect 2780 16662 2832 16668
rect 2688 16040 2740 16046
rect 2688 15982 2740 15988
rect 2884 15570 2912 19774
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 2976 18834 3004 19654
rect 3056 19236 3108 19242
rect 3056 19178 3108 19184
rect 2964 18828 3016 18834
rect 2964 18770 3016 18776
rect 3068 18426 3096 19178
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3344 18970 3372 19110
rect 3332 18964 3384 18970
rect 3332 18906 3384 18912
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 2976 17678 3004 17818
rect 3240 17740 3292 17746
rect 3240 17682 3292 17688
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 3068 16726 3096 17546
rect 3252 17202 3280 17682
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3056 16720 3108 16726
rect 3056 16662 3108 16668
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2976 15706 3004 16594
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 3344 15706 3372 15846
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 2872 15564 2924 15570
rect 2872 15506 2924 15512
rect 2884 15162 2912 15506
rect 3436 15502 3464 18702
rect 3528 18222 3556 18702
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3528 17785 3556 17818
rect 3514 17776 3570 17785
rect 3514 17711 3570 17720
rect 3620 17678 3648 19858
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2608 14793 2636 14962
rect 2964 14952 3016 14958
rect 2962 14920 2964 14929
rect 3016 14920 3018 14929
rect 2962 14855 3018 14864
rect 2964 14816 3016 14822
rect 2594 14784 2650 14793
rect 2964 14758 3016 14764
rect 2594 14719 2650 14728
rect 2778 14512 2834 14521
rect 2504 14476 2556 14482
rect 2778 14447 2834 14456
rect 2504 14418 2556 14424
rect 2412 14408 2464 14414
rect 2516 14385 2544 14418
rect 2688 14408 2740 14414
rect 2412 14350 2464 14356
rect 2502 14376 2558 14385
rect 2424 12986 2452 14350
rect 2688 14350 2740 14356
rect 2502 14311 2558 14320
rect 2700 13802 2728 14350
rect 2688 13796 2740 13802
rect 2688 13738 2740 13744
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2412 12980 2464 12986
rect 2412 12922 2464 12928
rect 2516 12442 2544 13262
rect 2700 12918 2728 13738
rect 2688 12912 2740 12918
rect 2688 12854 2740 12860
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 2700 12442 2728 12718
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2792 11898 2820 14447
rect 2870 13968 2926 13977
rect 2870 13903 2926 13912
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2424 10810 2452 11698
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2424 10130 2452 10746
rect 2884 10266 2912 13903
rect 2976 13841 3004 14758
rect 2962 13832 3018 13841
rect 2962 13767 3018 13776
rect 2964 13728 3016 13734
rect 2962 13696 2964 13705
rect 3016 13696 3018 13705
rect 2962 13631 3018 13640
rect 2976 12850 3004 13631
rect 3068 13394 3096 15302
rect 3332 14884 3384 14890
rect 3332 14826 3384 14832
rect 3344 14770 3372 14826
rect 3160 14742 3372 14770
rect 3160 14618 3188 14742
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3238 13560 3294 13569
rect 3238 13495 3294 13504
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 3252 12850 3280 13495
rect 3436 13462 3464 14010
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3240 12708 3292 12714
rect 3240 12650 3292 12656
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2332 9710 2636 9738
rect 1950 9616 2006 9625
rect 1950 9551 2006 9560
rect 2320 9580 2372 9586
rect 1676 9454 1728 9460
rect 1858 9480 1914 9489
rect 1688 8430 1716 9454
rect 1858 9415 1914 9424
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1872 9178 1900 9318
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1964 8974 1992 9551
rect 2320 9522 2372 9528
rect 2134 9344 2190 9353
rect 2134 9279 2190 9288
rect 2148 9110 2176 9279
rect 2136 9104 2188 9110
rect 2136 9046 2188 9052
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1688 7750 1716 8366
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 7342 1716 7686
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1688 6254 1716 7278
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1688 4690 1716 6190
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1872 5370 1900 5714
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1688 4146 1716 4626
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1124 3528 1176 3534
rect 1124 3470 1176 3476
rect 664 3460 716 3466
rect 664 3402 716 3408
rect 676 480 704 3402
rect 1136 480 1164 3470
rect 1964 1601 1992 8910
rect 2148 2553 2176 9046
rect 2332 8922 2360 9522
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 2516 9178 2544 9386
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2332 8906 2452 8922
rect 2332 8900 2464 8906
rect 2332 8894 2412 8900
rect 2412 8842 2464 8848
rect 2424 8634 2452 8842
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2424 8022 2452 8570
rect 2412 8016 2464 8022
rect 2412 7958 2464 7964
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 2332 5166 2360 5510
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2226 4176 2282 4185
rect 2226 4111 2282 4120
rect 2240 3097 2268 4111
rect 2410 3768 2466 3777
rect 2410 3703 2466 3712
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 2226 3088 2282 3097
rect 2226 3023 2282 3032
rect 2332 2650 2360 3538
rect 2424 3058 2452 3703
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2134 2544 2190 2553
rect 2134 2479 2190 2488
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 2424 2106 2452 2382
rect 2412 2100 2464 2106
rect 2412 2042 2464 2048
rect 2516 1902 2544 3470
rect 2608 3097 2636 9710
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2792 7274 2820 9590
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 8430 2912 8910
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2884 7342 2912 7686
rect 2872 7336 2924 7342
rect 2976 7313 3004 12310
rect 3056 12232 3108 12238
rect 3108 12192 3188 12220
rect 3252 12209 3280 12650
rect 3436 12646 3464 13262
rect 3528 13190 3556 16934
rect 3608 15972 3660 15978
rect 3608 15914 3660 15920
rect 3620 15609 3648 15914
rect 3606 15600 3662 15609
rect 3606 15535 3662 15544
rect 3620 15502 3648 15535
rect 3608 15496 3660 15502
rect 3608 15438 3660 15444
rect 3712 15366 3740 20046
rect 3700 15360 3752 15366
rect 3700 15302 3752 15308
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3606 14648 3662 14657
rect 3606 14583 3662 14592
rect 3620 14414 3648 14583
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 3608 14408 3660 14414
rect 3608 14350 3660 14356
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3620 13802 3648 14214
rect 3608 13796 3660 13802
rect 3608 13738 3660 13744
rect 3620 13326 3648 13738
rect 3712 13734 3740 14418
rect 3804 13734 3832 14758
rect 3700 13728 3752 13734
rect 3700 13670 3752 13676
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3804 13326 3832 13670
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3056 12174 3108 12180
rect 3056 11620 3108 11626
rect 3056 11562 3108 11568
rect 3068 10810 3096 11562
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3160 10010 3188 12192
rect 3238 12200 3294 12209
rect 3238 12135 3294 12144
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3344 11354 3372 11494
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3238 10704 3294 10713
rect 3238 10639 3294 10648
rect 3068 9982 3188 10010
rect 2872 7278 2924 7284
rect 2962 7304 3018 7313
rect 2780 7268 2832 7274
rect 2962 7239 3018 7248
rect 2780 7210 2832 7216
rect 2976 6798 3004 7239
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 3068 5642 3096 9982
rect 3252 9926 3280 10639
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3160 8974 3188 9862
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3252 7002 3280 9386
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3344 8090 3372 8910
rect 3528 8362 3556 12854
rect 3620 12238 3648 13262
rect 3700 12980 3752 12986
rect 3700 12922 3752 12928
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3620 10996 3648 11698
rect 3712 11694 3740 12922
rect 3896 12714 3924 22320
rect 4066 21584 4122 21593
rect 4066 21519 4122 21528
rect 3974 21176 4030 21185
rect 4080 21146 4108 21519
rect 3974 21111 4030 21120
rect 4068 21140 4120 21146
rect 3988 21010 4016 21111
rect 4068 21082 4120 21088
rect 3976 21004 4028 21010
rect 3976 20946 4028 20952
rect 4068 20256 4120 20262
rect 4066 20224 4068 20233
rect 4120 20224 4122 20233
rect 4066 20159 4122 20168
rect 4356 19802 4384 22320
rect 4264 19774 4384 19802
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4160 19712 4212 19718
rect 4066 19680 4122 19689
rect 4160 19654 4212 19660
rect 4066 19615 4122 19624
rect 4080 19514 4108 19615
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 4172 19394 4200 19654
rect 3988 19366 4200 19394
rect 4264 19394 4292 19774
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4264 19366 4476 19394
rect 3988 19310 4016 19366
rect 3976 19304 4028 19310
rect 4252 19304 4304 19310
rect 3976 19246 4028 19252
rect 4066 19272 4122 19281
rect 4122 19230 4200 19258
rect 4252 19246 4304 19252
rect 4066 19207 4122 19216
rect 4172 19174 4200 19230
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 4080 18766 4108 19110
rect 4264 18902 4292 19246
rect 4448 18902 4476 19366
rect 4252 18896 4304 18902
rect 4252 18838 4304 18844
rect 4436 18896 4488 18902
rect 4436 18838 4488 18844
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 4080 18154 4108 18702
rect 4264 18426 4292 18838
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 4724 17882 4752 19790
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 3976 16516 4028 16522
rect 3976 16458 4028 16464
rect 3988 16046 4016 16458
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 3988 13190 4016 14554
rect 4080 13258 4108 17070
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4172 16250 4200 16594
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 4172 14929 4200 15982
rect 4264 15162 4292 17138
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4158 14920 4214 14929
rect 4158 14855 4214 14864
rect 4172 14822 4200 14855
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4160 14340 4212 14346
rect 4160 14282 4212 14288
rect 4172 13462 4200 14282
rect 4264 13938 4292 15098
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4356 14414 4384 14758
rect 4724 14618 4752 14758
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4356 14260 4384 14350
rect 4325 14232 4384 14260
rect 4325 14056 4353 14232
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4325 14028 4384 14056
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4252 13796 4304 13802
rect 4356 13784 4384 14028
rect 4304 13756 4384 13784
rect 4252 13738 4304 13744
rect 4160 13456 4212 13462
rect 4160 13398 4212 13404
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3988 12617 4016 12922
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3974 12608 4030 12617
rect 3974 12543 4030 12552
rect 3974 12064 4030 12073
rect 3974 11999 4030 12008
rect 3988 11898 4016 11999
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3882 11656 3938 11665
rect 3700 11008 3752 11014
rect 3620 10968 3700 10996
rect 3700 10950 3752 10956
rect 3712 10674 3740 10950
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3516 8356 3568 8362
rect 3516 8298 3568 8304
rect 3620 8242 3648 8910
rect 3528 8214 3648 8242
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 3160 6458 3188 6802
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3160 5710 3188 6394
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2792 3942 2820 4626
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2594 3088 2650 3097
rect 2594 3023 2650 3032
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 2700 2650 2728 2858
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 2700 2038 2728 2450
rect 2792 2446 2820 3878
rect 2976 3534 3004 4422
rect 3068 4049 3096 5578
rect 3160 5234 3188 5646
rect 3252 5370 3280 6938
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3054 4040 3110 4049
rect 3054 3975 3110 3984
rect 3160 3602 3188 4626
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 2964 3528 3016 3534
rect 3016 3488 3096 3516
rect 2964 3470 3016 3476
rect 2962 3224 3018 3233
rect 2962 3159 3018 3168
rect 2976 3058 3004 3159
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 3068 2990 3096 3488
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 3252 2496 3280 4966
rect 3344 4078 3372 7142
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 5914 3464 6054
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3424 4616 3476 4622
rect 3422 4584 3424 4593
rect 3476 4584 3478 4593
rect 3422 4519 3478 4528
rect 3528 4468 3556 8214
rect 3804 7546 3832 11630
rect 3882 11591 3884 11600
rect 3936 11591 3938 11600
rect 3884 11562 3936 11568
rect 4080 11150 4108 12786
rect 4264 12374 4292 13738
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4724 12646 4752 13466
rect 4816 12714 4844 22320
rect 4988 20460 5040 20466
rect 4988 20402 5040 20408
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4908 19174 4936 19790
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4908 18154 4936 19110
rect 4896 18148 4948 18154
rect 4896 18090 4948 18096
rect 5000 15910 5028 20402
rect 5276 20058 5304 22320
rect 5736 20466 5764 22320
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5172 20052 5224 20058
rect 5172 19994 5224 20000
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 5184 19786 5212 19994
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 5172 19780 5224 19786
rect 5172 19722 5224 19728
rect 5644 19446 5672 19858
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 5632 19440 5684 19446
rect 5632 19382 5684 19388
rect 5448 19236 5500 19242
rect 5448 19178 5500 19184
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5368 18222 5396 18702
rect 5460 18698 5488 19178
rect 5448 18692 5500 18698
rect 5448 18634 5500 18640
rect 5356 18216 5408 18222
rect 5356 18158 5408 18164
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 5092 15706 5120 16934
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 4988 15564 5040 15570
rect 4988 15506 5040 15512
rect 4896 15428 4948 15434
rect 4896 15370 4948 15376
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4712 12640 4764 12646
rect 4816 12617 4844 12650
rect 4712 12582 4764 12588
rect 4802 12608 4858 12617
rect 4802 12543 4858 12552
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4804 11688 4856 11694
rect 4618 11656 4674 11665
rect 4252 11620 4304 11626
rect 4804 11630 4856 11636
rect 4618 11591 4674 11600
rect 4252 11562 4304 11568
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 10606 4108 10950
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4264 10198 4292 11562
rect 4632 11286 4660 11591
rect 4620 11280 4672 11286
rect 4620 11222 4672 11228
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4724 10674 4752 11018
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4080 9761 4108 9998
rect 4356 9908 4384 10542
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4448 10266 4476 10406
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4325 9880 4384 9908
rect 4066 9752 4122 9761
rect 4066 9687 4122 9696
rect 4325 9704 4353 9880
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4724 9722 4752 10610
rect 4816 9994 4844 11630
rect 4908 11218 4936 15370
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4804 9988 4856 9994
rect 4804 9930 4856 9936
rect 4712 9716 4764 9722
rect 4325 9676 4568 9704
rect 4252 9104 4304 9110
rect 4252 9046 4304 9052
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 3896 8634 3924 8978
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 3976 8832 4028 8838
rect 4080 8809 4108 8842
rect 3976 8774 4028 8780
rect 4066 8800 4122 8809
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3606 6896 3662 6905
rect 3606 6831 3662 6840
rect 3620 6118 3648 6831
rect 3792 6724 3844 6730
rect 3792 6666 3844 6672
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3712 6254 3740 6598
rect 3804 6361 3832 6666
rect 3790 6352 3846 6361
rect 3790 6287 3846 6296
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3436 4440 3556 4468
rect 3804 4457 3832 5306
rect 3790 4448 3846 4457
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3436 3602 3464 4440
rect 3790 4383 3846 4392
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3436 3505 3464 3538
rect 3516 3528 3568 3534
rect 3422 3496 3478 3505
rect 3516 3470 3568 3476
rect 3422 3431 3478 3440
rect 3424 2916 3476 2922
rect 3344 2876 3424 2904
rect 3344 2650 3372 2876
rect 3424 2858 3476 2864
rect 3528 2854 3556 3470
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3620 2666 3648 3878
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3528 2638 3648 2666
rect 3332 2508 3384 2514
rect 3252 2468 3332 2496
rect 3332 2450 3384 2456
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2688 2032 2740 2038
rect 2688 1974 2740 1980
rect 2504 1896 2556 1902
rect 2504 1838 2556 1844
rect 2964 1828 3016 1834
rect 2964 1770 3016 1776
rect 2504 1624 2556 1630
rect 1950 1592 2006 1601
rect 2504 1566 2556 1572
rect 1950 1527 2006 1536
rect 1584 1488 1636 1494
rect 1584 1430 1636 1436
rect 1596 480 1624 1430
rect 2044 1420 2096 1426
rect 2044 1362 2096 1368
rect 2056 480 2084 1362
rect 2516 480 2544 1566
rect 2976 480 3004 1770
rect 3344 649 3372 2450
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 3436 1698 3464 2382
rect 3528 1766 3556 2638
rect 3700 2576 3752 2582
rect 3698 2544 3700 2553
rect 3752 2544 3754 2553
rect 3698 2479 3754 2488
rect 3516 1760 3568 1766
rect 3516 1702 3568 1708
rect 3424 1692 3476 1698
rect 3424 1634 3476 1640
rect 3424 1556 3476 1562
rect 3424 1498 3476 1504
rect 3330 640 3386 649
rect 3330 575 3386 584
rect 3436 480 3464 1498
rect 3896 480 3924 7890
rect 3988 7410 4016 8774
rect 4066 8735 4122 8744
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4080 7970 4108 8230
rect 4172 8090 4200 8978
rect 4264 8265 4292 9046
rect 4540 8945 4568 9676
rect 4712 9658 4764 9664
rect 4816 9654 4844 9930
rect 4804 9648 4856 9654
rect 4804 9590 4856 9596
rect 4712 8968 4764 8974
rect 4526 8936 4582 8945
rect 4712 8910 4764 8916
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4908 8922 4936 11154
rect 5000 10742 5028 15506
rect 5184 15434 5212 17682
rect 5460 17678 5488 18634
rect 5736 18358 5764 19450
rect 5816 19304 5868 19310
rect 5816 19246 5868 19252
rect 5828 19009 5856 19246
rect 5814 19000 5870 19009
rect 5814 18935 5870 18944
rect 6012 18902 6040 19790
rect 5816 18896 5868 18902
rect 5816 18838 5868 18844
rect 6000 18896 6052 18902
rect 6000 18838 6052 18844
rect 5724 18352 5776 18358
rect 5724 18294 5776 18300
rect 5540 18148 5592 18154
rect 5540 18090 5592 18096
rect 5552 17882 5580 18090
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5828 17814 5856 18838
rect 6012 18426 6040 18838
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 5816 17808 5868 17814
rect 5816 17750 5868 17756
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5460 15978 5488 16390
rect 5552 16046 5580 16526
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 5460 15502 5488 15914
rect 5644 15706 5672 16934
rect 5920 16726 5948 17138
rect 6196 17082 6224 22320
rect 6276 21140 6328 21146
rect 6276 21082 6328 21088
rect 6288 19174 6316 21082
rect 6460 20732 6512 20738
rect 6460 20674 6512 20680
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 6472 18630 6500 20674
rect 6368 18624 6420 18630
rect 6368 18566 6420 18572
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6380 18426 6408 18566
rect 6368 18420 6420 18426
rect 6368 18362 6420 18368
rect 6656 18306 6684 22320
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 6012 17054 6224 17082
rect 6288 18278 6684 18306
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 5920 16250 5948 16662
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5172 15428 5224 15434
rect 5172 15370 5224 15376
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5092 14822 5120 15302
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 5368 14657 5396 14962
rect 5354 14648 5410 14657
rect 5354 14583 5410 14592
rect 5170 13832 5226 13841
rect 5170 13767 5226 13776
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 5092 12714 5120 13126
rect 5184 12850 5212 13767
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5080 12708 5132 12714
rect 5080 12650 5132 12656
rect 5092 12481 5120 12650
rect 5078 12472 5134 12481
rect 5078 12407 5134 12416
rect 5184 11529 5212 12786
rect 5276 12306 5304 13194
rect 5264 12300 5316 12306
rect 5316 12260 5396 12288
rect 5264 12242 5316 12248
rect 5262 11928 5318 11937
rect 5262 11863 5318 11872
rect 5170 11520 5226 11529
rect 5170 11455 5226 11464
rect 5276 11286 5304 11863
rect 5264 11280 5316 11286
rect 5264 11222 5316 11228
rect 4988 10736 5040 10742
rect 4988 10678 5040 10684
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5092 10282 5120 10610
rect 5000 10266 5120 10282
rect 4988 10260 5120 10266
rect 5040 10254 5120 10260
rect 4988 10202 5040 10208
rect 5172 10192 5224 10198
rect 5172 10134 5224 10140
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 5000 9110 5028 10066
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 4526 8871 4582 8880
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4724 8498 4752 8910
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4250 8256 4306 8265
rect 4250 8191 4306 8200
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4080 7942 4200 7970
rect 4066 7848 4122 7857
rect 4066 7783 4122 7792
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 4080 7206 4108 7783
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3988 5953 4016 6394
rect 3974 5944 4030 5953
rect 3974 5879 4030 5888
rect 4080 5846 4108 6598
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 3974 5400 4030 5409
rect 3974 5335 4030 5344
rect 3988 4758 4016 5335
rect 4080 5166 4108 5510
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4172 5098 4200 7942
rect 4724 7886 4752 8434
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4264 5166 4292 6190
rect 4724 6186 4752 6734
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4724 5846 4752 6122
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4724 5710 4752 5782
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4826 4108 4966
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4080 3505 4108 4082
rect 4172 3670 4200 4626
rect 4632 4468 4660 5102
rect 4724 4622 4752 5646
rect 4816 5001 4844 8910
rect 4908 8894 5028 8922
rect 4802 4992 4858 5001
rect 4802 4927 4858 4936
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4632 4440 4752 4468
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 4160 3528 4212 3534
rect 4066 3496 4122 3505
rect 4356 3516 4384 4082
rect 4724 4078 4752 4440
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4436 4004 4488 4010
rect 4436 3946 4488 3952
rect 4212 3488 4384 3516
rect 4160 3470 4212 3476
rect 4066 3431 4122 3440
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4080 2990 4108 3334
rect 4172 3233 4200 3470
rect 4448 3380 4476 3946
rect 4264 3352 4476 3380
rect 4158 3224 4214 3233
rect 4158 3159 4214 3168
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4172 1601 4200 2382
rect 4158 1592 4214 1601
rect 4158 1527 4214 1536
rect 4264 1442 4292 3352
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4632 2446 4660 2790
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4264 1414 4384 1442
rect 4068 1352 4120 1358
rect 4068 1294 4120 1300
rect 3976 1216 4028 1222
rect 3974 1184 3976 1193
rect 4028 1184 4030 1193
rect 3974 1119 4030 1128
rect 202 0 258 480
rect 662 0 718 480
rect 1122 0 1178 480
rect 1582 0 1638 480
rect 2042 0 2098 480
rect 2502 0 2558 480
rect 2962 0 3018 480
rect 3422 0 3478 480
rect 3882 0 3938 480
rect 4080 241 4108 1294
rect 4356 480 4384 1414
rect 4816 480 4844 4762
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4908 2428 4936 4694
rect 5000 2938 5028 8894
rect 5092 7002 5120 9862
rect 5184 8974 5212 10134
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5170 8800 5226 8809
rect 5170 8735 5226 8744
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5184 3369 5212 8735
rect 5276 4826 5304 11222
rect 5368 10062 5396 12260
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5356 9376 5408 9382
rect 5460 9353 5488 15302
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5552 13394 5580 15030
rect 5632 14544 5684 14550
rect 5632 14486 5684 14492
rect 5644 13462 5672 14486
rect 6012 14362 6040 17054
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6104 16250 6132 16934
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6104 15706 6132 16050
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 6092 15564 6144 15570
rect 6092 15506 6144 15512
rect 6104 14550 6132 15506
rect 6092 14544 6144 14550
rect 6092 14486 6144 14492
rect 5920 14334 6040 14362
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5828 13462 5856 13670
rect 5632 13456 5684 13462
rect 5632 13398 5684 13404
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5828 12850 5856 13398
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5644 12442 5672 12582
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5552 10690 5580 11630
rect 5644 10810 5672 12242
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5736 11200 5764 12038
rect 5920 11642 5948 14334
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 6012 14074 6040 14214
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6196 13870 6224 15982
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6012 13326 6040 13670
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 6012 12374 6040 13262
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6104 12782 6132 13126
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 6012 11762 6040 12310
rect 6196 12102 6224 12786
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 6196 11694 6224 12038
rect 6184 11688 6236 11694
rect 5920 11614 6132 11642
rect 6184 11630 6236 11636
rect 5906 11520 5962 11529
rect 5906 11455 5962 11464
rect 5920 11286 5948 11455
rect 5908 11280 5960 11286
rect 5908 11222 5960 11228
rect 5736 11172 5856 11200
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5552 10674 5672 10690
rect 5552 10668 5684 10674
rect 5552 10662 5632 10668
rect 5632 10610 5684 10616
rect 5736 9518 5764 11018
rect 5828 10198 5856 11172
rect 5998 11112 6054 11121
rect 5998 11047 6054 11056
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5920 10470 5948 10950
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5828 9722 5856 10134
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5356 9318 5408 9324
rect 5446 9344 5502 9353
rect 5368 8294 5396 9318
rect 5446 9279 5502 9288
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5460 7546 5488 8570
rect 5630 8528 5686 8537
rect 5630 8463 5686 8472
rect 5644 8430 5672 8463
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5460 7342 5488 7482
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5460 6798 5488 7278
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5368 4758 5396 5714
rect 5460 5710 5488 6734
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5460 5166 5488 5646
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5552 4826 5580 5102
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5460 3466 5488 3946
rect 5644 3652 5672 8230
rect 5736 7342 5764 9454
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5828 7546 5856 7822
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5828 6934 5856 7482
rect 5920 7274 5948 7822
rect 6012 7410 6040 11047
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 6104 7290 6132 11614
rect 6288 11506 6316 18278
rect 6644 18216 6696 18222
rect 6644 18158 6696 18164
rect 6368 17740 6420 17746
rect 6368 17682 6420 17688
rect 6380 16454 6408 17682
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6196 11478 6316 11506
rect 6196 10146 6224 11478
rect 6196 10118 6316 10146
rect 6182 8528 6238 8537
rect 6182 8463 6238 8472
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 6012 7262 6132 7290
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 5816 6112 5868 6118
rect 5920 6100 5948 7210
rect 5868 6072 5948 6100
rect 5816 6054 5868 6060
rect 5828 5234 5856 6054
rect 6012 5930 6040 7262
rect 5920 5902 6040 5930
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5644 3624 5764 3652
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5170 3360 5226 3369
rect 5170 3295 5226 3304
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 5000 2910 5120 2938
rect 5092 2689 5120 2910
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5078 2680 5134 2689
rect 5184 2650 5212 2790
rect 5078 2615 5134 2624
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 5092 2428 5120 2518
rect 4908 2400 5120 2428
rect 4908 1834 4936 2400
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 5092 2038 5120 2246
rect 5080 2032 5132 2038
rect 5080 1974 5132 1980
rect 4896 1828 4948 1834
rect 4896 1770 4948 1776
rect 5276 480 5304 3062
rect 5460 3058 5488 3402
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 5368 2650 5396 2858
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5460 2378 5488 2994
rect 5630 2816 5686 2825
rect 5630 2751 5686 2760
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 5644 2310 5672 2751
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 5644 1766 5672 2246
rect 5632 1760 5684 1766
rect 5632 1702 5684 1708
rect 5736 480 5764 3624
rect 5920 3233 5948 5902
rect 6090 5672 6146 5681
rect 6090 5607 6146 5616
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 6012 3942 6040 5034
rect 6104 4622 6132 5607
rect 6196 5370 6224 8463
rect 6288 8294 6316 10118
rect 6380 9042 6408 16390
rect 6552 15904 6604 15910
rect 6472 15864 6552 15892
rect 6472 11336 6500 15864
rect 6552 15846 6604 15852
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6564 13734 6592 14418
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6656 12374 6684 18158
rect 6748 15910 6776 19382
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 6840 15314 6868 20402
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6932 19514 6960 20334
rect 7012 19916 7064 19922
rect 7012 19858 7064 19864
rect 6920 19508 6972 19514
rect 6920 19450 6972 19456
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6932 17882 6960 19246
rect 7024 18970 7052 19858
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7012 18692 7064 18698
rect 7012 18634 7064 18640
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6920 17672 6972 17678
rect 7024 17660 7052 18634
rect 7116 18154 7144 22320
rect 7380 20868 7432 20874
rect 7380 20810 7432 20816
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7300 18766 7328 19654
rect 7288 18760 7340 18766
rect 7208 18720 7288 18748
rect 7208 18358 7236 18720
rect 7288 18702 7340 18708
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7104 18148 7156 18154
rect 7104 18090 7156 18096
rect 7208 17746 7236 18294
rect 7392 17785 7420 20810
rect 7576 20346 7604 22320
rect 7484 20318 7604 20346
rect 7484 19310 7512 20318
rect 8128 20244 8156 22320
rect 8588 22250 8616 22320
rect 8588 22222 8800 22250
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 7576 20216 8156 20244
rect 7472 19304 7524 19310
rect 7472 19246 7524 19252
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7378 17776 7434 17785
rect 7196 17740 7248 17746
rect 7378 17711 7434 17720
rect 7196 17682 7248 17688
rect 6972 17632 7052 17660
rect 6920 17614 6972 17620
rect 7208 17524 7236 17682
rect 7024 17496 7236 17524
rect 6920 17128 6972 17134
rect 7024 17116 7052 17496
rect 6972 17088 7052 17116
rect 6920 17070 6972 17076
rect 6932 15978 6960 17070
rect 7104 17060 7156 17066
rect 7208 17048 7236 17496
rect 7288 17060 7340 17066
rect 7208 17020 7288 17048
rect 7104 17002 7156 17008
rect 7288 17002 7340 17008
rect 7116 16794 7144 17002
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7392 16794 7420 16934
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7116 16522 7144 16730
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7104 16516 7156 16522
rect 7104 16458 7156 16464
rect 7116 16114 7144 16458
rect 7392 16250 7420 16594
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6748 15286 6868 15314
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6656 11898 6684 12174
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6656 11762 6684 11834
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6472 11308 6592 11336
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6472 10674 6500 11154
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6564 10606 6592 11308
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6656 9654 6684 10950
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6748 9586 6776 15286
rect 6932 15178 6960 15914
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 6840 15150 6960 15178
rect 7024 15162 7052 15438
rect 7012 15156 7064 15162
rect 6840 14958 6868 15150
rect 7012 15098 7064 15104
rect 6828 14952 6880 14958
rect 6826 14920 6828 14929
rect 6920 14952 6972 14958
rect 6880 14920 6882 14929
rect 6920 14894 6972 14900
rect 6826 14855 6882 14864
rect 6932 14414 6960 14894
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 7300 14346 7328 15506
rect 7484 14618 7512 18022
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7576 14498 7604 20216
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7668 18902 7696 19654
rect 7748 19440 7800 19446
rect 7748 19382 7800 19388
rect 7656 18896 7708 18902
rect 7656 18838 7708 18844
rect 7760 18358 7788 19382
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 8022 18728 8078 18737
rect 8022 18663 8078 18672
rect 7748 18352 7800 18358
rect 7748 18294 7800 18300
rect 7838 18320 7894 18329
rect 7838 18255 7840 18264
rect 7892 18255 7894 18264
rect 7840 18226 7892 18232
rect 8036 18154 8064 18663
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 8128 18193 8156 18226
rect 8114 18184 8170 18193
rect 8024 18148 8076 18154
rect 8114 18119 8170 18128
rect 8024 18090 8076 18096
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7668 16833 7696 16934
rect 7654 16824 7710 16833
rect 7654 16759 7710 16768
rect 7760 15162 7788 18022
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8220 17898 8248 20946
rect 8668 20868 8720 20874
rect 8668 20810 8720 20816
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 8312 18970 8340 19314
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8298 18864 8354 18873
rect 8298 18799 8354 18808
rect 8312 18086 8340 18799
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8220 17870 8340 17898
rect 7840 17808 7892 17814
rect 7838 17776 7840 17785
rect 7892 17776 7894 17785
rect 7838 17711 7894 17720
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 8220 17338 8248 17682
rect 8312 17542 8340 17870
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7838 16688 7894 16697
rect 7838 16623 7894 16632
rect 7852 16590 7880 16623
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 8404 16182 8432 19654
rect 8680 19496 8708 20810
rect 8671 19468 8708 19496
rect 8671 19428 8699 19468
rect 8671 19400 8708 19428
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8496 18698 8524 19110
rect 8484 18692 8536 18698
rect 8484 18634 8536 18640
rect 8482 18184 8538 18193
rect 8482 18119 8538 18128
rect 8392 16176 8444 16182
rect 8392 16118 8444 16124
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 7840 15496 7892 15502
rect 7838 15464 7840 15473
rect 7892 15464 7894 15473
rect 7838 15399 7894 15408
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7852 15042 7880 15399
rect 8220 15162 8248 15506
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 7760 15014 7880 15042
rect 7656 14952 7708 14958
rect 7760 14929 7788 15014
rect 7656 14894 7708 14900
rect 7746 14920 7802 14929
rect 7668 14618 7696 14894
rect 7746 14855 7802 14864
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7484 14470 7604 14498
rect 7288 14340 7340 14346
rect 7288 14282 7340 14288
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6932 11744 6960 13942
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 6932 11716 7052 11744
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6932 11218 6960 11562
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6828 9648 6880 9654
rect 6826 9616 6828 9625
rect 6880 9616 6882 9625
rect 6736 9580 6788 9586
rect 6826 9551 6882 9560
rect 6736 9522 6788 9528
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6472 8634 6500 9386
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6276 7948 6328 7954
rect 6564 7936 6592 8230
rect 6656 8090 6684 8774
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6564 7908 6684 7936
rect 6276 7890 6328 7896
rect 6288 5370 6316 7890
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6472 6866 6500 7142
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6564 4826 6592 5034
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 6012 3602 6040 3878
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 5906 3224 5962 3233
rect 5906 3159 5962 3168
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 5814 2680 5870 2689
rect 5814 2615 5816 2624
rect 5868 2615 5870 2624
rect 5816 2586 5868 2592
rect 6012 1494 6040 2926
rect 6104 2854 6132 4558
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6288 3738 6316 3878
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6472 3534 6500 3946
rect 6656 3777 6684 7908
rect 6748 7410 6776 8910
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6840 7546 6868 7890
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6748 6254 6776 7346
rect 6932 7342 6960 11154
rect 7024 8378 7052 11716
rect 7116 11608 7144 13126
rect 7300 11626 7328 13806
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7392 12850 7420 13262
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7484 12322 7512 14470
rect 7668 14396 7696 14554
rect 7576 14368 7696 14396
rect 7576 12442 7604 14368
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7668 13870 7696 14214
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7760 13326 7788 14855
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8220 14498 8248 15098
rect 8496 14890 8524 18119
rect 8484 14884 8536 14890
rect 8484 14826 8536 14832
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 8128 14470 8248 14498
rect 8036 14006 8064 14418
rect 8128 14414 8156 14470
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 8220 13190 8248 14350
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8312 13802 8340 13942
rect 8484 13932 8536 13938
rect 8484 13874 8536 13880
rect 8300 13796 8352 13802
rect 8300 13738 8352 13744
rect 8496 13394 8524 13874
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 7668 12782 7696 13126
rect 8312 12889 8340 13126
rect 8298 12880 8354 12889
rect 8298 12815 8354 12824
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7654 12472 7710 12481
rect 7564 12436 7616 12442
rect 7820 12464 8116 12484
rect 7654 12407 7656 12416
rect 7564 12378 7616 12384
rect 7708 12407 7710 12416
rect 7656 12378 7708 12384
rect 8404 12374 8432 12582
rect 8392 12368 8444 12374
rect 7196 11620 7248 11626
rect 7116 11580 7196 11608
rect 7196 11562 7248 11568
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7208 11150 7236 11562
rect 7300 11218 7328 11562
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7392 11150 7420 12310
rect 7484 12294 7604 12322
rect 8588 12322 8616 19110
rect 8680 18902 8708 19400
rect 8772 19174 8800 22222
rect 9048 20874 9076 22320
rect 9036 20868 9088 20874
rect 9036 20810 9088 20816
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8864 18970 8892 20198
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 8852 18964 8904 18970
rect 8852 18906 8904 18912
rect 8668 18896 8720 18902
rect 8668 18838 8720 18844
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8666 18320 8722 18329
rect 8666 18255 8722 18264
rect 8680 14498 8708 18255
rect 8772 17746 8800 18770
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 8956 16946 8984 19994
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9232 19174 9260 19790
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9232 18222 9260 19110
rect 9508 18358 9536 22320
rect 9772 20324 9824 20330
rect 9772 20266 9824 20272
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9692 18970 9720 19858
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9496 18352 9548 18358
rect 9496 18294 9548 18300
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 9784 17814 9812 20266
rect 9862 19272 9918 19281
rect 9862 19207 9918 19216
rect 9876 18766 9904 19207
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 8772 16918 8984 16946
rect 8772 16658 8800 16918
rect 8852 16788 8904 16794
rect 8852 16730 8904 16736
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 8760 16516 8812 16522
rect 8760 16458 8812 16464
rect 8772 16114 8800 16458
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8772 15609 8800 16050
rect 8758 15600 8814 15609
rect 8758 15535 8814 15544
rect 8680 14470 8800 14498
rect 8772 13734 8800 14470
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8772 12918 8800 13330
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8392 12310 8444 12316
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7484 11558 7512 12174
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7392 10606 7420 10950
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7300 9722 7328 10406
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 7116 9217 7144 9590
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7102 9208 7158 9217
rect 7102 9143 7158 9152
rect 7024 8362 7144 8378
rect 7024 8356 7156 8362
rect 7024 8350 7104 8356
rect 7104 8298 7156 8304
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 7208 6730 7236 9318
rect 7300 8090 7328 9318
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7392 8945 7420 9114
rect 7484 8974 7512 11494
rect 7576 9738 7604 12294
rect 8496 12294 8616 12322
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7668 11082 7696 11290
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7668 9926 7696 10542
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7576 9710 7696 9738
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7472 8968 7524 8974
rect 7378 8936 7434 8945
rect 7472 8910 7524 8916
rect 7378 8871 7434 8880
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 6748 5642 6776 6190
rect 7116 5710 7144 6190
rect 7104 5704 7156 5710
rect 7024 5664 7104 5692
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6748 4622 6776 5578
rect 6920 5568 6972 5574
rect 7024 5556 7052 5664
rect 7104 5646 7156 5652
rect 6972 5528 7052 5556
rect 6920 5510 6972 5516
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6932 4282 6960 4626
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 6642 3768 6698 3777
rect 6642 3703 6698 3712
rect 6460 3528 6512 3534
rect 6182 3496 6238 3505
rect 6460 3470 6512 3476
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6182 3431 6238 3440
rect 6092 2848 6144 2854
rect 6092 2790 6144 2796
rect 6000 1488 6052 1494
rect 6000 1430 6052 1436
rect 6104 1426 6132 2790
rect 6092 1420 6144 1426
rect 6092 1362 6144 1368
rect 6196 480 6224 3431
rect 6564 3058 6592 3470
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6656 2961 6684 3703
rect 7024 3534 7052 5528
rect 7392 5370 7420 8871
rect 7484 8362 7512 8910
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7484 7410 7512 8298
rect 7576 8022 7604 9386
rect 7668 9042 7696 9710
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7668 8022 7696 8774
rect 7564 8016 7616 8022
rect 7564 7958 7616 7964
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7576 4622 7604 7958
rect 7760 7954 7788 12038
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7944 11665 7972 11698
rect 7930 11656 7986 11665
rect 7930 11591 7986 11600
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8128 10606 8156 11086
rect 8116 10600 8168 10606
rect 8168 10560 8248 10588
rect 8116 10542 8168 10548
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 8220 10266 8248 10560
rect 8496 10470 8524 12294
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8588 11354 8616 12174
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8680 11354 8708 11630
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8666 11248 8722 11257
rect 8576 11212 8628 11218
rect 8666 11183 8722 11192
rect 8576 11154 8628 11160
rect 8588 10606 8616 11154
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8220 9586 8248 10202
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8312 9466 8340 9658
rect 8220 9438 8340 9466
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7852 8838 7880 8978
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8220 7002 8248 9438
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8312 9178 8340 9318
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8496 8974 8524 10066
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8404 8809 8432 8910
rect 8390 8800 8446 8809
rect 8390 8735 8446 8744
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8312 7886 8340 8230
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8312 6798 8340 7822
rect 8404 7002 8432 7822
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8496 6866 8524 7414
rect 8588 7274 8616 8230
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8390 5536 8446 5545
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7286 4448 7342 4457
rect 7286 4383 7342 4392
rect 7300 4078 7328 4383
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7470 4040 7526 4049
rect 7470 3975 7526 3984
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7116 3670 7144 3878
rect 7104 3664 7156 3670
rect 7104 3606 7156 3612
rect 7194 3632 7250 3641
rect 7194 3567 7250 3576
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 7024 3126 7052 3470
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 6642 2952 6698 2961
rect 6642 2887 6698 2896
rect 7208 1850 7236 3567
rect 7286 2816 7342 2825
rect 7286 2751 7342 2760
rect 7300 2553 7328 2751
rect 7286 2544 7342 2553
rect 7286 2479 7342 2488
rect 7116 1822 7236 1850
rect 6644 1760 6696 1766
rect 6644 1702 6696 1708
rect 6656 480 6684 1702
rect 7116 480 7144 1822
rect 7484 1306 7512 3975
rect 7564 2440 7616 2446
rect 7668 2428 7696 4762
rect 7746 4720 7802 4729
rect 7746 4655 7802 4664
rect 7760 3738 7788 4655
rect 8220 4622 8248 5510
rect 8390 5471 8446 5480
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8220 4214 8248 4558
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8312 4146 8340 4558
rect 8404 4486 8432 5471
rect 8482 4856 8538 4865
rect 8482 4791 8538 4800
rect 8496 4554 8524 4791
rect 8680 4690 8708 11183
rect 8772 9738 8800 11834
rect 8864 11393 8892 16730
rect 8956 14906 8984 16918
rect 9034 16688 9090 16697
rect 9034 16623 9036 16632
rect 9088 16623 9090 16632
rect 9036 16594 9088 16600
rect 9692 16538 9720 17206
rect 9784 17066 9812 17546
rect 9772 17060 9824 17066
rect 9772 17002 9824 17008
rect 9600 16510 9720 16538
rect 9784 16522 9812 17002
rect 9968 16794 9996 22320
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 10060 18834 10088 19790
rect 10140 19236 10192 19242
rect 10140 19178 10192 19184
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 10152 18766 10180 19178
rect 10244 19009 10272 19178
rect 10230 19000 10286 19009
rect 10230 18935 10286 18944
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10324 18692 10376 18698
rect 10324 18634 10376 18640
rect 10336 18426 10364 18634
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10428 18306 10456 22320
rect 10508 19916 10560 19922
rect 10508 19858 10560 19864
rect 10520 18426 10548 19858
rect 10888 18970 10916 22320
rect 11348 19802 11376 22320
rect 11808 20074 11836 22320
rect 11808 20046 11928 20074
rect 11796 19984 11848 19990
rect 11796 19926 11848 19932
rect 11164 19774 11376 19802
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 11072 18970 11100 19246
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 10692 18828 10744 18834
rect 10692 18770 10744 18776
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10428 18278 10548 18306
rect 10416 18216 10468 18222
rect 10416 18158 10468 18164
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10152 17202 10180 17614
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 9772 16516 9824 16522
rect 9600 16266 9628 16510
rect 9772 16458 9824 16464
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9508 16238 9628 16266
rect 9232 16114 9260 16186
rect 9508 16114 9536 16238
rect 9692 16130 9720 16390
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9600 16102 9720 16130
rect 9772 16176 9824 16182
rect 9772 16118 9824 16124
rect 9600 16046 9628 16102
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 9048 15473 9076 15506
rect 9034 15464 9090 15473
rect 9034 15399 9090 15408
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 9140 15026 9168 15302
rect 9416 15026 9444 15642
rect 9496 15156 9548 15162
rect 9548 15116 9628 15144
rect 9496 15098 9548 15104
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 9496 14952 9548 14958
rect 8956 14878 9168 14906
rect 9496 14894 9548 14900
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 8956 14618 8984 14758
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 9048 14074 9076 14758
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 8956 12782 8984 14010
rect 9140 13954 9168 14878
rect 9508 14550 9536 14894
rect 9496 14544 9548 14550
rect 9496 14486 9548 14492
rect 9600 14414 9628 15116
rect 9312 14408 9364 14414
rect 9588 14408 9640 14414
rect 9312 14350 9364 14356
rect 9494 14376 9550 14385
rect 9048 13926 9168 13954
rect 9324 13938 9352 14350
rect 9588 14350 9640 14356
rect 9494 14311 9550 14320
rect 9508 14278 9536 14311
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9312 13932 9364 13938
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 8956 11898 8984 12242
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 8850 11384 8906 11393
rect 8850 11319 8906 11328
rect 9048 11218 9076 13926
rect 9312 13874 9364 13880
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9140 13002 9168 13670
rect 9232 13530 9260 13670
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9140 12974 9260 13002
rect 9128 12912 9180 12918
rect 9128 12854 9180 12860
rect 9140 12238 9168 12854
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9232 11898 9260 12974
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9324 11762 9352 13874
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9416 12442 9444 12582
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9508 12322 9536 14214
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9600 12850 9628 13398
rect 9692 13326 9720 13670
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9416 12294 9536 12322
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 8956 10452 8984 11154
rect 8956 10424 9076 10452
rect 8772 9710 8984 9738
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8772 9042 8800 9522
rect 8956 9450 8984 9710
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8944 9444 8996 9450
rect 8944 9386 8996 9392
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8298 3904 8354 3913
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7760 3602 7788 3674
rect 7748 3596 7800 3602
rect 7800 3556 7880 3584
rect 7748 3538 7800 3544
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7760 3058 7788 3334
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7852 2904 7880 3556
rect 7760 2876 7880 2904
rect 7760 2446 7788 2876
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8220 2496 8248 3878
rect 8298 3839 8354 3848
rect 8312 3369 8340 3839
rect 8404 3738 8432 4082
rect 8588 4078 8616 4422
rect 8680 4185 8708 4626
rect 8666 4176 8722 4185
rect 8666 4111 8722 4120
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8298 3360 8354 3369
rect 8298 3295 8354 3304
rect 8404 2990 8432 3674
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8312 2582 8340 2790
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8128 2468 8248 2496
rect 7616 2400 7696 2428
rect 7748 2440 7800 2446
rect 7564 2382 7616 2388
rect 7748 2382 7800 2388
rect 7576 1630 7604 2382
rect 8128 2378 8156 2468
rect 8116 2372 8168 2378
rect 8116 2314 8168 2320
rect 8116 1692 8168 1698
rect 8116 1634 8168 1640
rect 7564 1624 7616 1630
rect 7564 1566 7616 1572
rect 7484 1278 7604 1306
rect 7576 480 7604 1278
rect 8128 480 8156 1634
rect 8588 480 8616 3674
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8680 2650 8708 2790
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8772 1698 8800 8978
rect 8864 2428 8892 9386
rect 9048 7206 9076 10424
rect 9232 10169 9260 11494
rect 9324 11150 9352 11698
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9218 10160 9274 10169
rect 9218 10095 9274 10104
rect 9126 8800 9182 8809
rect 9126 8735 9182 8744
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9048 6254 9076 7142
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8956 5778 8984 6054
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 8956 5234 8984 5714
rect 9048 5681 9076 5714
rect 9034 5672 9090 5681
rect 9034 5607 9090 5616
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8942 4448 8998 4457
rect 8942 4383 8998 4392
rect 8956 4146 8984 4383
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9140 3738 9168 8735
rect 9232 7342 9260 10095
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9220 6928 9272 6934
rect 9220 6870 9272 6876
rect 9232 4729 9260 6870
rect 9218 4720 9274 4729
rect 9218 4655 9274 4664
rect 9312 4684 9364 4690
rect 9232 4622 9260 4655
rect 9312 4626 9364 4632
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 9048 2922 9076 3538
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 8864 2400 9076 2428
rect 8760 1692 8812 1698
rect 8760 1634 8812 1640
rect 9048 480 9076 2400
rect 9324 1698 9352 4626
rect 9416 3618 9444 12294
rect 9600 11937 9628 12582
rect 9586 11928 9642 11937
rect 9586 11863 9642 11872
rect 9586 11792 9642 11801
rect 9586 11727 9642 11736
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9508 3738 9536 11154
rect 9600 11150 9628 11727
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9692 10606 9720 11630
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 5545 9628 10406
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 9926 9720 9998
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 8838 9720 9862
rect 9784 9761 9812 16118
rect 10060 15978 10088 16730
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 10152 14958 10180 17138
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10244 16726 10272 17070
rect 10232 16720 10284 16726
rect 10232 16662 10284 16668
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 10336 16114 10364 16526
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 10152 13462 10180 13738
rect 10140 13456 10192 13462
rect 10140 13398 10192 13404
rect 9862 12336 9918 12345
rect 9862 12271 9918 12280
rect 9876 12170 9904 12271
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 9770 9752 9826 9761
rect 9770 9687 9826 9696
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9784 9353 9812 9590
rect 9968 9586 9996 12106
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 9864 9376 9916 9382
rect 9770 9344 9826 9353
rect 9864 9318 9916 9324
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9770 9279 9826 9288
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9692 8430 9720 8774
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9692 7886 9720 8366
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9692 6798 9720 7822
rect 9784 6866 9812 8774
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9692 6100 9720 6734
rect 9772 6112 9824 6118
rect 9692 6072 9772 6100
rect 9772 6054 9824 6060
rect 9678 5944 9734 5953
rect 9678 5879 9734 5888
rect 9692 5846 9720 5879
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9680 5568 9732 5574
rect 9586 5536 9642 5545
rect 9680 5510 9732 5516
rect 9586 5471 9642 5480
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9600 4486 9628 5170
rect 9692 5166 9720 5510
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9784 5012 9812 6054
rect 9692 4984 9812 5012
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9692 3777 9720 4984
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9784 4078 9812 4694
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9772 3936 9824 3942
rect 9876 3924 9904 9318
rect 9968 8265 9996 9318
rect 10060 8634 10088 9454
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10152 8906 10180 9318
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 9954 8256 10010 8265
rect 9954 8191 10010 8200
rect 10060 8022 10088 8570
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10046 7304 10102 7313
rect 10046 7239 10048 7248
rect 10100 7239 10102 7248
rect 10048 7210 10100 7216
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 9954 6896 10010 6905
rect 9954 6831 10010 6840
rect 9968 6662 9996 6831
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 10060 6254 10088 6938
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 10060 5574 10088 5782
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10060 4758 10088 4966
rect 10152 4826 10180 4966
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 9968 4457 9996 4558
rect 9954 4448 10010 4457
rect 9954 4383 10010 4392
rect 9956 3936 10008 3942
rect 9876 3896 9956 3924
rect 9772 3878 9824 3884
rect 9956 3878 10008 3884
rect 9678 3768 9734 3777
rect 9496 3732 9548 3738
rect 9678 3703 9734 3712
rect 9496 3674 9548 3680
rect 9416 3590 9628 3618
rect 9600 2666 9628 3590
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9692 3194 9720 3538
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9508 2638 9628 2666
rect 9312 1692 9364 1698
rect 9312 1634 9364 1640
rect 9324 1562 9352 1634
rect 9312 1556 9364 1562
rect 9312 1498 9364 1504
rect 9508 480 9536 2638
rect 9692 2446 9720 3130
rect 9784 2582 9812 3878
rect 9862 3768 9918 3777
rect 9862 3703 9918 3712
rect 9956 3732 10008 3738
rect 9876 3534 9904 3703
rect 9956 3674 10008 3680
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 9876 2990 9904 3062
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9968 480 9996 3674
rect 10060 3126 10088 4558
rect 10244 4264 10272 15982
rect 10428 12918 10456 18158
rect 10520 16046 10548 18278
rect 10612 17678 10640 18702
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10704 16182 10732 18770
rect 11164 18170 11192 19774
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 11610 19000 11666 19009
rect 11610 18935 11666 18944
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11624 18290 11652 18935
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11164 18142 11652 18170
rect 11716 18154 11744 19246
rect 11808 18290 11836 19926
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10888 16794 10916 17478
rect 11072 17066 11100 17750
rect 11164 17202 11192 18022
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11624 17252 11652 18142
rect 11704 18148 11756 18154
rect 11704 18090 11756 18096
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11532 17224 11652 17252
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 11072 16590 11100 17002
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10508 15088 10560 15094
rect 10508 15030 10560 15036
rect 10520 14498 10548 15030
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10612 14822 10640 14894
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10612 14618 10640 14758
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10520 14470 10640 14498
rect 10612 14414 10640 14470
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10520 13938 10548 14350
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10428 11694 10456 12718
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10612 11830 10640 12174
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 10612 11558 10640 11766
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10152 4236 10272 4264
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 10152 2990 10180 4236
rect 10232 4004 10284 4010
rect 10232 3946 10284 3952
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 10152 2553 10180 2790
rect 10244 2650 10272 3946
rect 10336 3777 10364 11154
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10520 9217 10548 9318
rect 10506 9208 10562 9217
rect 10506 9143 10562 9152
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10428 8566 10456 8910
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 10428 6390 10456 8502
rect 10520 7206 10548 8842
rect 10612 7857 10640 8978
rect 10598 7848 10654 7857
rect 10598 7783 10654 7792
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10506 6760 10562 6769
rect 10506 6695 10562 6704
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10428 5710 10456 6054
rect 10520 5846 10548 6695
rect 10508 5840 10560 5846
rect 10508 5782 10560 5788
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10506 5672 10562 5681
rect 10506 5607 10562 5616
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10322 3768 10378 3777
rect 10322 3703 10378 3712
rect 10428 3670 10456 3878
rect 10416 3664 10468 3670
rect 10520 3641 10548 5607
rect 10612 3738 10640 7686
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10416 3606 10468 3612
rect 10506 3632 10562 3641
rect 10506 3567 10562 3576
rect 10704 3210 10732 15574
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11072 14890 11100 15302
rect 11060 14884 11112 14890
rect 11060 14826 11112 14832
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10796 14074 10824 14418
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10888 13734 10916 14554
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 11072 13977 11100 14486
rect 11058 13968 11114 13977
rect 11058 13903 11114 13912
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 13326 10916 13670
rect 10876 13320 10928 13326
rect 10796 13280 10876 13308
rect 10796 12782 10824 13280
rect 10876 13262 10928 13268
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10888 10713 10916 12922
rect 10874 10704 10930 10713
rect 10874 10639 10930 10648
rect 10980 10266 11008 13806
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 11072 12442 11100 13330
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11072 10810 11100 11562
rect 11164 11082 11192 16594
rect 11440 16538 11468 16934
rect 11532 16726 11560 17224
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11624 16794 11652 16934
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11520 16720 11572 16726
rect 11518 16688 11520 16697
rect 11572 16688 11574 16697
rect 11518 16623 11574 16632
rect 11440 16510 11652 16538
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11348 15706 11376 15982
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11518 13968 11574 13977
rect 11518 13903 11520 13912
rect 11572 13903 11574 13912
rect 11520 13874 11572 13880
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11256 13258 11284 13670
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 11532 13172 11560 13874
rect 11624 13326 11652 16510
rect 11716 16114 11744 17818
rect 11900 17762 11928 20046
rect 12164 19984 12216 19990
rect 12164 19926 12216 19932
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 11992 17882 12020 18770
rect 12084 18630 12112 19110
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 11900 17734 12020 17762
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11900 16794 11928 17614
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11704 15972 11756 15978
rect 11704 15914 11756 15920
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11612 13184 11664 13190
rect 11532 13144 11612 13172
rect 11612 13126 11664 13132
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11716 12424 11744 15914
rect 11624 12396 11744 12424
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11426 11384 11482 11393
rect 11426 11319 11482 11328
rect 11440 11286 11468 11319
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11336 11144 11388 11150
rect 11334 11112 11336 11121
rect 11388 11112 11390 11121
rect 11152 11076 11204 11082
rect 11532 11098 11560 11562
rect 11624 11234 11652 12396
rect 11808 12374 11836 16594
rect 11992 15910 12020 17734
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11888 15632 11940 15638
rect 12084 15620 12112 18022
rect 12176 15978 12204 19926
rect 12268 16794 12296 22320
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12360 18086 12388 19858
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12164 15972 12216 15978
rect 12164 15914 12216 15920
rect 11940 15592 12112 15620
rect 11888 15574 11940 15580
rect 12084 15026 12112 15592
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11992 14414 12020 14758
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 12268 13716 12296 16730
rect 12360 16658 12388 17546
rect 12452 17270 12480 18158
rect 12440 17264 12492 17270
rect 12440 17206 12492 17212
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12440 16040 12492 16046
rect 12544 16028 12572 19246
rect 12636 18290 12664 19858
rect 12728 19394 12756 22320
rect 13188 20058 13216 22320
rect 13648 20058 13676 22320
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 12728 19366 12848 19394
rect 12716 19236 12768 19242
rect 12716 19178 12768 19184
rect 12728 18698 12756 19178
rect 12820 18970 12848 19366
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12992 18896 13044 18902
rect 12992 18838 13044 18844
rect 12716 18692 12768 18698
rect 12716 18634 12768 18640
rect 13004 18630 13032 18838
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 12820 18358 12848 18566
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13188 16726 13216 17070
rect 13176 16720 13228 16726
rect 13082 16688 13138 16697
rect 12624 16652 12676 16658
rect 13176 16662 13228 16668
rect 13082 16623 13138 16632
rect 12624 16594 12676 16600
rect 12492 16000 12572 16028
rect 12440 15982 12492 15988
rect 12452 15570 12480 15982
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12452 14346 12480 15506
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12544 14074 12572 15642
rect 12636 15162 12664 16594
rect 12716 15972 12768 15978
rect 12716 15914 12768 15920
rect 12728 15638 12756 15914
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12268 13688 12388 13716
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11716 11354 11744 12242
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11624 11206 11744 11234
rect 11532 11070 11652 11098
rect 11334 11047 11390 11056
rect 11152 11018 11204 11024
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10980 9178 11008 10202
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10888 9058 10916 9114
rect 10784 9036 10836 9042
rect 10888 9030 11008 9058
rect 10784 8978 10836 8984
rect 10796 8838 10824 8978
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10980 8650 11008 9030
rect 11072 8809 11100 10542
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11164 9722 11192 10202
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11348 9081 11376 9318
rect 11532 9217 11560 9522
rect 11518 9208 11574 9217
rect 11518 9143 11574 9152
rect 11334 9072 11390 9081
rect 11334 9007 11390 9016
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11058 8800 11114 8809
rect 11058 8735 11114 8744
rect 10980 8622 11100 8650
rect 11072 8401 11100 8622
rect 11058 8392 11114 8401
rect 11164 8362 11192 8910
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11624 8480 11652 11070
rect 11716 10538 11744 11206
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11532 8452 11652 8480
rect 11058 8327 11114 8336
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10796 7546 10824 8026
rect 11532 7993 11560 8452
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11518 7984 11574 7993
rect 11518 7919 11574 7928
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10888 6934 10916 7686
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11520 7472 11572 7478
rect 11520 7414 11572 7420
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10796 6458 10824 6734
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10796 5778 10824 6054
rect 10888 5846 10916 6870
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10888 4622 10916 5646
rect 10980 5273 11008 7346
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 10966 5264 11022 5273
rect 10966 5199 10968 5208
rect 11020 5199 11022 5208
rect 10968 5170 11020 5176
rect 10966 4720 11022 4729
rect 10966 4655 10968 4664
rect 11020 4655 11022 4664
rect 10968 4626 11020 4632
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 11072 4554 11100 6666
rect 11164 6458 11192 7278
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11256 6730 11284 7142
rect 11532 7002 11560 7414
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11624 6458 11652 8298
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11426 6352 11482 6361
rect 11152 6316 11204 6322
rect 11624 6322 11652 6394
rect 11426 6287 11482 6296
rect 11612 6316 11664 6322
rect 11152 6258 11204 6264
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 10966 4448 11022 4457
rect 10966 4383 11022 4392
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 10428 3182 10732 3210
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10138 2544 10194 2553
rect 10138 2479 10194 2488
rect 10336 2417 10364 2994
rect 10322 2408 10378 2417
rect 10322 2343 10378 2352
rect 10428 480 10456 3182
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10612 2514 10640 2994
rect 10796 2514 10824 4150
rect 10980 4146 11008 4383
rect 11058 4312 11114 4321
rect 11058 4247 11114 4256
rect 11072 4214 11100 4247
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10980 4010 11008 4082
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 11164 3942 11192 6258
rect 11440 6186 11468 6287
rect 11612 6258 11664 6264
rect 11428 6180 11480 6186
rect 11428 6122 11480 6128
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11244 5772 11296 5778
rect 11348 5760 11376 6054
rect 11296 5732 11376 5760
rect 11244 5714 11296 5720
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11336 4004 11388 4010
rect 11256 3964 11336 3992
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11256 3754 11284 3964
rect 11336 3946 11388 3952
rect 10980 3738 11284 3754
rect 10968 3732 11284 3738
rect 11020 3726 11284 3732
rect 10968 3674 11020 3680
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 11518 3632 11574 3641
rect 10966 3224 11022 3233
rect 10966 3159 11022 3168
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10888 2650 10916 2926
rect 10980 2825 11008 3159
rect 10966 2816 11022 2825
rect 10966 2751 11022 2760
rect 11072 2650 11100 3606
rect 11164 3058 11192 3606
rect 11518 3567 11574 3576
rect 11532 3534 11560 3567
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11336 3052 11388 3058
rect 11336 2994 11388 3000
rect 11348 2650 11376 2994
rect 11624 2990 11652 5034
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10874 2272 10930 2281
rect 10874 2207 10930 2216
rect 10888 480 10916 2207
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11624 1834 11652 2518
rect 11716 2394 11744 10474
rect 11808 6746 11836 12310
rect 11900 12306 11928 12650
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11900 11898 11928 12242
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11900 11082 11928 11834
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11900 10130 11928 10202
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11900 9761 11928 10066
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11886 9752 11942 9761
rect 11886 9687 11942 9696
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 11900 8090 11928 9590
rect 11992 9586 12020 9862
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 12084 9364 12112 13194
rect 12176 12986 12204 13330
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12176 12238 12204 12922
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12176 11257 12204 11630
rect 12254 11384 12310 11393
rect 12254 11319 12256 11328
rect 12308 11319 12310 11328
rect 12256 11290 12308 11296
rect 12162 11248 12218 11257
rect 12162 11183 12218 11192
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12162 9752 12218 9761
rect 12162 9687 12218 9696
rect 12176 9518 12204 9687
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 11978 9344 12034 9353
rect 12084 9336 12204 9364
rect 11978 9279 12034 9288
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11992 7002 12020 9279
rect 12176 9178 12204 9336
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12084 7410 12112 8978
rect 12268 8129 12296 11086
rect 12254 8120 12310 8129
rect 12254 8055 12310 8064
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 12072 6792 12124 6798
rect 11808 6718 11928 6746
rect 12072 6734 12124 6740
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11808 5234 11836 6598
rect 11900 5658 11928 6718
rect 12084 5778 12112 6734
rect 12176 6118 12204 7890
rect 12256 7268 12308 7274
rect 12256 7210 12308 7216
rect 12268 6730 12296 7210
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 11900 5630 12204 5658
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11900 4622 11928 5170
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11808 4321 11836 4490
rect 11794 4312 11850 4321
rect 11794 4247 11850 4256
rect 11794 3768 11850 3777
rect 11794 3703 11850 3712
rect 11808 3233 11836 3703
rect 11794 3224 11850 3233
rect 11794 3159 11850 3168
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11808 2514 11836 3062
rect 11992 2514 12020 5510
rect 12070 5400 12126 5409
rect 12070 5335 12126 5344
rect 12084 5030 12112 5335
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 12070 4856 12126 4865
rect 12070 4791 12126 4800
rect 12084 4185 12112 4791
rect 12070 4176 12126 4185
rect 12070 4111 12126 4120
rect 12176 3652 12204 5630
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12268 4690 12296 5238
rect 12360 5137 12388 13688
rect 12636 12986 12664 14486
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12820 13938 12848 14214
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12912 13870 12940 14214
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12544 12442 12572 12582
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12440 12368 12492 12374
rect 12440 12310 12492 12316
rect 12452 11257 12480 12310
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12438 11248 12494 11257
rect 12438 11183 12494 11192
rect 12440 10192 12492 10198
rect 12438 10160 12440 10169
rect 12492 10160 12494 10169
rect 12438 10095 12494 10104
rect 12544 9586 12572 11562
rect 12636 10470 12664 12378
rect 12912 12102 12940 13670
rect 13004 12986 13032 14418
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 13004 12442 13032 12718
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12900 11824 12952 11830
rect 12900 11766 12952 11772
rect 12912 11286 12940 11766
rect 13004 11762 13032 12174
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 12728 10606 12756 11222
rect 12820 10810 12848 11222
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12990 11112 13046 11121
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12440 8968 12492 8974
rect 12636 8922 12664 10406
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12728 9178 12756 9318
rect 12912 9217 12940 11086
rect 12990 11047 13046 11056
rect 12898 9208 12954 9217
rect 12716 9172 12768 9178
rect 13004 9178 13032 11047
rect 12898 9143 12954 9152
rect 12992 9172 13044 9178
rect 12716 9114 12768 9120
rect 12992 9114 13044 9120
rect 12440 8910 12492 8916
rect 12452 8362 12480 8910
rect 12544 8894 12664 8922
rect 12900 8900 12952 8906
rect 12544 8430 12572 8894
rect 12900 8842 12952 8848
rect 12992 8900 13044 8906
rect 12992 8842 13044 8848
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12636 8430 12664 8774
rect 12912 8498 12940 8842
rect 13004 8634 13032 8842
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12544 7002 12572 7142
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12636 6934 12664 8026
rect 12728 8022 12756 8434
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12912 6780 12940 8298
rect 13004 8022 13032 8434
rect 12992 8016 13044 8022
rect 12992 7958 13044 7964
rect 13004 7410 13032 7958
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12992 6792 13044 6798
rect 12912 6752 12992 6780
rect 12992 6734 13044 6740
rect 13096 6746 13124 16623
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 13188 13530 13216 14826
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13280 12374 13308 18770
rect 13372 18290 13400 19858
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13372 13410 13400 15846
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13464 13938 13492 14418
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13464 13530 13492 13874
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13372 13382 13492 13410
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13188 11150 13216 12038
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13280 10169 13308 11086
rect 13372 11082 13400 11562
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13266 10160 13322 10169
rect 13266 10095 13322 10104
rect 13280 8974 13308 10095
rect 13360 9104 13412 9110
rect 13360 9046 13412 9052
rect 13268 8968 13320 8974
rect 13174 8936 13230 8945
rect 13268 8910 13320 8916
rect 13174 8871 13230 8880
rect 13188 8498 13216 8871
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13280 7546 13308 8910
rect 13372 8265 13400 9046
rect 13358 8256 13414 8265
rect 13358 8191 13414 8200
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13372 7750 13400 7890
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13372 7410 13400 7686
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13464 7002 13492 13382
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13556 12306 13584 12922
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13648 12186 13676 19178
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13832 19009 13860 19110
rect 13818 19000 13874 19009
rect 13818 18935 13874 18944
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13740 13734 13768 18362
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13556 12170 13676 12186
rect 13544 12164 13676 12170
rect 13596 12158 13676 12164
rect 13544 12106 13596 12112
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13634 10704 13690 10713
rect 13740 10674 13768 11630
rect 13832 11354 13860 18770
rect 14108 17338 14136 22320
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 14016 15638 14044 15982
rect 14004 15632 14056 15638
rect 14004 15574 14056 15580
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 13912 14816 13964 14822
rect 14016 14804 14044 14962
rect 13964 14776 14044 14804
rect 13912 14758 13964 14764
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13924 13870 13952 14350
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13924 12374 13952 12582
rect 14016 12458 14044 14776
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14108 13530 14136 14758
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14108 12594 14136 13194
rect 14200 12714 14228 19246
rect 14292 18902 14320 19246
rect 14568 19174 14596 22320
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 15028 19174 15056 22320
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 14280 18896 14332 18902
rect 14280 18838 14332 18844
rect 15108 18624 15160 18630
rect 15108 18566 15160 18572
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 14476 17202 14504 17682
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14384 15706 14412 15846
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14292 14346 14320 15506
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 14292 14074 14320 14282
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14384 13530 14412 13670
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14108 12566 14228 12594
rect 14016 12430 14136 12458
rect 13912 12368 13964 12374
rect 13912 12310 13964 12316
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13924 11150 13952 12310
rect 14016 11218 14044 12310
rect 14108 11626 14136 12430
rect 14200 11694 14228 12566
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14096 11620 14148 11626
rect 14096 11562 14148 11568
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13832 10674 13860 11086
rect 13634 10639 13690 10648
rect 13728 10668 13780 10674
rect 13648 10470 13676 10639
rect 13728 10610 13780 10616
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13556 8022 13584 10066
rect 13740 9586 13768 10610
rect 14200 10554 14228 11630
rect 14292 11354 14320 13126
rect 14384 12782 14412 13262
rect 14476 13258 14504 17138
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14568 14618 14596 14758
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 15028 13938 15056 14894
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 15120 13818 15148 18566
rect 15212 14346 15240 19246
rect 15580 19174 15608 22320
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15384 18828 15436 18834
rect 15384 18770 15436 18776
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 15304 14414 15332 14826
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15304 14006 15332 14214
rect 15292 14000 15344 14006
rect 15198 13968 15254 13977
rect 15292 13942 15344 13948
rect 15198 13903 15200 13912
rect 15252 13903 15254 13912
rect 15200 13874 15252 13880
rect 14648 13796 14700 13802
rect 14568 13756 14648 13784
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14384 11898 14412 12718
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14568 11676 14596 13756
rect 14648 13738 14700 13744
rect 15028 13790 15148 13818
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 14936 11694 14964 12174
rect 14476 11648 14596 11676
rect 14924 11688 14976 11694
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 13832 10526 14228 10554
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13728 9376 13780 9382
rect 13726 9344 13728 9353
rect 13780 9344 13782 9353
rect 13726 9279 13782 9288
rect 13832 8786 13860 10526
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 13648 8758 13860 8786
rect 13544 8016 13596 8022
rect 13544 7958 13596 7964
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13360 6792 13412 6798
rect 13096 6718 13308 6746
rect 13360 6734 13412 6740
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 12716 6180 12768 6186
rect 12716 6122 12768 6128
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12452 5846 12480 6054
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12452 5302 12480 5782
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12452 5166 12480 5238
rect 12544 5166 12572 5510
rect 12636 5370 12664 6054
rect 12728 5370 12756 6122
rect 13188 5930 13216 6598
rect 12912 5902 13216 5930
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12440 5160 12492 5166
rect 12346 5128 12402 5137
rect 12440 5102 12492 5108
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12346 5063 12402 5072
rect 12440 5024 12492 5030
rect 12438 4992 12440 5001
rect 12532 5024 12584 5030
rect 12492 4992 12494 5001
rect 12532 4966 12584 4972
rect 12438 4927 12494 4936
rect 12438 4856 12494 4865
rect 12544 4826 12572 4966
rect 12438 4791 12494 4800
rect 12532 4820 12584 4826
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12268 3777 12296 4626
rect 12452 4214 12480 4791
rect 12532 4762 12584 4768
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12636 4690 12664 4762
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 12532 4480 12584 4486
rect 12584 4440 12664 4468
rect 12532 4422 12584 4428
rect 12348 4208 12400 4214
rect 12348 4150 12400 4156
rect 12440 4208 12492 4214
rect 12440 4150 12492 4156
rect 12360 4049 12388 4150
rect 12346 4040 12402 4049
rect 12346 3975 12402 3984
rect 12636 3942 12664 4440
rect 12728 4214 12756 5306
rect 12912 5001 12940 5902
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 12992 5092 13044 5098
rect 12992 5034 13044 5040
rect 12898 4992 12954 5001
rect 12898 4927 12954 4936
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 12912 4146 12940 4422
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 13004 3942 13032 5034
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 12348 3936 12400 3942
rect 12624 3936 12676 3942
rect 12400 3896 12572 3924
rect 12348 3878 12400 3884
rect 12254 3768 12310 3777
rect 12254 3703 12310 3712
rect 12176 3624 12296 3652
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 12084 2553 12112 2926
rect 12070 2544 12126 2553
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11980 2508 12032 2514
rect 12070 2479 12126 2488
rect 11980 2450 12032 2456
rect 11716 2366 11836 2394
rect 11612 1828 11664 1834
rect 11612 1770 11664 1776
rect 11336 1420 11388 1426
rect 11336 1362 11388 1368
rect 11348 480 11376 1362
rect 11808 480 11836 2366
rect 12176 1630 12204 3334
rect 12164 1624 12216 1630
rect 12164 1566 12216 1572
rect 12268 480 12296 3624
rect 12440 3392 12492 3398
rect 12360 3340 12440 3346
rect 12360 3334 12492 3340
rect 12360 3318 12480 3334
rect 12360 1426 12388 3318
rect 12544 3058 12572 3896
rect 12624 3878 12676 3884
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 12714 3768 12770 3777
rect 12990 3768 13046 3777
rect 12714 3703 12770 3712
rect 12808 3732 12860 3738
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12636 3194 12664 3334
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 12636 2825 12664 2858
rect 12622 2816 12678 2825
rect 12622 2751 12678 2760
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 12636 1902 12664 2246
rect 12624 1896 12676 1902
rect 12624 1838 12676 1844
rect 12348 1420 12400 1426
rect 12348 1362 12400 1368
rect 12728 480 12756 3703
rect 13096 3738 13124 4626
rect 13188 4078 13216 5714
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 12990 3703 13046 3712
rect 13084 3732 13136 3738
rect 12808 3674 12860 3680
rect 12820 3194 12848 3674
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 13004 2961 13032 3703
rect 13084 3674 13136 3680
rect 13280 3670 13308 6718
rect 13372 6458 13400 6734
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13372 4214 13400 5646
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13450 5400 13506 5409
rect 13450 5335 13506 5344
rect 13464 5302 13492 5335
rect 13452 5296 13504 5302
rect 13452 5238 13504 5244
rect 13452 5092 13504 5098
rect 13452 5034 13504 5040
rect 13464 4729 13492 5034
rect 13450 4720 13506 4729
rect 13450 4655 13506 4664
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13372 3534 13400 3878
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 12990 2952 13046 2961
rect 12990 2887 13046 2896
rect 13004 2553 13032 2887
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 12990 2544 13046 2553
rect 12990 2479 13046 2488
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13188 1766 13216 2382
rect 13280 2106 13308 2790
rect 13464 2582 13492 3606
rect 13556 2802 13584 5510
rect 13648 5114 13676 8758
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13832 7342 13860 8570
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13924 6866 13952 10406
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14016 8090 14044 9318
rect 14108 8673 14136 9522
rect 14200 9450 14228 10406
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 14292 9178 14320 10406
rect 14384 10266 14412 11494
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14476 9568 14504 11648
rect 14924 11630 14976 11636
rect 15028 11642 15056 13790
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15304 12442 15332 13330
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15028 11614 15240 11642
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 14568 11286 14596 11494
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14568 9586 14596 11018
rect 14660 10606 14688 11086
rect 15028 10810 15056 11494
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14384 9540 14504 9568
rect 14556 9580 14608 9586
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14094 8664 14150 8673
rect 14200 8634 14228 8910
rect 14094 8599 14150 8608
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 14004 7268 14056 7274
rect 14004 7210 14056 7216
rect 14016 6905 14044 7210
rect 14002 6896 14058 6905
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13912 6860 13964 6866
rect 14002 6831 14058 6840
rect 13912 6802 13964 6808
rect 13832 6322 13860 6802
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13832 5352 13860 5714
rect 13912 5364 13964 5370
rect 13832 5324 13912 5352
rect 13832 5273 13860 5324
rect 13912 5306 13964 5312
rect 13818 5264 13874 5273
rect 14016 5250 14044 6734
rect 14108 5817 14136 8230
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14094 5808 14150 5817
rect 14094 5743 14150 5752
rect 14094 5672 14150 5681
rect 14094 5607 14150 5616
rect 13818 5199 13874 5208
rect 13924 5222 14044 5250
rect 13648 5086 13860 5114
rect 13832 3942 13860 5086
rect 13924 4826 13952 5222
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 13924 4729 13952 4762
rect 13910 4720 13966 4729
rect 13910 4655 13966 4664
rect 13910 4584 13966 4593
rect 14016 4554 14044 4966
rect 13910 4519 13966 4528
rect 14004 4548 14056 4554
rect 13924 4146 13952 4519
rect 14004 4490 14056 4496
rect 14108 4434 14136 5607
rect 14016 4406 14136 4434
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13726 3768 13782 3777
rect 13726 3703 13782 3712
rect 13740 3670 13768 3703
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13556 2774 13676 2802
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13268 2100 13320 2106
rect 13268 2042 13320 2048
rect 13176 1760 13228 1766
rect 13176 1702 13228 1708
rect 13372 1698 13400 2450
rect 13360 1692 13412 1698
rect 13360 1634 13412 1640
rect 13176 1624 13228 1630
rect 13176 1566 13228 1572
rect 13188 480 13216 1566
rect 13648 480 13676 2774
rect 13924 1970 13952 3946
rect 14016 3516 14044 4406
rect 14200 3720 14228 7142
rect 14292 6225 14320 9114
rect 14384 9042 14412 9540
rect 14556 9522 14608 9528
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 14462 9480 14518 9489
rect 14568 9466 14596 9522
rect 14568 9450 14688 9466
rect 14568 9444 14700 9450
rect 14568 9438 14648 9444
rect 14462 9415 14518 9424
rect 14476 9382 14504 9415
rect 14648 9386 14700 9392
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14372 9036 14424 9042
rect 14372 8978 14424 8984
rect 14568 7857 14596 9318
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 15028 8974 15056 9522
rect 15120 9518 15148 11494
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 15014 8528 15070 8537
rect 15014 8463 15016 8472
rect 15068 8463 15070 8472
rect 15016 8434 15068 8440
rect 15016 8356 15068 8362
rect 15016 8298 15068 8304
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14554 7848 14610 7857
rect 14554 7783 14610 7792
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14476 6769 14504 7142
rect 14462 6760 14518 6769
rect 14462 6695 14518 6704
rect 14464 6248 14516 6254
rect 14278 6216 14334 6225
rect 14464 6190 14516 6196
rect 14278 6151 14334 6160
rect 14476 5846 14504 6190
rect 14464 5840 14516 5846
rect 14464 5782 14516 5788
rect 14568 5370 14596 7686
rect 15028 7410 15056 8298
rect 15212 8294 15240 11614
rect 15396 9081 15424 18770
rect 15764 14550 15792 19246
rect 16040 19174 16068 22320
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16028 19168 16080 19174
rect 16028 19110 16080 19116
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 16212 14544 16264 14550
rect 16212 14486 16264 14492
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15856 13938 15884 14350
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15382 9072 15438 9081
rect 15382 9007 15438 9016
rect 15488 8956 15516 12378
rect 15396 8928 15516 8956
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 15028 5681 15056 7346
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15014 5672 15070 5681
rect 15014 5607 15070 5616
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 14752 5234 14780 5306
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14292 4865 14320 5102
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14278 4856 14334 4865
rect 14684 4848 14980 4868
rect 14278 4791 14334 4800
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14384 4486 14412 4762
rect 14646 4720 14702 4729
rect 14646 4655 14702 4664
rect 14660 4622 14688 4655
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14372 3936 14424 3942
rect 14370 3904 14372 3913
rect 14424 3904 14426 3913
rect 14370 3839 14426 3848
rect 14108 3692 14228 3720
rect 14278 3768 14334 3777
rect 14278 3703 14334 3712
rect 14372 3732 14424 3738
rect 14108 3641 14136 3692
rect 14094 3632 14150 3641
rect 14292 3602 14320 3703
rect 14372 3674 14424 3680
rect 14094 3567 14150 3576
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14016 3488 14136 3516
rect 14004 2984 14056 2990
rect 14002 2952 14004 2961
rect 14056 2952 14058 2961
rect 14002 2887 14058 2896
rect 13912 1964 13964 1970
rect 13912 1906 13964 1912
rect 14016 1222 14044 2887
rect 14108 2428 14136 3488
rect 14200 2650 14228 3538
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14188 2440 14240 2446
rect 14108 2400 14188 2428
rect 14188 2382 14240 2388
rect 14096 1964 14148 1970
rect 14096 1906 14148 1912
rect 14004 1216 14056 1222
rect 14004 1158 14056 1164
rect 14108 480 14136 1906
rect 14292 1358 14320 3538
rect 14384 3505 14412 3674
rect 14476 3534 14504 4558
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14660 4146 14688 4218
rect 14648 4140 14700 4146
rect 14568 4100 14648 4128
rect 14464 3528 14516 3534
rect 14370 3496 14426 3505
rect 14464 3470 14516 3476
rect 14568 3466 14596 4100
rect 14648 4082 14700 4088
rect 14646 4040 14702 4049
rect 14646 3975 14648 3984
rect 14700 3975 14702 3984
rect 14648 3946 14700 3952
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14370 3431 14426 3440
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 14372 3052 14424 3058
rect 14568 3040 14596 3402
rect 14424 3012 14596 3040
rect 14646 3088 14702 3097
rect 14646 3023 14648 3032
rect 14372 2994 14424 3000
rect 14700 3023 14702 3032
rect 14648 2994 14700 3000
rect 14372 2916 14424 2922
rect 14372 2858 14424 2864
rect 14384 2038 14412 2858
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14476 2650 14504 2790
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14372 2032 14424 2038
rect 14372 1974 14424 1980
rect 14556 1760 14608 1766
rect 14556 1702 14608 1708
rect 14280 1352 14332 1358
rect 14280 1294 14332 1300
rect 14568 480 14596 1702
rect 15028 480 15056 4966
rect 15108 4004 15160 4010
rect 15108 3946 15160 3952
rect 15120 2378 15148 3946
rect 15212 3942 15240 7142
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15304 5166 15332 6598
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15304 4826 15332 4966
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15198 3632 15254 3641
rect 15198 3567 15200 3576
rect 15252 3567 15254 3576
rect 15200 3538 15252 3544
rect 15396 2961 15424 8928
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15580 6186 15608 6598
rect 15568 6180 15620 6186
rect 15568 6122 15620 6128
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15488 5234 15516 5782
rect 15580 5574 15608 6122
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15474 5128 15530 5137
rect 15474 5063 15530 5072
rect 15488 2990 15516 5063
rect 15580 4622 15608 5510
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15672 4026 15700 13466
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15856 11626 15884 12174
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15750 8392 15806 8401
rect 15750 8327 15806 8336
rect 15764 5234 15792 8327
rect 15934 7304 15990 7313
rect 15934 7239 15936 7248
rect 15988 7239 15990 7248
rect 15936 7210 15988 7216
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15764 4826 15792 4966
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15571 3998 15700 4026
rect 15571 3942 15599 3998
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15580 3058 15608 3878
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15476 2984 15528 2990
rect 15382 2952 15438 2961
rect 15476 2926 15528 2932
rect 15382 2887 15438 2896
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15212 2417 15240 2790
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15198 2408 15254 2417
rect 15108 2372 15160 2378
rect 15198 2343 15254 2352
rect 15108 2314 15160 2320
rect 15488 2106 15516 2586
rect 15476 2100 15528 2106
rect 15476 2042 15528 2048
rect 15764 2020 15792 3878
rect 15856 2514 15884 6938
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15948 5778 15976 6054
rect 16028 5840 16080 5846
rect 16028 5782 16080 5788
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 16040 5370 16068 5782
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 16026 5128 16082 5137
rect 16026 5063 16082 5072
rect 16040 5030 16068 5063
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 15948 4214 15976 4558
rect 16040 4321 16068 4626
rect 16026 4312 16082 4321
rect 16026 4247 16082 4256
rect 15936 4208 15988 4214
rect 15936 4150 15988 4156
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15948 3670 15976 4014
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 16132 2854 16160 5170
rect 16224 4434 16252 14486
rect 16316 12442 16344 19246
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16408 10470 16436 19858
rect 16500 19174 16528 22320
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16868 18902 16896 19246
rect 16960 19174 16988 22320
rect 17420 20058 17448 22320
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17316 19236 17368 19242
rect 17316 19178 17368 19184
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16856 18896 16908 18902
rect 16856 18838 16908 18844
rect 17328 12850 17356 19178
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 17052 12345 17080 12718
rect 17038 12336 17094 12345
rect 17038 12271 17094 12280
rect 17512 10742 17540 19246
rect 17880 19174 17908 22320
rect 18340 19700 18368 22320
rect 18696 19712 18748 19718
rect 18340 19672 18552 19700
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18524 19174 18552 19672
rect 18696 19654 18748 19660
rect 18708 19242 18736 19654
rect 18696 19236 18748 19242
rect 18696 19178 18748 19184
rect 18800 19174 18828 22320
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18800 9625 18828 18770
rect 19168 14482 19196 19246
rect 19260 19174 19288 22320
rect 19340 19984 19392 19990
rect 19340 19926 19392 19932
rect 19352 19718 19380 19926
rect 19720 19854 19748 22320
rect 20180 19990 20208 22320
rect 20168 19984 20220 19990
rect 20168 19926 20220 19932
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19720 18902 19748 19246
rect 20640 19174 20668 22320
rect 20628 19168 20680 19174
rect 20628 19110 20680 19116
rect 19708 18896 19760 18902
rect 19708 18838 19760 18844
rect 21100 18834 21128 22320
rect 21560 19242 21588 22320
rect 21548 19236 21600 19242
rect 21548 19178 21600 19184
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 19352 17882 19380 18770
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 22020 17610 22048 22320
rect 22008 17604 22060 17610
rect 22008 17546 22060 17552
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 22480 14346 22508 22320
rect 22468 14340 22520 14346
rect 22468 14282 22520 14288
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19156 13320 19208 13326
rect 19156 13262 19208 13268
rect 19168 12986 19196 13262
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19444 11529 19472 13330
rect 19430 11520 19486 11529
rect 19430 11455 19486 11464
rect 18786 9616 18842 9625
rect 18786 9551 18842 9560
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 16316 4826 16344 7278
rect 16500 6254 16528 8502
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16592 6186 16620 7142
rect 16580 6180 16632 6186
rect 16580 6122 16632 6128
rect 16394 5808 16450 5817
rect 16394 5743 16450 5752
rect 16408 5642 16436 5743
rect 16396 5636 16448 5642
rect 16396 5578 16448 5584
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16394 4448 16450 4457
rect 16224 4406 16344 4434
rect 16210 4176 16266 4185
rect 16210 4111 16266 4120
rect 16224 4078 16252 4111
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16316 3738 16344 4406
rect 16394 4383 16450 4392
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16408 2990 16436 4383
rect 16580 4208 16632 4214
rect 16580 4150 16632 4156
rect 16396 2984 16448 2990
rect 16396 2926 16448 2932
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 16118 2544 16174 2553
rect 15844 2508 15896 2514
rect 16118 2479 16120 2488
rect 15844 2450 15896 2456
rect 16172 2479 16174 2488
rect 16120 2450 16172 2456
rect 16028 2372 16080 2378
rect 16028 2314 16080 2320
rect 15580 1992 15792 2020
rect 15580 480 15608 1992
rect 16040 480 16068 2314
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16500 480 16528 2246
rect 16592 1970 16620 4150
rect 16684 3602 16712 8230
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 16762 6352 16818 6361
rect 16762 6287 16764 6296
rect 16816 6287 16818 6296
rect 16764 6258 16816 6264
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 19800 5704 19852 5710
rect 19800 5646 19852 5652
rect 17498 5536 17554 5545
rect 17498 5471 17554 5480
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16764 4752 16816 4758
rect 16764 4694 16816 4700
rect 16776 3942 16804 4694
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16868 2446 16896 4966
rect 17420 4622 17448 5170
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17408 3460 17460 3466
rect 17408 3402 17460 3408
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 16580 1964 16632 1970
rect 16580 1906 16632 1912
rect 16960 480 16988 3334
rect 17328 1766 17356 3334
rect 17316 1760 17368 1766
rect 17316 1702 17368 1708
rect 17420 480 17448 3402
rect 17512 2514 17540 5471
rect 17972 4690 18000 5646
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 19812 5166 19840 5646
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 17960 4684 18012 4690
rect 17960 4626 18012 4632
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 17788 2650 17816 2858
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 17880 480 17908 2790
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17972 1170 18000 2246
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1142 18368 1170
rect 18340 480 18368 1142
rect 18800 480 18828 4422
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 19708 3120 19760 3126
rect 19708 3062 19760 3068
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 19260 480 19288 2790
rect 19720 480 19748 3062
rect 20180 480 20208 3470
rect 20640 480 20668 4966
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 21548 2916 21600 2922
rect 21548 2858 21600 2864
rect 21088 2100 21140 2106
rect 21088 2042 21140 2048
rect 21100 480 21128 2042
rect 21560 480 21588 2858
rect 22020 480 22048 3130
rect 22480 480 22508 3878
rect 4066 232 4122 241
rect 4066 167 4122 176
rect 4342 0 4398 480
rect 4802 0 4858 480
rect 5262 0 5318 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6642 0 6698 480
rect 7102 0 7158 480
rect 7562 0 7618 480
rect 8114 0 8170 480
rect 8574 0 8630 480
rect 9034 0 9090 480
rect 9494 0 9550 480
rect 9954 0 10010 480
rect 10414 0 10470 480
rect 10874 0 10930 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12254 0 12310 480
rect 12714 0 12770 480
rect 13174 0 13230 480
rect 13634 0 13690 480
rect 14094 0 14150 480
rect 14554 0 14610 480
rect 15014 0 15070 480
rect 15566 0 15622 480
rect 16026 0 16082 480
rect 16486 0 16542 480
rect 16946 0 17002 480
rect 17406 0 17462 480
rect 17866 0 17922 480
rect 18326 0 18382 480
rect 18786 0 18842 480
rect 19246 0 19302 480
rect 19706 0 19762 480
rect 20166 0 20222 480
rect 20626 0 20682 480
rect 21086 0 21142 480
rect 21546 0 21602 480
rect 22006 0 22062 480
rect 22466 0 22522 480
<< via2 >>
rect 3514 22480 3570 22536
rect 1858 18672 1914 18728
rect 1766 18264 1822 18320
rect 2318 18944 2374 19000
rect 1950 17312 2006 17368
rect 1674 16768 1730 16824
rect 1674 16396 1676 16416
rect 1676 16396 1728 16416
rect 1728 16396 1730 16416
rect 1674 16360 1730 16396
rect 1582 15816 1638 15872
rect 1582 15408 1638 15464
rect 1582 14864 1638 14920
rect 2410 18808 2466 18864
rect 2502 18708 2504 18728
rect 2504 18708 2556 18728
rect 2556 18708 2558 18728
rect 2502 18672 2558 18708
rect 3330 22072 3386 22128
rect 3330 20576 3386 20632
rect 2594 18264 2650 18320
rect 2042 13640 2098 13696
rect 1950 11736 2006 11792
rect 2042 10648 2098 10704
rect 2778 16768 2834 16824
rect 3514 17720 3570 17776
rect 2962 14900 2964 14920
rect 2964 14900 3016 14920
rect 3016 14900 3018 14920
rect 2962 14864 3018 14900
rect 2594 14728 2650 14784
rect 2778 14456 2834 14512
rect 2502 14320 2558 14376
rect 2870 13912 2926 13968
rect 2962 13776 3018 13832
rect 2962 13676 2964 13696
rect 2964 13676 3016 13696
rect 3016 13676 3018 13696
rect 2962 13640 3018 13676
rect 3238 13504 3294 13560
rect 1950 9560 2006 9616
rect 1858 9424 1914 9480
rect 2134 9288 2190 9344
rect 2226 4120 2282 4176
rect 2410 3712 2466 3768
rect 2226 3032 2282 3088
rect 2134 2488 2190 2544
rect 3606 15544 3662 15600
rect 3606 14592 3662 14648
rect 3238 12144 3294 12200
rect 3238 10648 3294 10704
rect 2962 7248 3018 7304
rect 4066 21528 4122 21584
rect 3974 21120 4030 21176
rect 4066 20204 4068 20224
rect 4068 20204 4120 20224
rect 4120 20204 4122 20224
rect 4066 20168 4122 20204
rect 4066 19624 4122 19680
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4066 19216 4122 19272
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4158 14864 4214 14920
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 3974 12552 4030 12608
rect 3974 12008 4030 12064
rect 2594 3032 2650 3088
rect 3054 3984 3110 4040
rect 2962 3168 3018 3224
rect 3422 4564 3424 4584
rect 3424 4564 3476 4584
rect 3476 4564 3478 4584
rect 3422 4528 3478 4564
rect 3882 11620 3938 11656
rect 3882 11600 3884 11620
rect 3884 11600 3936 11620
rect 3936 11600 3938 11620
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4802 12552 4858 12608
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4618 11600 4674 11656
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4066 9696 4122 9752
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 3606 6840 3662 6896
rect 3790 6296 3846 6352
rect 3790 4392 3846 4448
rect 3422 3440 3478 3496
rect 1950 1536 2006 1592
rect 3698 2524 3700 2544
rect 3700 2524 3752 2544
rect 3752 2524 3754 2544
rect 3698 2488 3754 2524
rect 3330 584 3386 640
rect 4066 8744 4122 8800
rect 4526 8880 4582 8936
rect 5814 18944 5870 19000
rect 5354 14592 5410 14648
rect 5170 13776 5226 13832
rect 5078 12416 5134 12472
rect 5262 11872 5318 11928
rect 5170 11464 5226 11520
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4250 8200 4306 8256
rect 4066 7792 4122 7848
rect 3974 5888 4030 5944
rect 3974 5344 4030 5400
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4802 4936 4858 4992
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4066 3440 4122 3496
rect 4158 3168 4214 3224
rect 4158 1536 4214 1592
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 3974 1164 3976 1184
rect 3976 1164 4028 1184
rect 4028 1164 4030 1184
rect 3974 1128 4030 1164
rect 5170 8744 5226 8800
rect 5906 11464 5962 11520
rect 5998 11056 6054 11112
rect 5446 9288 5502 9344
rect 5630 8472 5686 8528
rect 6182 8472 6238 8528
rect 5170 3304 5226 3360
rect 5078 2624 5134 2680
rect 5630 2760 5686 2816
rect 6090 5616 6146 5672
rect 7378 17720 7434 17776
rect 6826 14900 6828 14920
rect 6828 14900 6880 14920
rect 6880 14900 6882 14920
rect 6826 14864 6882 14900
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 8022 18672 8078 18728
rect 7838 18284 7894 18320
rect 7838 18264 7840 18284
rect 7840 18264 7892 18284
rect 7892 18264 7894 18284
rect 8114 18128 8170 18184
rect 7654 16768 7710 16824
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 8298 18808 8354 18864
rect 7838 17756 7840 17776
rect 7840 17756 7892 17776
rect 7892 17756 7894 17776
rect 7838 17720 7894 17756
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7838 16632 7894 16688
rect 8482 18128 8538 18184
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7838 15444 7840 15464
rect 7840 15444 7892 15464
rect 7892 15444 7894 15464
rect 7838 15408 7894 15444
rect 7746 14864 7802 14920
rect 6826 9596 6828 9616
rect 6828 9596 6880 9616
rect 6880 9596 6882 9616
rect 6826 9560 6882 9596
rect 5906 3168 5962 3224
rect 5814 2644 5870 2680
rect 5814 2624 5816 2644
rect 5816 2624 5868 2644
rect 5868 2624 5870 2644
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 8298 12824 8354 12880
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7654 12436 7710 12472
rect 7654 12416 7656 12436
rect 7656 12416 7708 12436
rect 7708 12416 7710 12436
rect 8666 18264 8722 18320
rect 9862 19216 9918 19272
rect 8758 15544 8814 15600
rect 7102 9152 7158 9208
rect 7378 8880 7434 8936
rect 6642 3712 6698 3768
rect 6182 3440 6238 3496
rect 7930 11600 7986 11656
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 8666 11192 8722 11248
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 8390 8744 8446 8800
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7286 4392 7342 4448
rect 7470 3984 7526 4040
rect 7194 3576 7250 3632
rect 6642 2896 6698 2952
rect 7286 2760 7342 2816
rect 7286 2488 7342 2544
rect 7746 4664 7802 4720
rect 8390 5480 8446 5536
rect 8482 4800 8538 4856
rect 9034 16652 9090 16688
rect 9034 16632 9036 16652
rect 9036 16632 9088 16652
rect 9088 16632 9090 16652
rect 10230 18944 10286 19000
rect 9034 15408 9090 15464
rect 9494 14320 9550 14376
rect 8850 11328 8906 11384
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 8298 3848 8354 3904
rect 8666 4120 8722 4176
rect 8298 3304 8354 3360
rect 9218 10104 9274 10160
rect 9126 8744 9182 8800
rect 9034 5616 9090 5672
rect 8942 4392 8998 4448
rect 9218 4664 9274 4720
rect 9586 11872 9642 11928
rect 9586 11736 9642 11792
rect 9862 12280 9918 12336
rect 9770 9696 9826 9752
rect 9770 9288 9826 9344
rect 9678 5888 9734 5944
rect 9586 5480 9642 5536
rect 9954 8200 10010 8256
rect 10046 7268 10102 7304
rect 10046 7248 10048 7268
rect 10048 7248 10100 7268
rect 10100 7248 10102 7268
rect 9954 6840 10010 6896
rect 9954 4392 10010 4448
rect 9678 3712 9734 3768
rect 9862 3712 9918 3768
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 11610 18944 11666 19000
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 10506 9152 10562 9208
rect 10598 7792 10654 7848
rect 10506 6704 10562 6760
rect 10506 5616 10562 5672
rect 10322 3712 10378 3768
rect 10506 3576 10562 3632
rect 11058 13912 11114 13968
rect 10874 10648 10930 10704
rect 11518 16668 11520 16688
rect 11520 16668 11572 16688
rect 11572 16668 11574 16688
rect 11518 16632 11574 16668
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11518 13932 11574 13968
rect 11518 13912 11520 13932
rect 11520 13912 11572 13932
rect 11572 13912 11574 13932
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11426 11328 11482 11384
rect 11334 11092 11336 11112
rect 11336 11092 11388 11112
rect 11388 11092 11390 11112
rect 11334 11056 11390 11092
rect 13082 16632 13138 16688
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11518 9152 11574 9208
rect 11334 9016 11390 9072
rect 11058 8744 11114 8800
rect 11058 8336 11114 8392
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11518 7928 11574 7984
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 10966 5228 11022 5264
rect 10966 5208 10968 5228
rect 10968 5208 11020 5228
rect 11020 5208 11022 5228
rect 10966 4684 11022 4720
rect 10966 4664 10968 4684
rect 10968 4664 11020 4684
rect 11020 4664 11022 4684
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11426 6296 11482 6352
rect 10966 4392 11022 4448
rect 10138 2488 10194 2544
rect 10322 2352 10378 2408
rect 11058 4256 11114 4312
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 10966 3168 11022 3224
rect 10966 2760 11022 2816
rect 11518 3576 11574 3632
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 10874 2216 10930 2272
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 11886 9696 11942 9752
rect 12254 11348 12310 11384
rect 12254 11328 12256 11348
rect 12256 11328 12308 11348
rect 12308 11328 12310 11348
rect 12162 11192 12218 11248
rect 12162 9696 12218 9752
rect 11978 9288 12034 9344
rect 12254 8064 12310 8120
rect 11794 4256 11850 4312
rect 11794 3712 11850 3768
rect 11794 3168 11850 3224
rect 12070 5344 12126 5400
rect 12070 4800 12126 4856
rect 12070 4120 12126 4176
rect 12438 11192 12494 11248
rect 12438 10140 12440 10160
rect 12440 10140 12492 10160
rect 12492 10140 12494 10160
rect 12438 10104 12494 10140
rect 12990 11056 13046 11112
rect 12898 9152 12954 9208
rect 13266 10104 13322 10160
rect 13174 8880 13230 8936
rect 13358 8200 13414 8256
rect 13818 18944 13874 19000
rect 13634 10648 13690 10704
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 15198 13932 15254 13968
rect 15198 13912 15200 13932
rect 15200 13912 15252 13932
rect 15252 13912 15254 13932
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 13726 9324 13728 9344
rect 13728 9324 13780 9344
rect 13780 9324 13782 9344
rect 13726 9288 13782 9324
rect 12346 5072 12402 5128
rect 12438 4972 12440 4992
rect 12440 4972 12492 4992
rect 12492 4972 12494 4992
rect 12438 4936 12494 4972
rect 12438 4800 12494 4856
rect 12346 3984 12402 4040
rect 12898 4936 12954 4992
rect 12254 3712 12310 3768
rect 12070 2488 12126 2544
rect 12714 3712 12770 3768
rect 12622 2760 12678 2816
rect 12990 3712 13046 3768
rect 13450 5344 13506 5400
rect 13450 4664 13506 4720
rect 12990 2896 13046 2952
rect 12990 2488 13046 2544
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14094 8608 14150 8664
rect 14002 6840 14058 6896
rect 13818 5208 13874 5264
rect 14094 5752 14150 5808
rect 14094 5616 14150 5672
rect 13910 4664 13966 4720
rect 13910 4528 13966 4584
rect 13726 3712 13782 3768
rect 14462 9424 14518 9480
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 15014 8492 15070 8528
rect 15014 8472 15016 8492
rect 15016 8472 15068 8492
rect 15068 8472 15070 8492
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14554 7792 14610 7848
rect 14462 6704 14518 6760
rect 14278 6160 14334 6216
rect 15382 9016 15438 9072
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 15014 5616 15070 5672
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14278 4800 14334 4856
rect 14646 4664 14702 4720
rect 14370 3884 14372 3904
rect 14372 3884 14424 3904
rect 14424 3884 14426 3904
rect 14370 3848 14426 3884
rect 14278 3712 14334 3768
rect 14094 3576 14150 3632
rect 14002 2932 14004 2952
rect 14004 2932 14056 2952
rect 14056 2932 14058 2952
rect 14002 2896 14058 2932
rect 14370 3440 14426 3496
rect 14646 4004 14702 4040
rect 14646 3984 14648 4004
rect 14648 3984 14700 4004
rect 14700 3984 14702 4004
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14646 3052 14702 3088
rect 14646 3032 14648 3052
rect 14648 3032 14700 3052
rect 14700 3032 14702 3052
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 15198 3596 15254 3632
rect 15198 3576 15200 3596
rect 15200 3576 15252 3596
rect 15252 3576 15254 3596
rect 15474 5072 15530 5128
rect 15750 8336 15806 8392
rect 15934 7268 15990 7304
rect 15934 7248 15936 7268
rect 15936 7248 15988 7268
rect 15988 7248 15990 7268
rect 15382 2896 15438 2952
rect 15198 2352 15254 2408
rect 16026 5072 16082 5128
rect 16026 4256 16082 4312
rect 17038 12280 17094 12336
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 19430 11464 19486 11520
rect 18786 9560 18842 9616
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 16394 5752 16450 5808
rect 16210 4120 16266 4176
rect 16394 4392 16450 4448
rect 16118 2508 16174 2544
rect 16118 2488 16120 2508
rect 16120 2488 16172 2508
rect 16172 2488 16174 2508
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 16762 6316 16818 6352
rect 16762 6296 16764 6316
rect 16764 6296 16816 6316
rect 16816 6296 16818 6316
rect 17498 5480 17554 5536
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 4066 176 4122 232
<< metal3 >>
rect 0 22538 480 22568
rect 3509 22538 3575 22541
rect 0 22536 3575 22538
rect 0 22480 3514 22536
rect 3570 22480 3575 22536
rect 0 22478 3575 22480
rect 0 22448 480 22478
rect 3509 22475 3575 22478
rect 0 22130 480 22160
rect 3325 22130 3391 22133
rect 0 22128 3391 22130
rect 0 22072 3330 22128
rect 3386 22072 3391 22128
rect 0 22070 3391 22072
rect 0 22040 480 22070
rect 3325 22067 3391 22070
rect 0 21586 480 21616
rect 4061 21586 4127 21589
rect 0 21584 4127 21586
rect 0 21528 4066 21584
rect 4122 21528 4127 21584
rect 0 21526 4127 21528
rect 0 21496 480 21526
rect 4061 21523 4127 21526
rect 0 21178 480 21208
rect 3969 21178 4035 21181
rect 0 21176 4035 21178
rect 0 21120 3974 21176
rect 4030 21120 4035 21176
rect 0 21118 4035 21120
rect 0 21088 480 21118
rect 3969 21115 4035 21118
rect 0 20634 480 20664
rect 3325 20634 3391 20637
rect 0 20632 3391 20634
rect 0 20576 3330 20632
rect 3386 20576 3391 20632
rect 0 20574 3391 20576
rect 0 20544 480 20574
rect 3325 20571 3391 20574
rect 0 20226 480 20256
rect 4061 20226 4127 20229
rect 0 20224 4127 20226
rect 0 20168 4066 20224
rect 4122 20168 4127 20224
rect 0 20166 4127 20168
rect 0 20136 480 20166
rect 4061 20163 4127 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 20095 14992 20096
rect 0 19682 480 19712
rect 4061 19682 4127 19685
rect 0 19680 4127 19682
rect 0 19624 4066 19680
rect 4122 19624 4127 19680
rect 0 19622 4127 19624
rect 0 19592 480 19622
rect 4061 19619 4127 19622
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 480 19304
rect 4061 19274 4127 19277
rect 0 19272 4127 19274
rect 0 19216 4066 19272
rect 4122 19216 4127 19272
rect 0 19214 4127 19216
rect 0 19184 480 19214
rect 4061 19211 4127 19214
rect 9857 19274 9923 19277
rect 9857 19272 15210 19274
rect 9857 19216 9862 19272
rect 9918 19216 15210 19272
rect 9857 19214 15210 19216
rect 9857 19211 9923 19214
rect 15150 19138 15210 19214
rect 22320 19138 22800 19168
rect 15150 19078 22800 19138
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 22320 19048 22800 19078
rect 14672 19007 14992 19008
rect 2313 19002 2379 19005
rect 5809 19002 5875 19005
rect 2313 19000 5875 19002
rect 2313 18944 2318 19000
rect 2374 18944 5814 19000
rect 5870 18944 5875 19000
rect 2313 18942 5875 18944
rect 2313 18939 2379 18942
rect 5809 18939 5875 18942
rect 10225 19002 10291 19005
rect 11605 19002 11671 19005
rect 13813 19002 13879 19005
rect 10225 19000 13879 19002
rect 10225 18944 10230 19000
rect 10286 18944 11610 19000
rect 11666 18944 13818 19000
rect 13874 18944 13879 19000
rect 10225 18942 13879 18944
rect 10225 18939 10291 18942
rect 11605 18939 11671 18942
rect 13813 18939 13879 18942
rect 2405 18866 2471 18869
rect 8293 18866 8359 18869
rect 2405 18864 8359 18866
rect 2405 18808 2410 18864
rect 2466 18808 8298 18864
rect 8354 18808 8359 18864
rect 2405 18806 8359 18808
rect 2405 18803 2471 18806
rect 8293 18803 8359 18806
rect 0 18730 480 18760
rect 1853 18730 1919 18733
rect 0 18728 1919 18730
rect 0 18672 1858 18728
rect 1914 18672 1919 18728
rect 0 18670 1919 18672
rect 0 18640 480 18670
rect 1853 18667 1919 18670
rect 2497 18730 2563 18733
rect 8017 18730 8083 18733
rect 2497 18728 8083 18730
rect 2497 18672 2502 18728
rect 2558 18672 8022 18728
rect 8078 18672 8083 18728
rect 2497 18670 8083 18672
rect 2497 18667 2563 18670
rect 8017 18667 8083 18670
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 480 18352
rect 1761 18322 1827 18325
rect 0 18320 1827 18322
rect 0 18264 1766 18320
rect 1822 18264 1827 18320
rect 0 18262 1827 18264
rect 0 18232 480 18262
rect 1761 18259 1827 18262
rect 2589 18322 2655 18325
rect 7833 18322 7899 18325
rect 8661 18322 8727 18325
rect 2589 18320 8727 18322
rect 2589 18264 2594 18320
rect 2650 18264 7838 18320
rect 7894 18264 8666 18320
rect 8722 18264 8727 18320
rect 2589 18262 8727 18264
rect 2589 18259 2655 18262
rect 7833 18259 7899 18262
rect 8661 18259 8727 18262
rect 8109 18186 8175 18189
rect 8477 18186 8543 18189
rect 8109 18184 8543 18186
rect 8109 18128 8114 18184
rect 8170 18128 8482 18184
rect 8538 18128 8543 18184
rect 8109 18126 8543 18128
rect 8109 18123 8175 18126
rect 8477 18123 8543 18126
rect 7808 17984 8128 17985
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 0 17778 480 17808
rect 3509 17778 3575 17781
rect 0 17776 3575 17778
rect 0 17720 3514 17776
rect 3570 17720 3575 17776
rect 0 17718 3575 17720
rect 0 17688 480 17718
rect 3509 17715 3575 17718
rect 7373 17778 7439 17781
rect 7833 17778 7899 17781
rect 7373 17776 7899 17778
rect 7373 17720 7378 17776
rect 7434 17720 7838 17776
rect 7894 17720 7899 17776
rect 7373 17718 7899 17720
rect 7373 17715 7439 17718
rect 7833 17715 7899 17718
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 1945 17370 2011 17373
rect 0 17368 2011 17370
rect 0 17312 1950 17368
rect 2006 17312 2011 17368
rect 0 17310 2011 17312
rect 0 17280 480 17310
rect 1945 17307 2011 17310
rect 7808 16896 8128 16897
rect 0 16826 480 16856
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 1669 16826 1735 16829
rect 0 16824 1735 16826
rect 0 16768 1674 16824
rect 1730 16768 1735 16824
rect 0 16766 1735 16768
rect 0 16736 480 16766
rect 1669 16763 1735 16766
rect 2773 16826 2839 16829
rect 7649 16826 7715 16829
rect 2773 16824 7715 16826
rect 2773 16768 2778 16824
rect 2834 16768 7654 16824
rect 7710 16768 7715 16824
rect 2773 16766 7715 16768
rect 2773 16763 2839 16766
rect 7649 16763 7715 16766
rect 7833 16690 7899 16693
rect 9029 16690 9095 16693
rect 7833 16688 9095 16690
rect 7833 16632 7838 16688
rect 7894 16632 9034 16688
rect 9090 16632 9095 16688
rect 7833 16630 9095 16632
rect 7833 16627 7899 16630
rect 9029 16627 9095 16630
rect 11513 16690 11579 16693
rect 13077 16690 13143 16693
rect 11513 16688 13143 16690
rect 11513 16632 11518 16688
rect 11574 16632 13082 16688
rect 13138 16632 13143 16688
rect 11513 16630 13143 16632
rect 11513 16627 11579 16630
rect 13077 16627 13143 16630
rect 0 16418 480 16448
rect 1669 16418 1735 16421
rect 0 16416 1735 16418
rect 0 16360 1674 16416
rect 1730 16360 1735 16416
rect 0 16358 1735 16360
rect 0 16328 480 16358
rect 1669 16355 1735 16358
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 0 15874 480 15904
rect 1577 15874 1643 15877
rect 0 15872 1643 15874
rect 0 15816 1582 15872
rect 1638 15816 1643 15872
rect 0 15814 1643 15816
rect 0 15784 480 15814
rect 1577 15811 1643 15814
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 3601 15602 3667 15605
rect 8753 15602 8819 15605
rect 3601 15600 8819 15602
rect 3601 15544 3606 15600
rect 3662 15544 8758 15600
rect 8814 15544 8819 15600
rect 3601 15542 8819 15544
rect 3601 15539 3667 15542
rect 8753 15539 8819 15542
rect 0 15466 480 15496
rect 1577 15466 1643 15469
rect 0 15464 1643 15466
rect 0 15408 1582 15464
rect 1638 15408 1643 15464
rect 0 15406 1643 15408
rect 0 15376 480 15406
rect 1577 15403 1643 15406
rect 7833 15466 7899 15469
rect 9029 15466 9095 15469
rect 7833 15464 9095 15466
rect 7833 15408 7838 15464
rect 7894 15408 9034 15464
rect 9090 15408 9095 15464
rect 7833 15406 9095 15408
rect 7833 15403 7899 15406
rect 9029 15403 9095 15406
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 14922 480 14952
rect 1577 14922 1643 14925
rect 0 14920 1643 14922
rect 0 14864 1582 14920
rect 1638 14864 1643 14920
rect 0 14862 1643 14864
rect 0 14832 480 14862
rect 1577 14859 1643 14862
rect 2957 14922 3023 14925
rect 4153 14922 4219 14925
rect 2957 14920 4219 14922
rect 2957 14864 2962 14920
rect 3018 14864 4158 14920
rect 4214 14864 4219 14920
rect 2957 14862 4219 14864
rect 2957 14859 3023 14862
rect 4153 14859 4219 14862
rect 6821 14922 6887 14925
rect 7741 14922 7807 14925
rect 6821 14920 7807 14922
rect 6821 14864 6826 14920
rect 6882 14864 7746 14920
rect 7802 14864 7807 14920
rect 6821 14862 7807 14864
rect 6821 14859 6887 14862
rect 7741 14859 7807 14862
rect 2589 14786 2655 14789
rect 2589 14784 3434 14786
rect 2589 14728 2594 14784
rect 2650 14728 3434 14784
rect 2589 14726 3434 14728
rect 2589 14723 2655 14726
rect 3374 14650 3434 14726
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 3601 14650 3667 14653
rect 5349 14650 5415 14653
rect 3374 14648 5415 14650
rect 3374 14592 3606 14648
rect 3662 14592 5354 14648
rect 5410 14592 5415 14648
rect 3374 14590 5415 14592
rect 3601 14587 3667 14590
rect 5349 14587 5415 14590
rect 0 14514 480 14544
rect 2773 14514 2839 14517
rect 0 14512 2839 14514
rect 0 14456 2778 14512
rect 2834 14456 2839 14512
rect 0 14454 2839 14456
rect 0 14424 480 14454
rect 2773 14451 2839 14454
rect 2497 14378 2563 14381
rect 9489 14378 9555 14381
rect 2497 14376 9555 14378
rect 2497 14320 2502 14376
rect 2558 14320 9494 14376
rect 9550 14320 9555 14376
rect 2497 14318 9555 14320
rect 2497 14315 2563 14318
rect 9489 14315 9555 14318
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 0 13970 480 14000
rect 2865 13970 2931 13973
rect 0 13968 2931 13970
rect 0 13912 2870 13968
rect 2926 13912 2931 13968
rect 0 13910 2931 13912
rect 0 13880 480 13910
rect 2865 13907 2931 13910
rect 11053 13970 11119 13973
rect 11513 13970 11579 13973
rect 15193 13970 15259 13973
rect 11053 13968 15259 13970
rect 11053 13912 11058 13968
rect 11114 13912 11518 13968
rect 11574 13912 15198 13968
rect 15254 13912 15259 13968
rect 11053 13910 15259 13912
rect 11053 13907 11119 13910
rect 11513 13907 11579 13910
rect 15193 13907 15259 13910
rect 2957 13834 3023 13837
rect 5165 13834 5231 13837
rect 2957 13832 5231 13834
rect 2957 13776 2962 13832
rect 3018 13776 5170 13832
rect 5226 13776 5231 13832
rect 2957 13774 5231 13776
rect 2957 13771 3023 13774
rect 5165 13771 5231 13774
rect 2037 13698 2103 13701
rect 2957 13698 3023 13701
rect 2037 13696 3023 13698
rect 2037 13640 2042 13696
rect 2098 13640 2962 13696
rect 3018 13640 3023 13696
rect 2037 13638 3023 13640
rect 2037 13635 2103 13638
rect 2957 13635 3023 13638
rect 7808 13632 8128 13633
rect 0 13562 480 13592
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 3233 13562 3299 13565
rect 0 13560 3299 13562
rect 0 13504 3238 13560
rect 3294 13504 3299 13560
rect 0 13502 3299 13504
rect 0 13472 480 13502
rect 3233 13499 3299 13502
rect 4376 13088 4696 13089
rect 0 13018 480 13048
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 0 12958 4170 13018
rect 0 12928 480 12958
rect 4110 12882 4170 12958
rect 8293 12882 8359 12885
rect 4110 12880 8359 12882
rect 4110 12824 8298 12880
rect 8354 12824 8359 12880
rect 4110 12822 8359 12824
rect 8293 12819 8359 12822
rect 0 12610 480 12640
rect 3969 12610 4035 12613
rect 0 12608 4035 12610
rect 0 12552 3974 12608
rect 4030 12552 4035 12608
rect 0 12550 4035 12552
rect 0 12520 480 12550
rect 3969 12547 4035 12550
rect 4797 12610 4863 12613
rect 5022 12610 5028 12612
rect 4797 12608 5028 12610
rect 4797 12552 4802 12608
rect 4858 12552 5028 12608
rect 4797 12550 5028 12552
rect 4797 12547 4863 12550
rect 5022 12548 5028 12550
rect 5092 12548 5098 12612
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 5073 12474 5139 12477
rect 7649 12474 7715 12477
rect 5073 12472 7715 12474
rect 5073 12416 5078 12472
rect 5134 12416 7654 12472
rect 7710 12416 7715 12472
rect 5073 12414 7715 12416
rect 5073 12411 5139 12414
rect 7649 12411 7715 12414
rect 9857 12338 9923 12341
rect 17033 12338 17099 12341
rect 9857 12336 17099 12338
rect 9857 12280 9862 12336
rect 9918 12280 17038 12336
rect 17094 12280 17099 12336
rect 9857 12278 17099 12280
rect 9857 12275 9923 12278
rect 17033 12275 17099 12278
rect 3233 12202 3299 12205
rect 3233 12200 4906 12202
rect 3233 12144 3238 12200
rect 3294 12144 4906 12200
rect 3233 12142 4906 12144
rect 3233 12139 3299 12142
rect 0 12066 480 12096
rect 3969 12066 4035 12069
rect 0 12064 4035 12066
rect 0 12008 3974 12064
rect 4030 12008 4035 12064
rect 0 12006 4035 12008
rect 0 11976 480 12006
rect 3969 12003 4035 12006
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 4846 11930 4906 12142
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 5257 11930 5323 11933
rect 9581 11930 9647 11933
rect 4846 11928 9647 11930
rect 4846 11872 5262 11928
rect 5318 11872 9586 11928
rect 9642 11872 9647 11928
rect 4846 11870 9647 11872
rect 5257 11867 5323 11870
rect 9581 11867 9647 11870
rect 1945 11794 2011 11797
rect 9581 11794 9647 11797
rect 1945 11792 9647 11794
rect 1945 11736 1950 11792
rect 2006 11736 9586 11792
rect 9642 11736 9647 11792
rect 1945 11734 9647 11736
rect 1945 11731 2011 11734
rect 9581 11731 9647 11734
rect 0 11658 480 11688
rect 3877 11658 3943 11661
rect 0 11656 3943 11658
rect 0 11600 3882 11656
rect 3938 11600 3943 11656
rect 0 11598 3943 11600
rect 0 11568 480 11598
rect 3877 11595 3943 11598
rect 4613 11658 4679 11661
rect 7925 11658 7991 11661
rect 4613 11656 7991 11658
rect 4613 11600 4618 11656
rect 4674 11600 7930 11656
rect 7986 11600 7991 11656
rect 4613 11598 7991 11600
rect 4613 11595 4679 11598
rect 7925 11595 7991 11598
rect 5165 11522 5231 11525
rect 5901 11522 5967 11525
rect 5165 11520 5967 11522
rect 5165 11464 5170 11520
rect 5226 11464 5906 11520
rect 5962 11464 5967 11520
rect 5165 11462 5967 11464
rect 5165 11459 5231 11462
rect 5901 11459 5967 11462
rect 19425 11522 19491 11525
rect 22320 11522 22800 11552
rect 19425 11520 22800 11522
rect 19425 11464 19430 11520
rect 19486 11464 22800 11520
rect 19425 11462 22800 11464
rect 19425 11459 19491 11462
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 22320 11432 22800 11462
rect 14672 11391 14992 11392
rect 8845 11386 8911 11389
rect 8710 11384 8911 11386
rect 8710 11328 8850 11384
rect 8906 11328 8911 11384
rect 8710 11326 8911 11328
rect 8710 11253 8770 11326
rect 8845 11323 8911 11326
rect 11421 11386 11487 11389
rect 12249 11386 12315 11389
rect 11421 11384 12315 11386
rect 11421 11328 11426 11384
rect 11482 11328 12254 11384
rect 12310 11328 12315 11384
rect 11421 11326 12315 11328
rect 11421 11323 11487 11326
rect 12249 11323 12315 11326
rect 8661 11248 8770 11253
rect 8661 11192 8666 11248
rect 8722 11192 8770 11248
rect 8661 11190 8770 11192
rect 12157 11250 12223 11253
rect 12433 11250 12499 11253
rect 12157 11248 12499 11250
rect 12157 11192 12162 11248
rect 12218 11192 12438 11248
rect 12494 11192 12499 11248
rect 12157 11190 12499 11192
rect 8661 11187 8727 11190
rect 12157 11187 12223 11190
rect 12433 11187 12499 11190
rect 0 11114 480 11144
rect 5993 11114 6059 11117
rect 0 11112 6059 11114
rect 0 11056 5998 11112
rect 6054 11056 6059 11112
rect 0 11054 6059 11056
rect 0 11024 480 11054
rect 5993 11051 6059 11054
rect 11329 11114 11395 11117
rect 12985 11114 13051 11117
rect 11329 11112 13051 11114
rect 11329 11056 11334 11112
rect 11390 11056 12990 11112
rect 13046 11056 13051 11112
rect 11329 11054 13051 11056
rect 11329 11051 11395 11054
rect 12985 11051 13051 11054
rect 4376 10912 4696 10913
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 0 10706 480 10736
rect 2037 10706 2103 10709
rect 3233 10706 3299 10709
rect 0 10704 3299 10706
rect 0 10648 2042 10704
rect 2098 10648 3238 10704
rect 3294 10648 3299 10704
rect 0 10646 3299 10648
rect 0 10616 480 10646
rect 2037 10643 2103 10646
rect 3233 10643 3299 10646
rect 10869 10706 10935 10709
rect 13629 10706 13695 10709
rect 10869 10704 13695 10706
rect 10869 10648 10874 10704
rect 10930 10648 13634 10704
rect 13690 10648 13695 10704
rect 10869 10646 13695 10648
rect 10869 10643 10935 10646
rect 13629 10643 13695 10646
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 0 10162 480 10192
rect 9213 10162 9279 10165
rect 0 10160 9279 10162
rect 0 10104 9218 10160
rect 9274 10104 9279 10160
rect 0 10102 9279 10104
rect 0 10072 480 10102
rect 9213 10099 9279 10102
rect 12433 10162 12499 10165
rect 13261 10162 13327 10165
rect 12433 10160 13327 10162
rect 12433 10104 12438 10160
rect 12494 10104 13266 10160
rect 13322 10104 13327 10160
rect 12433 10102 13327 10104
rect 12433 10099 12499 10102
rect 13261 10099 13327 10102
rect 4376 9824 4696 9825
rect 0 9754 480 9784
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 4061 9754 4127 9757
rect 9765 9754 9831 9757
rect 0 9752 4127 9754
rect 0 9696 4066 9752
rect 4122 9696 4127 9752
rect 0 9694 4127 9696
rect 0 9664 480 9694
rect 4061 9691 4127 9694
rect 5030 9752 9831 9754
rect 5030 9696 9770 9752
rect 9826 9696 9831 9752
rect 5030 9694 9831 9696
rect 1945 9618 2011 9621
rect 5030 9618 5090 9694
rect 9765 9691 9831 9694
rect 11881 9754 11947 9757
rect 12157 9754 12223 9757
rect 11881 9752 12223 9754
rect 11881 9696 11886 9752
rect 11942 9696 12162 9752
rect 12218 9696 12223 9752
rect 11881 9694 12223 9696
rect 11881 9691 11947 9694
rect 12157 9691 12223 9694
rect 1945 9616 5090 9618
rect 1945 9560 1950 9616
rect 2006 9560 5090 9616
rect 1945 9558 5090 9560
rect 6821 9618 6887 9621
rect 18781 9618 18847 9621
rect 6821 9616 18847 9618
rect 6821 9560 6826 9616
rect 6882 9560 18786 9616
rect 18842 9560 18847 9616
rect 6821 9558 18847 9560
rect 1945 9555 2011 9558
rect 6821 9555 6887 9558
rect 18781 9555 18847 9558
rect 1853 9482 1919 9485
rect 14457 9482 14523 9485
rect 1853 9480 14523 9482
rect 1853 9424 1858 9480
rect 1914 9424 14462 9480
rect 14518 9424 14523 9480
rect 1853 9422 14523 9424
rect 1853 9419 1919 9422
rect 14457 9419 14523 9422
rect 2129 9346 2195 9349
rect 5441 9346 5507 9349
rect 2129 9344 5507 9346
rect 2129 9288 2134 9344
rect 2190 9288 5446 9344
rect 5502 9288 5507 9344
rect 2129 9286 5507 9288
rect 2129 9283 2195 9286
rect 5441 9283 5507 9286
rect 9765 9346 9831 9349
rect 11973 9346 12039 9349
rect 13721 9346 13787 9349
rect 9765 9344 13787 9346
rect 9765 9288 9770 9344
rect 9826 9288 11978 9344
rect 12034 9288 13726 9344
rect 13782 9288 13787 9344
rect 9765 9286 13787 9288
rect 9765 9283 9831 9286
rect 11973 9283 12039 9286
rect 13721 9283 13787 9286
rect 7808 9280 8128 9281
rect 0 9210 480 9240
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 7097 9210 7163 9213
rect 0 9208 7163 9210
rect 0 9152 7102 9208
rect 7158 9152 7163 9208
rect 0 9150 7163 9152
rect 0 9120 480 9150
rect 7097 9147 7163 9150
rect 10501 9210 10567 9213
rect 11513 9210 11579 9213
rect 10501 9208 11579 9210
rect 10501 9152 10506 9208
rect 10562 9152 11518 9208
rect 11574 9152 11579 9208
rect 10501 9150 11579 9152
rect 10501 9147 10567 9150
rect 11513 9147 11579 9150
rect 12750 9148 12756 9212
rect 12820 9210 12826 9212
rect 12893 9210 12959 9213
rect 12820 9208 12959 9210
rect 12820 9152 12898 9208
rect 12954 9152 12959 9208
rect 12820 9150 12959 9152
rect 12820 9148 12826 9150
rect 12893 9147 12959 9150
rect 11329 9074 11395 9077
rect 15377 9074 15443 9077
rect 11329 9072 15443 9074
rect 11329 9016 11334 9072
rect 11390 9016 15382 9072
rect 15438 9016 15443 9072
rect 11329 9014 15443 9016
rect 11329 9011 11395 9014
rect 15377 9011 15443 9014
rect 4521 8938 4587 8941
rect 4838 8938 4844 8940
rect 4521 8936 4844 8938
rect 4521 8880 4526 8936
rect 4582 8880 4844 8936
rect 4521 8878 4844 8880
rect 4521 8875 4587 8878
rect 4838 8876 4844 8878
rect 4908 8876 4914 8940
rect 7373 8938 7439 8941
rect 13169 8938 13235 8941
rect 7373 8936 13235 8938
rect 7373 8880 7378 8936
rect 7434 8880 13174 8936
rect 13230 8880 13235 8936
rect 7373 8878 13235 8880
rect 7373 8875 7439 8878
rect 13169 8875 13235 8878
rect 0 8802 480 8832
rect 4061 8802 4127 8805
rect 0 8800 4127 8802
rect 0 8744 4066 8800
rect 4122 8744 4127 8800
rect 0 8742 4127 8744
rect 0 8712 480 8742
rect 4061 8739 4127 8742
rect 5022 8740 5028 8804
rect 5092 8802 5098 8804
rect 5165 8802 5231 8805
rect 5092 8800 5231 8802
rect 5092 8744 5170 8800
rect 5226 8744 5231 8800
rect 5092 8742 5231 8744
rect 5092 8740 5098 8742
rect 5165 8739 5231 8742
rect 8385 8802 8451 8805
rect 9121 8802 9187 8805
rect 11053 8802 11119 8805
rect 8385 8800 11119 8802
rect 8385 8744 8390 8800
rect 8446 8744 9126 8800
rect 9182 8744 11058 8800
rect 11114 8744 11119 8800
rect 8385 8742 11119 8744
rect 8385 8739 8451 8742
rect 9121 8739 9187 8742
rect 11053 8739 11119 8742
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 14089 8666 14155 8669
rect 14222 8666 14228 8668
rect 14089 8664 14228 8666
rect 14089 8608 14094 8664
rect 14150 8608 14228 8664
rect 14089 8606 14228 8608
rect 14089 8603 14155 8606
rect 14222 8604 14228 8606
rect 14292 8604 14298 8668
rect 5625 8530 5691 8533
rect 6177 8530 6243 8533
rect 15009 8530 15075 8533
rect 5625 8528 15075 8530
rect 5625 8472 5630 8528
rect 5686 8472 6182 8528
rect 6238 8472 15014 8528
rect 15070 8472 15075 8528
rect 5625 8470 15075 8472
rect 5625 8467 5691 8470
rect 6177 8467 6243 8470
rect 15009 8467 15075 8470
rect 11053 8394 11119 8397
rect 15745 8394 15811 8397
rect 11053 8392 15811 8394
rect 11053 8336 11058 8392
rect 11114 8336 15750 8392
rect 15806 8336 15811 8392
rect 11053 8334 15811 8336
rect 11053 8331 11119 8334
rect 15745 8331 15811 8334
rect 0 8258 480 8288
rect 4245 8258 4311 8261
rect 0 8256 4311 8258
rect 0 8200 4250 8256
rect 4306 8200 4311 8256
rect 0 8198 4311 8200
rect 0 8168 480 8198
rect 4245 8195 4311 8198
rect 9949 8258 10015 8261
rect 13353 8258 13419 8261
rect 9949 8256 13419 8258
rect 9949 8200 9954 8256
rect 10010 8200 13358 8256
rect 13414 8200 13419 8256
rect 9949 8198 13419 8200
rect 9949 8195 10015 8198
rect 13353 8195 13419 8198
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 10910 8060 10916 8124
rect 10980 8122 10986 8124
rect 12249 8122 12315 8125
rect 10980 8120 12315 8122
rect 10980 8064 12254 8120
rect 12310 8064 12315 8120
rect 10980 8062 12315 8064
rect 10980 8060 10986 8062
rect 12249 8059 12315 8062
rect 11513 7986 11579 7989
rect 13854 7986 13860 7988
rect 11513 7984 13860 7986
rect 11513 7928 11518 7984
rect 11574 7928 13860 7984
rect 11513 7926 13860 7928
rect 11513 7923 11579 7926
rect 13854 7924 13860 7926
rect 13924 7924 13930 7988
rect 0 7850 480 7880
rect 4061 7850 4127 7853
rect 0 7848 4127 7850
rect 0 7792 4066 7848
rect 4122 7792 4127 7848
rect 0 7790 4127 7792
rect 0 7760 480 7790
rect 4061 7787 4127 7790
rect 10593 7850 10659 7853
rect 14549 7850 14615 7853
rect 10593 7848 14615 7850
rect 10593 7792 10598 7848
rect 10654 7792 14554 7848
rect 14610 7792 14615 7848
rect 10593 7790 14615 7792
rect 10593 7787 10659 7790
rect 14549 7787 14615 7790
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 0 7306 480 7336
rect 2957 7306 3023 7309
rect 0 7304 3023 7306
rect 0 7248 2962 7304
rect 3018 7248 3023 7304
rect 0 7246 3023 7248
rect 0 7216 480 7246
rect 2957 7243 3023 7246
rect 10041 7306 10107 7309
rect 15929 7306 15995 7309
rect 10041 7304 15995 7306
rect 10041 7248 10046 7304
rect 10102 7248 15934 7304
rect 15990 7248 15995 7304
rect 10041 7246 15995 7248
rect 10041 7243 10107 7246
rect 15929 7243 15995 7246
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 0 6898 480 6928
rect 3601 6898 3667 6901
rect 0 6896 3667 6898
rect 0 6840 3606 6896
rect 3662 6840 3667 6896
rect 0 6838 3667 6840
rect 0 6808 480 6838
rect 3601 6835 3667 6838
rect 9949 6898 10015 6901
rect 13997 6898 14063 6901
rect 9949 6896 14063 6898
rect 9949 6840 9954 6896
rect 10010 6840 14002 6896
rect 14058 6840 14063 6896
rect 9949 6838 14063 6840
rect 9949 6835 10015 6838
rect 13997 6835 14063 6838
rect 10501 6762 10567 6765
rect 14457 6762 14523 6765
rect 10501 6760 14523 6762
rect 10501 6704 10506 6760
rect 10562 6704 14462 6760
rect 14518 6704 14523 6760
rect 10501 6702 14523 6704
rect 10501 6699 10567 6702
rect 14457 6699 14523 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 0 6354 480 6384
rect 3785 6354 3851 6357
rect 0 6352 3851 6354
rect 0 6296 3790 6352
rect 3846 6296 3851 6352
rect 0 6294 3851 6296
rect 0 6264 480 6294
rect 3785 6291 3851 6294
rect 11421 6354 11487 6357
rect 16757 6354 16823 6357
rect 11421 6352 16823 6354
rect 11421 6296 11426 6352
rect 11482 6296 16762 6352
rect 16818 6296 16823 6352
rect 11421 6294 16823 6296
rect 11421 6291 11487 6294
rect 16757 6291 16823 6294
rect 12198 6156 12204 6220
rect 12268 6218 12274 6220
rect 14273 6218 14339 6221
rect 12268 6216 14339 6218
rect 12268 6160 14278 6216
rect 14334 6160 14339 6216
rect 12268 6158 14339 6160
rect 12268 6156 12274 6158
rect 14273 6155 14339 6158
rect 7808 6016 8128 6017
rect 0 5946 480 5976
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 3969 5946 4035 5949
rect 0 5944 4035 5946
rect 0 5888 3974 5944
rect 4030 5888 4035 5944
rect 0 5886 4035 5888
rect 0 5856 480 5886
rect 3969 5883 4035 5886
rect 9673 5946 9739 5949
rect 9673 5944 14290 5946
rect 9673 5888 9678 5944
rect 9734 5888 14290 5944
rect 9673 5886 14290 5888
rect 9673 5883 9739 5886
rect 14089 5810 14155 5813
rect 10550 5808 14155 5810
rect 10550 5752 14094 5808
rect 14150 5752 14155 5808
rect 10550 5750 14155 5752
rect 14230 5810 14290 5886
rect 16389 5810 16455 5813
rect 14230 5808 16455 5810
rect 14230 5752 16394 5808
rect 16450 5752 16455 5808
rect 14230 5750 16455 5752
rect 10550 5677 10610 5750
rect 14089 5747 14155 5750
rect 16389 5747 16455 5750
rect 6085 5674 6151 5677
rect 9029 5674 9095 5677
rect 6085 5672 9095 5674
rect 6085 5616 6090 5672
rect 6146 5616 9034 5672
rect 9090 5616 9095 5672
rect 6085 5614 9095 5616
rect 6085 5611 6151 5614
rect 9029 5611 9095 5614
rect 10501 5672 10610 5677
rect 14089 5674 14155 5677
rect 15009 5674 15075 5677
rect 10501 5616 10506 5672
rect 10562 5616 10610 5672
rect 10501 5614 10610 5616
rect 11102 5614 11714 5674
rect 10501 5611 10567 5614
rect 8385 5538 8451 5541
rect 9581 5538 9647 5541
rect 11102 5538 11162 5614
rect 8385 5536 11162 5538
rect 8385 5480 8390 5536
rect 8446 5480 9586 5536
rect 9642 5480 11162 5536
rect 8385 5478 11162 5480
rect 11654 5538 11714 5614
rect 14089 5672 15075 5674
rect 14089 5616 14094 5672
rect 14150 5616 15014 5672
rect 15070 5616 15075 5672
rect 14089 5614 15075 5616
rect 14089 5611 14155 5614
rect 15009 5611 15075 5614
rect 17493 5538 17559 5541
rect 11654 5536 17559 5538
rect 11654 5480 17498 5536
rect 17554 5480 17559 5536
rect 11654 5478 17559 5480
rect 8385 5475 8451 5478
rect 9581 5475 9647 5478
rect 17493 5475 17559 5478
rect 4376 5472 4696 5473
rect 0 5402 480 5432
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 3969 5402 4035 5405
rect 0 5400 4035 5402
rect 0 5344 3974 5400
rect 4030 5344 4035 5400
rect 0 5342 4035 5344
rect 0 5312 480 5342
rect 3969 5339 4035 5342
rect 12065 5402 12131 5405
rect 13445 5402 13511 5405
rect 12065 5400 13511 5402
rect 12065 5344 12070 5400
rect 12126 5344 13450 5400
rect 13506 5344 13511 5400
rect 12065 5342 13511 5344
rect 12065 5339 12131 5342
rect 13445 5339 13511 5342
rect 10961 5266 11027 5269
rect 13813 5266 13879 5269
rect 10961 5264 13879 5266
rect 10961 5208 10966 5264
rect 11022 5208 13818 5264
rect 13874 5208 13879 5264
rect 10961 5206 13879 5208
rect 10961 5203 11027 5206
rect 13813 5203 13879 5206
rect 12341 5130 12407 5133
rect 15469 5130 15535 5133
rect 16021 5130 16087 5133
rect 12341 5128 16087 5130
rect 12341 5072 12346 5128
rect 12402 5072 15474 5128
rect 15530 5072 16026 5128
rect 16082 5072 16087 5128
rect 12341 5070 16087 5072
rect 12341 5067 12407 5070
rect 15469 5067 15535 5070
rect 16021 5067 16087 5070
rect 0 4994 480 5024
rect 4797 4994 4863 4997
rect 0 4992 4863 4994
rect 0 4936 4802 4992
rect 4858 4936 4863 4992
rect 0 4934 4863 4936
rect 0 4904 480 4934
rect 4797 4931 4863 4934
rect 12433 4994 12499 4997
rect 12893 4994 12959 4997
rect 12433 4992 12959 4994
rect 12433 4936 12438 4992
rect 12494 4936 12898 4992
rect 12954 4936 12959 4992
rect 12433 4934 12959 4936
rect 12433 4931 12499 4934
rect 12893 4931 12959 4934
rect 7808 4928 8128 4929
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 8477 4858 8543 4861
rect 12065 4858 12131 4861
rect 8477 4856 12131 4858
rect 8477 4800 8482 4856
rect 8538 4800 12070 4856
rect 12126 4800 12131 4856
rect 8477 4798 12131 4800
rect 8477 4795 8543 4798
rect 12065 4795 12131 4798
rect 12433 4858 12499 4861
rect 14273 4858 14339 4861
rect 12433 4856 14339 4858
rect 12433 4800 12438 4856
rect 12494 4800 14278 4856
rect 14334 4800 14339 4856
rect 12433 4798 14339 4800
rect 12433 4795 12499 4798
rect 14273 4795 14339 4798
rect 7741 4722 7807 4725
rect 9213 4722 9279 4725
rect 7741 4720 9279 4722
rect 7741 4664 7746 4720
rect 7802 4664 9218 4720
rect 9274 4664 9279 4720
rect 7741 4662 9279 4664
rect 7741 4659 7807 4662
rect 9213 4659 9279 4662
rect 10961 4722 11027 4725
rect 13445 4722 13511 4725
rect 10961 4720 13511 4722
rect 10961 4664 10966 4720
rect 11022 4664 13450 4720
rect 13506 4664 13511 4720
rect 10961 4662 13511 4664
rect 10961 4659 11027 4662
rect 13445 4659 13511 4662
rect 13905 4722 13971 4725
rect 14641 4722 14707 4725
rect 13905 4720 14707 4722
rect 13905 4664 13910 4720
rect 13966 4664 14646 4720
rect 14702 4664 14707 4720
rect 13905 4662 14707 4664
rect 13905 4659 13971 4662
rect 14641 4659 14707 4662
rect 3417 4586 3483 4589
rect 13905 4586 13971 4589
rect 3417 4584 13971 4586
rect 3417 4528 3422 4584
rect 3478 4528 13910 4584
rect 13966 4528 13971 4584
rect 3417 4526 13971 4528
rect 3417 4523 3483 4526
rect 13905 4523 13971 4526
rect 0 4450 480 4480
rect 3785 4450 3851 4453
rect 0 4448 3851 4450
rect 0 4392 3790 4448
rect 3846 4392 3851 4448
rect 0 4390 3851 4392
rect 0 4360 480 4390
rect 3785 4387 3851 4390
rect 7281 4450 7347 4453
rect 8937 4450 9003 4453
rect 7281 4448 9003 4450
rect 7281 4392 7286 4448
rect 7342 4392 8942 4448
rect 8998 4392 9003 4448
rect 7281 4390 9003 4392
rect 7281 4387 7347 4390
rect 8937 4387 9003 4390
rect 9949 4450 10015 4453
rect 10961 4450 11027 4453
rect 16389 4450 16455 4453
rect 9949 4448 11027 4450
rect 9949 4392 9954 4448
rect 10010 4392 10966 4448
rect 11022 4392 11027 4448
rect 9949 4390 11027 4392
rect 9949 4387 10015 4390
rect 10961 4387 11027 4390
rect 11654 4448 16455 4450
rect 11654 4392 16394 4448
rect 16450 4392 16455 4448
rect 11654 4390 16455 4392
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 4838 4314 4844 4316
rect 4800 4252 4844 4314
rect 4908 4314 4914 4316
rect 11053 4314 11119 4317
rect 4908 4312 11119 4314
rect 4908 4256 11058 4312
rect 11114 4256 11119 4312
rect 4908 4254 11119 4256
rect 4908 4252 4914 4254
rect 2221 4178 2287 4181
rect 4800 4178 4860 4252
rect 11053 4251 11119 4254
rect 2221 4176 4860 4178
rect 2221 4120 2226 4176
rect 2282 4120 4860 4176
rect 2221 4118 4860 4120
rect 8661 4178 8727 4181
rect 11654 4178 11714 4390
rect 16389 4387 16455 4390
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 11789 4314 11855 4317
rect 16021 4314 16087 4317
rect 11789 4312 16087 4314
rect 11789 4256 11794 4312
rect 11850 4256 16026 4312
rect 16082 4256 16087 4312
rect 11789 4254 16087 4256
rect 11789 4251 11855 4254
rect 16021 4251 16087 4254
rect 8661 4176 11714 4178
rect 8661 4120 8666 4176
rect 8722 4120 11714 4176
rect 8661 4118 11714 4120
rect 12065 4178 12131 4181
rect 16205 4178 16271 4181
rect 12065 4176 16271 4178
rect 12065 4120 12070 4176
rect 12126 4120 16210 4176
rect 16266 4120 16271 4176
rect 12065 4118 16271 4120
rect 2221 4115 2287 4118
rect 8661 4115 8727 4118
rect 12065 4115 12131 4118
rect 16205 4115 16271 4118
rect 0 4042 480 4072
rect 3049 4042 3115 4045
rect 0 4040 3115 4042
rect 0 3984 3054 4040
rect 3110 3984 3115 4040
rect 0 3982 3115 3984
rect 0 3952 480 3982
rect 3049 3979 3115 3982
rect 7465 4042 7531 4045
rect 12198 4042 12204 4044
rect 7465 4040 12204 4042
rect 7465 3984 7470 4040
rect 7526 3984 12204 4040
rect 7465 3982 12204 3984
rect 7465 3979 7531 3982
rect 12198 3980 12204 3982
rect 12268 3980 12274 4044
rect 12341 4042 12407 4045
rect 14641 4042 14707 4045
rect 12341 4040 14707 4042
rect 12341 3984 12346 4040
rect 12402 3984 14646 4040
rect 14702 3984 14707 4040
rect 12341 3982 14707 3984
rect 12341 3979 12407 3982
rect 14641 3979 14707 3982
rect 8293 3906 8359 3909
rect 14365 3906 14431 3909
rect 22320 3906 22800 3936
rect 8293 3904 14431 3906
rect 8293 3848 8298 3904
rect 8354 3848 14370 3904
rect 14426 3848 14431 3904
rect 8293 3846 14431 3848
rect 8293 3843 8359 3846
rect 14365 3843 14431 3846
rect 17358 3846 22800 3906
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 2405 3770 2471 3773
rect 6637 3770 6703 3773
rect 2405 3768 6703 3770
rect 2405 3712 2410 3768
rect 2466 3712 6642 3768
rect 6698 3712 6703 3768
rect 2405 3710 6703 3712
rect 2405 3707 2471 3710
rect 6637 3707 6703 3710
rect 9673 3770 9739 3773
rect 9857 3770 9923 3773
rect 9673 3768 9923 3770
rect 9673 3712 9678 3768
rect 9734 3712 9862 3768
rect 9918 3712 9923 3768
rect 9673 3710 9923 3712
rect 9673 3707 9739 3710
rect 9857 3707 9923 3710
rect 10317 3770 10383 3773
rect 11789 3770 11855 3773
rect 10317 3768 11855 3770
rect 10317 3712 10322 3768
rect 10378 3712 11794 3768
rect 11850 3712 11855 3768
rect 10317 3710 11855 3712
rect 10317 3707 10383 3710
rect 11789 3707 11855 3710
rect 12249 3768 12315 3773
rect 12709 3772 12775 3773
rect 12709 3770 12756 3772
rect 12249 3712 12254 3768
rect 12310 3712 12315 3768
rect 12249 3707 12315 3712
rect 12664 3768 12756 3770
rect 12664 3712 12714 3768
rect 12664 3710 12756 3712
rect 12709 3708 12756 3710
rect 12820 3708 12826 3772
rect 12985 3770 13051 3773
rect 13721 3770 13787 3773
rect 14273 3772 14339 3773
rect 14222 3770 14228 3772
rect 12985 3768 13787 3770
rect 12985 3712 12990 3768
rect 13046 3712 13726 3768
rect 13782 3712 13787 3768
rect 12985 3710 13787 3712
rect 14182 3710 14228 3770
rect 14292 3768 14339 3772
rect 14334 3712 14339 3768
rect 12709 3707 12775 3708
rect 12985 3707 13051 3710
rect 13721 3707 13787 3710
rect 14222 3708 14228 3710
rect 14292 3708 14339 3712
rect 14273 3707 14339 3708
rect 7189 3634 7255 3637
rect 10501 3634 10567 3637
rect 7189 3632 10567 3634
rect 7189 3576 7194 3632
rect 7250 3576 10506 3632
rect 10562 3576 10567 3632
rect 7189 3574 10567 3576
rect 7189 3571 7255 3574
rect 10501 3571 10567 3574
rect 11513 3634 11579 3637
rect 12252 3634 12312 3707
rect 11513 3632 12312 3634
rect 11513 3576 11518 3632
rect 11574 3576 12312 3632
rect 11513 3574 12312 3576
rect 14089 3634 14155 3637
rect 15193 3634 15259 3637
rect 14089 3632 15259 3634
rect 14089 3576 14094 3632
rect 14150 3576 15198 3632
rect 15254 3576 15259 3632
rect 14089 3574 15259 3576
rect 11513 3571 11579 3574
rect 14089 3571 14155 3574
rect 15193 3571 15259 3574
rect 0 3498 480 3528
rect 3417 3498 3483 3501
rect 0 3496 3483 3498
rect 0 3440 3422 3496
rect 3478 3440 3483 3496
rect 0 3438 3483 3440
rect 0 3408 480 3438
rect 3417 3435 3483 3438
rect 4061 3498 4127 3501
rect 6177 3498 6243 3501
rect 14365 3498 14431 3501
rect 4061 3496 4906 3498
rect 4061 3440 4066 3496
rect 4122 3440 4906 3496
rect 4061 3438 4906 3440
rect 4061 3435 4127 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 2957 3226 3023 3229
rect 4153 3226 4219 3229
rect 2957 3224 4219 3226
rect 2957 3168 2962 3224
rect 3018 3168 4158 3224
rect 4214 3168 4219 3224
rect 2957 3166 4219 3168
rect 4846 3226 4906 3438
rect 6177 3496 14431 3498
rect 6177 3440 6182 3496
rect 6238 3440 14370 3496
rect 14426 3440 14431 3496
rect 6177 3438 14431 3440
rect 6177 3435 6243 3438
rect 14365 3435 14431 3438
rect 5165 3362 5231 3365
rect 8293 3362 8359 3365
rect 5165 3360 8359 3362
rect 5165 3304 5170 3360
rect 5226 3304 8298 3360
rect 8354 3304 8359 3360
rect 5165 3302 8359 3304
rect 5165 3299 5231 3302
rect 8293 3299 8359 3302
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 5901 3226 5967 3229
rect 10961 3226 11027 3229
rect 4846 3224 11027 3226
rect 4846 3168 5906 3224
rect 5962 3168 10966 3224
rect 11022 3168 11027 3224
rect 4846 3166 11027 3168
rect 2957 3163 3023 3166
rect 4153 3163 4219 3166
rect 5901 3163 5967 3166
rect 10961 3163 11027 3166
rect 11789 3226 11855 3229
rect 17358 3226 17418 3846
rect 22320 3816 22800 3846
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 11789 3224 17418 3226
rect 11789 3168 11794 3224
rect 11850 3168 17418 3224
rect 11789 3166 17418 3168
rect 11789 3163 11855 3166
rect 0 3090 480 3120
rect 2221 3090 2287 3093
rect 0 3088 2287 3090
rect 0 3032 2226 3088
rect 2282 3032 2287 3088
rect 0 3030 2287 3032
rect 0 3000 480 3030
rect 2221 3027 2287 3030
rect 2589 3090 2655 3093
rect 14641 3090 14707 3093
rect 2589 3088 14707 3090
rect 2589 3032 2594 3088
rect 2650 3032 14646 3088
rect 14702 3032 14707 3088
rect 2589 3030 14707 3032
rect 2589 3027 2655 3030
rect 14641 3027 14707 3030
rect 6637 2954 6703 2957
rect 12985 2954 13051 2957
rect 6637 2952 13051 2954
rect 6637 2896 6642 2952
rect 6698 2896 12990 2952
rect 13046 2896 13051 2952
rect 6637 2894 13051 2896
rect 6637 2891 6703 2894
rect 12985 2891 13051 2894
rect 13854 2892 13860 2956
rect 13924 2954 13930 2956
rect 13997 2954 14063 2957
rect 15377 2954 15443 2957
rect 13924 2952 14063 2954
rect 13924 2896 14002 2952
rect 14058 2896 14063 2952
rect 13924 2894 14063 2896
rect 13924 2892 13930 2894
rect 13997 2891 14063 2894
rect 14414 2952 15443 2954
rect 14414 2896 15382 2952
rect 15438 2896 15443 2952
rect 14414 2894 15443 2896
rect 5625 2818 5691 2821
rect 7281 2818 7347 2821
rect 10961 2818 11027 2821
rect 12617 2818 12683 2821
rect 14414 2818 14474 2894
rect 15377 2891 15443 2894
rect 5625 2816 7347 2818
rect 5625 2760 5630 2816
rect 5686 2760 7286 2816
rect 7342 2760 7347 2816
rect 5625 2758 7347 2760
rect 5625 2755 5691 2758
rect 7281 2755 7347 2758
rect 8342 2758 10426 2818
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 5073 2682 5139 2685
rect 5809 2682 5875 2685
rect 3926 2680 5875 2682
rect 3926 2624 5078 2680
rect 5134 2624 5814 2680
rect 5870 2624 5875 2680
rect 3926 2622 5875 2624
rect 0 2546 480 2576
rect 2129 2546 2195 2549
rect 3693 2546 3759 2549
rect 0 2544 3759 2546
rect 0 2488 2134 2544
rect 2190 2488 3698 2544
rect 3754 2488 3759 2544
rect 0 2486 3759 2488
rect 0 2456 480 2486
rect 2129 2483 2195 2486
rect 3693 2483 3759 2486
rect 0 2138 480 2168
rect 3926 2138 3986 2622
rect 5073 2619 5139 2622
rect 5809 2619 5875 2622
rect 7281 2546 7347 2549
rect 8342 2546 8402 2758
rect 10366 2682 10426 2758
rect 10961 2816 12683 2818
rect 10961 2760 10966 2816
rect 11022 2760 12622 2816
rect 12678 2760 12683 2816
rect 10961 2758 12683 2760
rect 10961 2755 11027 2758
rect 12617 2755 12683 2758
rect 12758 2758 14474 2818
rect 12758 2682 12818 2758
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 10366 2622 12818 2682
rect 7281 2544 8402 2546
rect 7281 2488 7286 2544
rect 7342 2488 8402 2544
rect 7281 2486 8402 2488
rect 10133 2546 10199 2549
rect 12065 2546 12131 2549
rect 10133 2544 12131 2546
rect 10133 2488 10138 2544
rect 10194 2488 12070 2544
rect 12126 2488 12131 2544
rect 10133 2486 12131 2488
rect 7281 2483 7347 2486
rect 10133 2483 10199 2486
rect 12065 2483 12131 2486
rect 12985 2546 13051 2549
rect 16113 2546 16179 2549
rect 12985 2544 16179 2546
rect 12985 2488 12990 2544
rect 13046 2488 16118 2544
rect 16174 2488 16179 2544
rect 12985 2486 16179 2488
rect 12985 2483 13051 2486
rect 16113 2483 16179 2486
rect 10317 2410 10383 2413
rect 15193 2410 15259 2413
rect 10317 2408 15259 2410
rect 10317 2352 10322 2408
rect 10378 2352 15198 2408
rect 15254 2352 15259 2408
rect 10317 2350 15259 2352
rect 10317 2347 10383 2350
rect 15193 2347 15259 2350
rect 10869 2276 10935 2277
rect 10869 2274 10916 2276
rect 10824 2272 10916 2274
rect 10824 2216 10874 2272
rect 10824 2214 10916 2216
rect 10869 2212 10916 2214
rect 10980 2212 10986 2276
rect 10869 2211 10935 2212
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2078 3986 2138
rect 0 2048 480 2078
rect 0 1594 480 1624
rect 1945 1594 2011 1597
rect 4153 1594 4219 1597
rect 0 1592 4219 1594
rect 0 1536 1950 1592
rect 2006 1536 4158 1592
rect 4214 1536 4219 1592
rect 0 1534 4219 1536
rect 0 1504 480 1534
rect 1945 1531 2011 1534
rect 4153 1531 4219 1534
rect 0 1186 480 1216
rect 3969 1186 4035 1189
rect 0 1184 4035 1186
rect 0 1128 3974 1184
rect 4030 1128 4035 1184
rect 0 1126 4035 1128
rect 0 1096 480 1126
rect 3969 1123 4035 1126
rect 0 642 480 672
rect 3325 642 3391 645
rect 0 640 3391 642
rect 0 584 3330 640
rect 3386 584 3391 640
rect 0 582 3391 584
rect 0 552 480 582
rect 3325 579 3391 582
rect 0 234 480 264
rect 4061 234 4127 237
rect 0 232 4127 234
rect 0 176 4066 232
rect 4122 176 4127 232
rect 0 174 4127 176
rect 0 144 480 174
rect 4061 171 4127 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 5028 12548 5092 12612
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 12756 9148 12820 9212
rect 4844 8876 4908 8940
rect 5028 8740 5092 8804
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 14228 8604 14292 8668
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 10916 8060 10980 8124
rect 13860 7924 13924 7988
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 12204 6156 12268 6220
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 4844 4252 4908 4316
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 12204 3980 12268 4044
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 12756 3768 12820 3772
rect 12756 3712 12770 3768
rect 12770 3712 12820 3768
rect 12756 3708 12820 3712
rect 14228 3768 14292 3772
rect 14228 3712 14278 3768
rect 14278 3712 14292 3768
rect 14228 3708 14292 3712
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 13860 2892 13924 2956
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 10916 2272 10980 2276
rect 10916 2216 10930 2272
rect 10930 2216 10980 2272
rect 10916 2212 10980 2216
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 5027 12612 5093 12613
rect 5027 12548 5028 12612
rect 5092 12548 5093 12612
rect 5027 12547 5093 12548
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4843 8940 4909 8941
rect 4843 8876 4844 8940
rect 4908 8876 4909 8940
rect 4843 8875 4909 8876
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4846 4317 4906 8875
rect 5030 8805 5090 12547
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 5027 8804 5093 8805
rect 5027 8740 5028 8804
rect 5092 8740 5093 8804
rect 5027 8739 5093 8740
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 12755 9212 12821 9213
rect 12755 9148 12756 9212
rect 12820 9148 12821 9212
rect 12755 9147 12821 9148
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 10915 8124 10981 8125
rect 10915 8060 10916 8124
rect 10980 8060 10981 8124
rect 10915 8059 10981 8060
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 4843 4316 4909 4317
rect 4843 4252 4844 4316
rect 4908 4252 4909 4316
rect 4843 4251 4909 4252
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 10918 2277 10978 8059
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 12203 6220 12269 6221
rect 12203 6156 12204 6220
rect 12268 6156 12269 6220
rect 12203 6155 12269 6156
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 12206 4045 12266 6155
rect 12203 4044 12269 4045
rect 12203 3980 12204 4044
rect 12268 3980 12269 4044
rect 12203 3979 12269 3980
rect 12758 3773 12818 9147
rect 14227 8668 14293 8669
rect 14227 8604 14228 8668
rect 14292 8604 14293 8668
rect 14227 8603 14293 8604
rect 13859 7988 13925 7989
rect 13859 7924 13860 7988
rect 13924 7924 13925 7988
rect 13859 7923 13925 7924
rect 12755 3772 12821 3773
rect 12755 3708 12756 3772
rect 12820 3708 12821 3772
rect 12755 3707 12821 3708
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 10915 2276 10981 2277
rect 10915 2212 10916 2276
rect 10980 2212 10981 2276
rect 10915 2211 10981 2212
rect 11240 2208 11560 3232
rect 13862 2957 13922 7923
rect 14230 3773 14290 8603
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14227 3772 14293 3773
rect 14227 3708 14228 3772
rect 14292 3708 14293 3772
rect 14227 3707 14293 3708
rect 13859 2956 13925 2957
rect 13859 2892 13860 2956
rect 13924 2892 13925 2956
rect 13859 2891 13925 2892
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__decap_6  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1932 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 1932 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_18 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18
timestamp 1605641404
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1605641404
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2944 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_2_
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1605641404
transform 1 0 4692 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1605641404
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41
timestamp 1605641404
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_36
timestamp 1605641404
transform 1 0 4416 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1605641404
transform 1 0 5704 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5060 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5888 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1605641404
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_48
timestamp 1605641404
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1605641404
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 8280 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_4_
timestamp 1605641404
transform 1 0 7084 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 7268 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 8648 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74
timestamp 1605641404
transform 1 0 7912 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 7176 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_76
timestamp 1605641404
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 9936 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1605641404
transform 1 0 10488 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1605641404
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1605641404
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_94
timestamp 1605641404
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_100
timestamp 1605641404
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_111
timestamp 1605641404
transform 1 0 11316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1605641404
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10764 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11592 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1605641404
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1605641404
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11776 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13616 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1605641404
transform 1 0 13432 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1605641404
transform 1 0 14444 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1605641404
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1605641404
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1605641404
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_143
timestamp 1605641404
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1605641404
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1605641404
transform 1 0 14628 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1605641404
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1605641404
transform 1 0 15456 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_160
timestamp 1605641404
transform 1 0 15824 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1605641404
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_160
timestamp 1605641404
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1605641404
transform 1 0 16008 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1605641404
transform 1 0 16376 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_176
timestamp 1605641404
transform 1 0 17296 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_170
timestamp 1605641404
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_172
timestamp 1605641404
transform 1 0 16928 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1605641404
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1605641404
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_184
timestamp 1605641404
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1605641404
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1605641404
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1605641404
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1605641404
transform 1 0 18400 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1605641404
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_192
timestamp 1605641404
transform 1 0 18768 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_204
timestamp 1605641404
transform 1 0 19872 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1605641404
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1605641404
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_216
timestamp 1605641404
transform 1 0 20976 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 1932 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_3_
timestamp 1605641404
transform 1 0 2944 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_18
timestamp 1605641404
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4140 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1605641404
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_32
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1605641404
transform 1 0 5980 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_49
timestamp 1605641404
transform 1 0 5612 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_62
timestamp 1605641404
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6992 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_2_80
timestamp 1605641404
transform 1 0 8464 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1605641404
transform 1 0 9016 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 9844 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1605641404
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11500 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_111
timestamp 1605641404
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13156 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1605641404
transform 1 0 14168 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1605641404
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_140
timestamp 1605641404
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1605641404
transform 1 0 16008 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1605641404
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_160
timestamp 1605641404
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_166
timestamp 1605641404
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1605641404
transform 1 0 16560 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1605641404
transform 1 0 17112 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_172
timestamp 1605641404
transform 1 0 16928 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1605641404
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1605641404
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1605641404
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1605641404
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1605641404
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 1748 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4600 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 3588 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_23
timestamp 1605641404
transform 1 0 3220 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_36
timestamp 1605641404
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6256 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1605641404
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1605641404
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1605641404
transform 1 0 7820 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1605641404
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_82
timestamp 1605641404
transform 1 0 8648 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1605641404
transform 1 0 10396 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1605641404
transform 1 0 9384 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_99
timestamp 1605641404
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11592 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_110
timestamp 1605641404
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1605641404
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1605641404
transform 1 0 14168 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_132
timestamp 1605641404
transform 1 0 13248 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1605641404
transform 1 0 16192 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15180 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_151
timestamp 1605641404
transform 1 0 14996 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_162
timestamp 1605641404
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1605641404
transform 1 0 16744 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_168
timestamp 1605641404
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_174
timestamp 1605641404
transform 1 0 17112 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1605641404
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1605641404
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1605641404
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1605641404
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1564 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1605641404
transform 1 0 3404 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1605641404
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_21
timestamp 1605641404
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1605641404
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_41
timestamp 1605641404
transform 1 0 4876 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6532 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 5520 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_47
timestamp 1605641404
transform 1 0 5428 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_57
timestamp 1605641404
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7544 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_5_
timestamp 1605641404
transform 1 0 8556 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_68
timestamp 1605641404
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_79
timestamp 1605641404
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1605641404
transform 1 0 9752 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10212 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1605641404
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_97
timestamp 1605641404
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12512 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11224 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_108
timestamp 1605641404
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_119
timestamp 1605641404
transform 1 0 12052 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_123
timestamp 1605641404
transform 1 0 12420 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13984 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1605641404
transform 1 0 16284 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1605641404
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1605641404
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1605641404
transform 1 0 17940 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_174
timestamp 1605641404
transform 1 0 17112 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_182
timestamp 1605641404
transform 1 0 17848 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_187
timestamp 1605641404
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_199
timestamp 1605641404
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_211
timestamp 1605641404
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1605641404
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1605641404
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2852 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1605641404
transform 1 0 1840 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1605641404
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_17
timestamp 1605641404
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4784 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_5_28
timestamp 1605641404
transform 1 0 3680 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_56
timestamp 1605641404
transform 1 0 6256 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1605641404
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1605641404
transform 1 0 8280 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_71
timestamp 1605641404
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_77
timestamp 1605641404
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1605641404
transform 1 0 10028 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_87
timestamp 1605641404
transform 1 0 9108 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_95
timestamp 1605641404
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1605641404
transform 1 0 11316 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_106
timestamp 1605641404
transform 1 0 10856 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_110
timestamp 1605641404
transform 1 0 11224 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1605641404
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1605641404
transform 1 0 13892 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14260 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15824 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1605641404
transform 1 0 14812 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_158
timestamp 1605641404
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1605641404
transform 1 0 16836 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1605641404
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_180
timestamp 1605641404
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1605641404
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1605641404
transform 1 0 19780 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_196
timestamp 1605641404
transform 1 0 19136 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_202
timestamp 1605641404
transform 1 0 19688 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_207
timestamp 1605641404
transform 1 0 20148 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1605641404
transform 1 0 21252 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 1748 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1605641404
transform 1 0 2300 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1605641404
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_28
timestamp 1605641404
transform 1 0 3680 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_23
timestamp 1605641404
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_30
timestamp 1605641404
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_22
timestamp 1605641404
transform 1 0 3128 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1605641404
transform 1 0 3404 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_34
timestamp 1605641404
transform 1 0 4232 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_41
timestamp 1605641404
transform 1 0 4876 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4324 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5428 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1605641404
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1605641404
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 7544 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7084 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_63
timestamp 1605641404
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_81
timestamp 1605641404
transform 1 0 8556 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9200 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1605641404
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_102
timestamp 1605641404
transform 1 0 10488 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_86
timestamp 1605641404
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_104
timestamp 1605641404
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 11224 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1605641404
transform 1 0 10856 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_115
timestamp 1605641404
transform 1 0 11684 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1605641404
transform 1 0 14076 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1605641404
transform 1 0 12880 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13524 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_126
timestamp 1605641404
transform 1 0 12696 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_132
timestamp 1605641404
transform 1 0 13248 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_139
timestamp 1605641404
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_144
timestamp 1605641404
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 14536 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1605641404
transform 1 0 16192 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1605641404
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_162
timestamp 1605641404
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17112 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_170
timestamp 1605641404
transform 1 0 16744 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_180
timestamp 1605641404
transform 1 0 17664 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_173
timestamp 1605641404
transform 1 0 17020 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1605641404
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1605641404
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18952 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_192
timestamp 1605641404
transform 1 0 18768 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_200
timestamp 1605641404
transform 1 0 19504 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1605641404
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1605641404
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1605641404
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1605641404
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1605641404
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1932 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_25
timestamp 1605641404
transform 1 0 3404 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp 1605641404
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1605641404
transform 1 0 5152 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5888 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_47
timestamp 1605641404
transform 1 0 5428 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_51
timestamp 1605641404
transform 1 0 5796 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1605641404
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_68
timestamp 1605641404
transform 1 0 7360 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_74
timestamp 1605641404
transform 1 0 7912 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1605641404
transform 1 0 9016 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1605641404
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1605641404
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12420 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1605641404
transform 1 0 11408 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_109
timestamp 1605641404
transform 1 0 11132 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_121
timestamp 1605641404
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1605641404
transform 1 0 13432 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_132
timestamp 1605641404
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_143
timestamp 1605641404
transform 1 0 14260 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1605641404
transform 1 0 14720 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_147
timestamp 1605641404
transform 1 0 14628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1605641404
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_163
timestamp 1605641404
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_175
timestamp 1605641404
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_187
timestamp 1605641404
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_199
timestamp 1605641404
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_211
timestamp 1605641404
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1605641404
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1605641404
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 1840 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1605641404
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 4692 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 3496 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_24
timestamp 1605641404
transform 1 0 3312 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_35
timestamp 1605641404
transform 1 0 4324 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1605641404
transform 1 0 6348 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_55
timestamp 1605641404
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1605641404
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1605641404
transform 1 0 7820 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1605641404
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1605641404
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1605641404
transform 1 0 9752 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_103
timestamp 1605641404
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1605641404
transform 1 0 11868 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1605641404
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_114
timestamp 1605641404
transform 1 0 11592 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1605641404
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14444 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1605641404
transform 1 0 13432 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1605641404
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_143
timestamp 1605641404
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1605641404
transform 1 0 15456 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_154
timestamp 1605641404
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_165
timestamp 1605641404
transform 1 0 16284 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_177
timestamp 1605641404
transform 1 0 17388 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1605641404
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1605641404
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1605641404
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_19
timestamp 1605641404
transform 1 0 2852 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1605641404
transform 1 0 3036 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_24
timestamp 1605641404
transform 1 0 3312 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1605641404
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_41
timestamp 1605641404
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1605641404
transform 1 0 6164 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1605641404
transform 1 0 5152 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_53
timestamp 1605641404
transform 1 0 5980 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1605641404
transform 1 0 8740 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7728 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_64
timestamp 1605641404
transform 1 0 6992 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_81
timestamp 1605641404
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_86
timestamp 1605641404
transform 1 0 9016 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 11408 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_10_109
timestamp 1605641404
transform 1 0 11132 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13064 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_128
timestamp 1605641404
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_146
timestamp 1605641404
transform 1 0 14536 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1605641404
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1605641404
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1605641404
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1605641404
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1605641404
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1605641404
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1605641404
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 2208 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1472 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_10
timestamp 1605641404
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 3864 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_28
timestamp 1605641404
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_39
timestamp 1605641404
transform 1 0 4692 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5060 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1605641404
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6992 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 8648 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1605641404
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10672 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1605641404
transform 1 0 10396 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_98
timestamp 1605641404
transform 1 0 10120 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1605641404
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1605641404
transform 1 0 13432 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14444 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_132
timestamp 1605641404
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_143
timestamp 1605641404
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_154
timestamp 1605641404
transform 1 0 15272 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_166
timestamp 1605641404
transform 1 0 16376 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1605641404
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1605641404
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1605641404
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1605641404
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1605641404
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1605641404
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1605641404
transform 1 0 1840 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2852 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1605641404
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_17
timestamp 1605641404
transform 1 0 2668 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_28
timestamp 1605641404
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1605641404
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1605641404
transform 1 0 6072 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1605641404
transform 1 0 5060 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1605641404
transform 1 0 6716 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_52
timestamp 1605641404
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_57
timestamp 1605641404
transform 1 0 6348 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7912 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1605641404
transform 1 0 7728 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_70
timestamp 1605641404
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_83
timestamp 1605641404
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1605641404
transform 1 0 10120 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1605641404
transform 1 0 10580 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1605641404
transform 1 0 8924 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1605641404
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1605641404
transform 1 0 10028 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_101
timestamp 1605641404
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_3_
timestamp 1605641404
transform 1 0 11684 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_112
timestamp 1605641404
transform 1 0 11408 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_124
timestamp 1605641404
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13708 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_3_
timestamp 1605641404
transform 1 0 12696 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_135
timestamp 1605641404
transform 1 0 13524 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1605641404
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1605641404
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1605641404
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1605641404
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1605641404
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1605641404
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1605641404
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1605641404
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1605641404
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2760 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 1748 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 1748 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1605641404
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1605641404
transform 1 0 3404 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4876 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1605641404
transform 1 0 4600 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1605641404
transform 1 0 4600 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_34
timestamp 1605641404
transform 1 0 4232 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1605641404
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_28
timestamp 1605641404
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_32
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5796 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1605641404
transform 1 0 6348 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_47
timestamp 1605641404
transform 1 0 5428 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7452 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7820 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1605641404
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_82
timestamp 1605641404
transform 1 0 8648 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_67
timestamp 1605641404
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_6_
timestamp 1605641404
transform 1 0 9660 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10488 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_90
timestamp 1605641404
transform 1 0 9384 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1605641404
transform 1 0 8924 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1605641404
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 11316 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1605641404
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_109
timestamp 1605641404
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12972 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1605641404
transform 1 0 14444 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1605641404
transform 1 0 13432 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1605641404
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1605641404
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_127
timestamp 1605641404
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1605641404
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_154
timestamp 1605641404
transform 1 0 15272 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_166
timestamp 1605641404
transform 1 0 16376 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1605641404
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1605641404
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1605641404
transform 1 0 17480 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1605641404
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1605641404
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1605641404
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1605641404
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1605641404
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1605641404
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1605641404
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1605641404
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1605641404
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1605641404
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1605641404
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1605641404
transform 1 0 4048 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 3036 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1605641404
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_41
timestamp 1605641404
transform 1 0 4876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1605641404
transform 1 0 6072 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1605641404
transform 1 0 5060 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_52
timestamp 1605641404
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1605641404
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7820 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1605641404
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1605641404
transform 1 0 9384 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9660 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_89
timestamp 1605641404
transform 1 0 9292 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11132 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 12604 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1605641404
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1605641404
transform 1 0 14168 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1605641404
transform 1 0 13156 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_128
timestamp 1605641404
transform 1 0 12880 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_140
timestamp 1605641404
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_151
timestamp 1605641404
transform 1 0 14996 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_163
timestamp 1605641404
transform 1 0 16100 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1605641404
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_175
timestamp 1605641404
transform 1 0 17204 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1605641404
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1605641404
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1605641404
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 2300 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1564 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1605641404
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1605641404
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1605641404
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1605641404
transform 1 0 5060 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_3_
timestamp 1605641404
transform 1 0 6072 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_52
timestamp 1605641404
transform 1 0 5888 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_1_
timestamp 1605641404
transform 1 0 7360 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1605641404
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1605641404
transform 1 0 7084 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_63
timestamp 1605641404
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_77
timestamp 1605641404
transform 1 0 8188 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10304 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1605641404
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_93
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_99
timestamp 1605641404
transform 1 0 10212 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12144 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12972 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1605641404
transform 1 0 13800 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1605641404
transform 1 0 14628 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1605641404
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1605641404
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1605641404
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_190
timestamp 1605641404
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1605641404
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1605641404
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1605641404
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1605641404
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2944 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 1932 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1605641404
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_18
timestamp 1605641404
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4784 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 3956 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_29
timestamp 1605641404
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_37
timestamp 1605641404
transform 1 0 4508 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_56
timestamp 1605641404
transform 1 0 6256 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1605641404
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 8464 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_78
timestamp 1605641404
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_83
timestamp 1605641404
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1605641404
transform 1 0 9936 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10580 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1605641404
transform 1 0 8924 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_94
timestamp 1605641404
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_99
timestamp 1605641404
transform 1 0 10212 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_119
timestamp 1605641404
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_123
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12972 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_145
timestamp 1605641404
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1605641404
transform 1 0 14628 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_156
timestamp 1605641404
transform 1 0 15456 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1605641404
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_168
timestamp 1605641404
transform 1 0 16560 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1605641404
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1605641404
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1605641404
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1605641404
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1605641404
transform 1 0 1472 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1605641404
transform 1 0 2484 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_13
timestamp 1605641404
transform 1 0 2300 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1605641404
transform 1 0 3496 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4416 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_24
timestamp 1605641404
transform 1 0 3312 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1605641404
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6072 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1605641404
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1605641404
transform 1 0 8556 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7176 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_63
timestamp 1605641404
transform 1 0 6900 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_75
timestamp 1605641404
transform 1 0 8004 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1605641404
transform 1 0 9936 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1605641404
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_93
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_1_
timestamp 1605641404
transform 1 0 11960 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l3_in_0_
timestamp 1605641404
transform 1 0 10948 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_105
timestamp 1605641404
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_116
timestamp 1605641404
transform 1 0 11776 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13524 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_127
timestamp 1605641404
transform 1 0 12788 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1605641404
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_163
timestamp 1605641404
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_175
timestamp 1605641404
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_187
timestamp 1605641404
transform 1 0 18308 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_199
timestamp 1605641404
transform 1 0 19412 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1605641404
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_211
timestamp 1605641404
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1605641404
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1605641404
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp 1605641404
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1605641404
transform 1 0 1932 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1605641404
transform 1 0 1564 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_18
timestamp 1605641404
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 2392 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4600 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1605641404
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp 1605641404
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1605641404
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1605641404
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_41
timestamp 1605641404
transform 1 0 4876 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6164 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5152 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5612 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_47
timestamp 1605641404
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_58
timestamp 1605641404
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_53
timestamp 1605641404
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7360 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 7912 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_19_66
timestamp 1605641404
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_71
timestamp 1605641404
transform 1 0 7636 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 10672 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1605641404
transform 1 0 9016 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_84
timestamp 1605641404
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_95
timestamp 1605641404
transform 1 0 9844 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_103
timestamp 1605641404
transform 1 0 10580 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1605641404
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12052 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11316 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1605641404
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_109
timestamp 1605641404
transform 1 0 11132 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_117
timestamp 1605641404
transform 1 0 11868 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 13248 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1605641404
transform 1 0 13708 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 12880 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_126
timestamp 1605641404
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_131
timestamp 1605641404
transform 1 0 13156 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_135
timestamp 1605641404
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_148
timestamp 1605641404
transform 1 0 14720 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_160
timestamp 1605641404
transform 1 0 15824 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_146
timestamp 1605641404
transform 1 0 14536 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1605641404
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1605641404
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17020 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1605641404
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_172
timestamp 1605641404
transform 1 0 16928 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1605641404
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1605641404
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1605641404
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 19136 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1605641404
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1605641404
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1605641404
transform 1 0 18584 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1605641404
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1605641404
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1605641404
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1605641404
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 2392 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_12
timestamp 1605641404
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4416 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_21_30
timestamp 1605641404
transform 1 0 3864 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1605641404
transform 1 0 6072 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_52
timestamp 1605641404
transform 1 0 5888 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1605641404
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_62
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8740 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 7728 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1605641404
transform 1 0 7084 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_68
timestamp 1605641404
transform 1 0 7360 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_81
timestamp 1605641404
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1605641404
transform 1 0 9844 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_92
timestamp 1605641404
transform 1 0 9568 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_104
timestamp 1605641404
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12512 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_6_
timestamp 1605641404
transform 1 0 10856 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_115
timestamp 1605641404
transform 1 0 11684 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1605641404
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_123
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13524 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_133
timestamp 1605641404
transform 1 0 13340 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_144
timestamp 1605641404
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_5_
timestamp 1605641404
transform 1 0 14536 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_155
timestamp 1605641404
transform 1 0 15364 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1605641404
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_167
timestamp 1605641404
transform 1 0 16468 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1605641404
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1605641404
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1605641404
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1605641404
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 1932 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1605641404
transform 1 0 2944 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1605641404
transform 1 0 1748 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_18
timestamp 1605641404
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4508 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1605641404
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_32
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_36
timestamp 1605641404
transform 1 0 4416 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1605641404
transform 1 0 6164 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 6624 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_53
timestamp 1605641404
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_58
timestamp 1605641404
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 7636 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_69
timestamp 1605641404
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_80
timestamp 1605641404
transform 1 0 8464 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1605641404
transform 1 0 9108 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1605641404
transform 1 0 9936 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1605641404
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_86
timestamp 1605641404
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1605641404
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11316 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1605641404
transform 1 0 10948 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1605641404
transform 1 0 12604 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_105
timestamp 1605641404
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_110
timestamp 1605641404
transform 1 0 11224 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_120
timestamp 1605641404
transform 1 0 12144 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_124
timestamp 1605641404
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12880 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_144
timestamp 1605641404
transform 1 0 14352 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_4_
timestamp 1605641404
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1605641404
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1605641404
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_163
timestamp 1605641404
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_175
timestamp 1605641404
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_187
timestamp 1605641404
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_199
timestamp 1605641404
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1605641404
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1605641404
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1605641404
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1605641404
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1605641404
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2944 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 1932 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1605641404
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1605641404
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_18
timestamp 1605641404
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1605641404
transform 1 0 4692 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_23_36
timestamp 1605641404
transform 1 0 4416 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1605641404
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_48
timestamp 1605641404
transform 1 0 5520 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1605641404
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1605641404
transform 1 0 8556 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_23_78
timestamp 1605641404
transform 1 0 8280 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10580 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1605641404
transform 1 0 9568 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_90
timestamp 1605641404
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1605641404
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12420 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1605641404
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_119
timestamp 1605641404
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14076 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_139
timestamp 1605641404
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_150
timestamp 1605641404
transform 1 0 14904 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_162
timestamp 1605641404
transform 1 0 16008 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1605641404
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_174
timestamp 1605641404
transform 1 0 17112 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1605641404
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1605641404
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1605641404
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1605641404
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1605641404
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1605641404
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1605641404
transform 1 0 2944 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 1932 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1605641404
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1605641404
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_18
timestamp 1605641404
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_1_
timestamp 1605641404
transform 1 0 4784 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1605641404
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1605641404
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_38
timestamp 1605641404
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5796 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_49
timestamp 1605641404
transform 1 0 5612 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_60
timestamp 1605641404
transform 1 0 6624 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7912 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6900 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_72
timestamp 1605641404
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 9660 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1605641404
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1605641404
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12328 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11316 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_109
timestamp 1605641404
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_120
timestamp 1605641404
transform 1 0 12144 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13984 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1605641404
transform 1 0 13800 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1605641404
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1605641404
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1605641404
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1605641404
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1605641404
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1605641404
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1605641404
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1605641404
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1605641404
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1605641404
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1605641404
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1605641404
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 2576 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1840 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1605641404
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_6
timestamp 1605641404
transform 1 0 1656 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_14
timestamp 1605641404
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4232 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_32
timestamp 1605641404
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1605641404
transform 1 0 5888 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_1_
timestamp 1605641404
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1605641404
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1605641404
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_50
timestamp 1605641404
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_56
timestamp 1605641404
transform 1 0 6256 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1605641404
transform 1 0 7820 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1605641404
transform 1 0 8280 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8740 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_71
timestamp 1605641404
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_76
timestamp 1605641404
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_81
timestamp 1605641404
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10580 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_92
timestamp 1605641404
transform 1 0 9568 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_100
timestamp 1605641404
transform 1 0 10304 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12420 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11592 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1605641404
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_112
timestamp 1605641404
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1605641404
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1605641404
transform 1 0 14076 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1605641404
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_144
timestamp 1605641404
transform 1 0 14352 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_156
timestamp 1605641404
transform 1 0 15456 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1605641404
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_168
timestamp 1605641404
transform 1 0 16560 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1605641404
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1605641404
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1605641404
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1605641404
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1605641404
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1605641404
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_8
timestamp 1605641404
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1605641404
transform 1 0 1380 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1605641404
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1605641404
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1472 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1605641404
transform 1 0 1472 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_18
timestamp 1605641404
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_10
timestamp 1605641404
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_16
timestamp 1605641404
transform 1 0 2576 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2024 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2208 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2944 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4048 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4692 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1605641404
transform 1 0 3680 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1605641404
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1605641404
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_26
timestamp 1605641404
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_37
timestamp 1605641404
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5704 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6808 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1605641404
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_48
timestamp 1605641404
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_48
timestamp 1605641404
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1605641404
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8464 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8372 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7360 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_66
timestamp 1605641404
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_77
timestamp 1605641404
transform 1 0 8188 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_78
timestamp 1605641404
transform 1 0 8280 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10120 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_1_
timestamp 1605641404
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1605641404
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1605641404
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_102
timestamp 1605641404
transform 1 0 10488 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_96
timestamp 1605641404
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1605641404
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1605641404
transform 1 0 11776 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11868 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1605641404
transform 1 0 10856 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1605641404
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_115
timestamp 1605641404
transform 1 0 11684 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1605641404
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_119
timestamp 1605641404
transform 1 0 12052 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1605641404
transform 1 0 13432 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12880 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_126
timestamp 1605641404
transform 1 0 12696 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_134
timestamp 1605641404
transform 1 0 13432 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_126
timestamp 1605641404
transform 1 0 12696 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_138
timestamp 1605641404
transform 1 0 13800 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1605641404
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_146
timestamp 1605641404
transform 1 0 14536 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1605641404
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1605641404
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1605641404
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_150
timestamp 1605641404
transform 1 0 14904 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_162
timestamp 1605641404
transform 1 0 16008 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1605641404
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1605641404
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_174
timestamp 1605641404
transform 1 0 17112 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1605641404
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1605641404
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1605641404
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1605641404
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1605641404
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1605641404
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1605641404
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1605641404
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1605641404
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1605641404
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1605641404
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1605641404
transform 1 0 1472 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2760 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2024 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1605641404
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1605641404
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_8
timestamp 1605641404
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_16
timestamp 1605641404
transform 1 0 2576 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1605641404
transform 1 0 3496 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1605641404
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4784 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1605641404
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_24
timestamp 1605641404
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1605641404
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_36
timestamp 1605641404
transform 1 0 4416 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1605641404
transform 1 0 6072 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_49
timestamp 1605641404
transform 1 0 5612 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_53
timestamp 1605641404
transform 1 0 5980 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1605641404
transform 1 0 8740 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7084 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_63
timestamp 1605641404
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_81
timestamp 1605641404
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1605641404
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10580 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1605641404
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_87
timestamp 1605641404
transform 1 0 9108 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1605641404
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_97
timestamp 1605641404
transform 1 0 10028 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12236 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_119
timestamp 1605641404
transform 1 0 12052 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1605641404
transform 1 0 13248 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_130
timestamp 1605641404
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_136
timestamp 1605641404
transform 1 0 13616 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_144
timestamp 1605641404
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1605641404
transform 1 0 14536 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1605641404
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_150
timestamp 1605641404
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1605641404
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1605641404
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1605641404
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1605641404
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1605641404
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1605641404
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1605641404
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1605641404
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1605641404
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1605641404
transform 1 0 2300 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1605641404
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 2760 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1605641404
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1605641404
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1605641404
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_16
timestamp 1605641404
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4692 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_34
timestamp 1605641404
transform 1 0 4232 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_38
timestamp 1605641404
transform 1 0 4600 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1605641404
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1605641404
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_55
timestamp 1605641404
transform 1 0 6164 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 8464 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1605641404
transform 1 0 7452 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_66
timestamp 1605641404
transform 1 0 7176 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1605641404
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1605641404
transform 1 0 10120 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_96
timestamp 1605641404
transform 1 0 9936 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_102
timestamp 1605641404
transform 1 0 10488 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1605641404
transform 1 0 11776 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12420 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1605641404
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1605641404
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_119
timestamp 1605641404
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13156 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_129
timestamp 1605641404
transform 1 0 12972 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1605641404
transform 1 0 13708 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1605641404
transform 1 0 14812 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_161
timestamp 1605641404
transform 1 0 15916 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1605641404
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_173
timestamp 1605641404
transform 1 0 17020 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1605641404
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1605641404
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1605641404
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1605641404
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1605641404
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1472 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2208 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1605641404
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1605641404
transform 1 0 1380 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_10
timestamp 1605641404
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1605641404
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4048 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1605641404
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1605641404
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5704 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_48
timestamp 1605641404
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7360 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_66
timestamp 1605641404
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1605641404
transform 1 0 9016 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9844 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1605641404
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_84
timestamp 1605641404
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1605641404
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1605641404
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_104
timestamp 1605641404
transform 1 0 10672 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11132 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_30_108
timestamp 1605641404
transform 1 0 11040 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_125
timestamp 1605641404
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12788 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13800 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_136
timestamp 1605641404
transform 1 0 13616 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_144
timestamp 1605641404
transform 1 0 14352 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15272 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1605641404
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1605641404
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_160
timestamp 1605641404
transform 1 0 15824 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_172
timestamp 1605641404
transform 1 0 16928 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_184
timestamp 1605641404
transform 1 0 18032 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18768 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_198
timestamp 1605641404
transform 1 0 19320 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1605641404
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1605641404
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1605641404
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1605641404
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1605641404
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1605641404
transform 1 0 1564 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2852 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2116 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1605641404
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1605641404
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_9
timestamp 1605641404
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_17
timestamp 1605641404
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4140 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_28
timestamp 1605641404
transform 1 0 3680 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_32
timestamp 1605641404
transform 1 0 4048 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1605641404
transform 1 0 5796 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1605641404
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_49
timestamp 1605641404
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_55
timestamp 1605641404
transform 1 0 6164 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_62
timestamp 1605641404
transform 1 0 6808 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1605641404
transform 1 0 7912 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8372 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6900 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_72
timestamp 1605641404
transform 1 0 7728 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_77
timestamp 1605641404
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10028 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_95
timestamp 1605641404
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1605641404
transform 1 0 11684 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1605641404
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1605641404
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1605641404
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1605641404
transform 1 0 14076 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1605641404
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_145
timestamp 1605641404
transform 1 0 14444 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1605641404
transform 1 0 16284 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1605641404
transform 1 0 15732 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1605641404
transform 1 0 15180 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1605641404
transform 1 0 14628 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_151
timestamp 1605641404
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_157
timestamp 1605641404
transform 1 0 15548 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_163
timestamp 1605641404
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1605641404
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1605641404
transform 1 0 17388 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1605641404
transform 1 0 16836 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1605641404
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1605641404
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1605641404
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1605641404
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1605641404
transform 1 0 19688 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1605641404
transform 1 0 19136 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1605641404
transform 1 0 18584 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_188
timestamp 1605641404
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_194
timestamp 1605641404
transform 1 0 18952 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_200
timestamp 1605641404
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_206
timestamp 1605641404
transform 1 0 20056 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1605641404
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_218
timestamp 1605641404
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1605641404
transform 1 0 1656 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2208 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1605641404
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1605641404
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_10
timestamp 1605641404
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_18
timestamp 1605641404
transform 1 0 2760 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4232 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1605641404
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1605641404
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_32
timestamp 1605641404
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1605641404
transform 1 0 6348 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5336 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1605641404
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_43
timestamp 1605641404
transform 1 0 5060 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_55
timestamp 1605641404
transform 1 0 6164 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_60
timestamp 1605641404
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6900 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8648 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_32_79
timestamp 1605641404
transform 1 0 8372 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 10488 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 9752 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1605641404
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_91
timestamp 1605641404
transform 1 0 9476 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_100
timestamp 1605641404
transform 1 0 10304 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1605641404
transform 1 0 11316 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1605641404
transform 1 0 11868 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1605641404
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1605641404
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_108
timestamp 1605641404
transform 1 0 11040 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_115
timestamp 1605641404
transform 1 0 11684 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_121
timestamp 1605641404
transform 1 0 12236 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1605641404
transform 1 0 13708 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1605641404
transform 1 0 13156 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_129
timestamp 1605641404
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_135
timestamp 1605641404
transform 1 0 13524 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1605641404
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1605641404
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_153
timestamp 1605641404
transform 1 0 15180 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_156
timestamp 1605641404
transform 1 0 15456 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_164
timestamp 1605641404
transform 1 0 16192 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1605641404
transform 1 0 16468 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1605641404
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_171
timestamp 1605641404
transform 1 0 16836 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_183
timestamp 1605641404
transform 1 0 17940 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1605641404
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1605641404
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1605641404
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1605641404
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_211
timestamp 1605641404
transform 1 0 20516 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1605641404
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 0 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_43_
port 1 nsew default input
rlabel metal2 s 1122 0 1178 480 6 bottom_left_grid_pin_44_
port 2 nsew default input
rlabel metal2 s 1582 0 1638 480 6 bottom_left_grid_pin_45_
port 3 nsew default input
rlabel metal2 s 2042 0 2098 480 6 bottom_left_grid_pin_46_
port 4 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_47_
port 5 nsew default input
rlabel metal2 s 2962 0 3018 480 6 bottom_left_grid_pin_48_
port 6 nsew default input
rlabel metal2 s 3422 0 3478 480 6 bottom_left_grid_pin_49_
port 7 nsew default input
rlabel metal2 s 22466 0 22522 480 6 bottom_right_grid_pin_1_
port 8 nsew default input
rlabel metal3 s 22320 11432 22800 11552 6 ccff_head
port 9 nsew default input
rlabel metal3 s 22320 19048 22800 19168 6 ccff_tail
port 10 nsew default tristate
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[0]
port 11 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[10]
port 12 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[11]
port 13 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_left_in[12]
port 14 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[13]
port 15 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[14]
port 16 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[15]
port 17 nsew default input
rlabel metal3 s 0 11568 480 11688 6 chanx_left_in[16]
port 18 nsew default input
rlabel metal3 s 0 11976 480 12096 6 chanx_left_in[17]
port 19 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[18]
port 20 nsew default input
rlabel metal3 s 0 12928 480 13048 6 chanx_left_in[19]
port 21 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[1]
port 22 nsew default input
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[2]
port 23 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[3]
port 24 nsew default input
rlabel metal3 s 0 5856 480 5976 6 chanx_left_in[4]
port 25 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[5]
port 26 nsew default input
rlabel metal3 s 0 6808 480 6928 6 chanx_left_in[6]
port 27 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[7]
port 28 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[8]
port 29 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[9]
port 30 nsew default input
rlabel metal3 s 0 13472 480 13592 6 chanx_left_out[0]
port 31 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[10]
port 32 nsew default tristate
rlabel metal3 s 0 18640 480 18760 6 chanx_left_out[11]
port 33 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[12]
port 34 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chanx_left_out[13]
port 35 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[14]
port 36 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[15]
port 37 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[16]
port 38 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[17]
port 39 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[18]
port 40 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[19]
port 41 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[1]
port 42 nsew default tristate
rlabel metal3 s 0 14424 480 14544 6 chanx_left_out[2]
port 43 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 chanx_left_out[3]
port 44 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[4]
port 45 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 chanx_left_out[5]
port 46 nsew default tristate
rlabel metal3 s 0 16328 480 16448 6 chanx_left_out[6]
port 47 nsew default tristate
rlabel metal3 s 0 16736 480 16856 6 chanx_left_out[7]
port 48 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[8]
port 49 nsew default tristate
rlabel metal3 s 0 17688 480 17808 6 chanx_left_out[9]
port 50 nsew default tristate
rlabel metal2 s 3882 0 3938 480 6 chany_bottom_in[0]
port 51 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[10]
port 52 nsew default input
rlabel metal2 s 9034 0 9090 480 6 chany_bottom_in[11]
port 53 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[12]
port 54 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[13]
port 55 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[14]
port 56 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[15]
port 57 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[16]
port 58 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[17]
port 59 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[18]
port 60 nsew default input
rlabel metal2 s 12714 0 12770 480 6 chany_bottom_in[19]
port 61 nsew default input
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_in[1]
port 62 nsew default input
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_in[2]
port 63 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[3]
port 64 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[4]
port 65 nsew default input
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[5]
port 66 nsew default input
rlabel metal2 s 6642 0 6698 480 6 chany_bottom_in[6]
port 67 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[7]
port 68 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[8]
port 69 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_in[9]
port 70 nsew default input
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_out[0]
port 71 nsew default tristate
rlabel metal2 s 17866 0 17922 480 6 chany_bottom_out[10]
port 72 nsew default tristate
rlabel metal2 s 18326 0 18382 480 6 chany_bottom_out[11]
port 73 nsew default tristate
rlabel metal2 s 18786 0 18842 480 6 chany_bottom_out[12]
port 74 nsew default tristate
rlabel metal2 s 19246 0 19302 480 6 chany_bottom_out[13]
port 75 nsew default tristate
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[14]
port 76 nsew default tristate
rlabel metal2 s 20166 0 20222 480 6 chany_bottom_out[15]
port 77 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 chany_bottom_out[16]
port 78 nsew default tristate
rlabel metal2 s 21086 0 21142 480 6 chany_bottom_out[17]
port 79 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[18]
port 80 nsew default tristate
rlabel metal2 s 22006 0 22062 480 6 chany_bottom_out[19]
port 81 nsew default tristate
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_out[1]
port 82 nsew default tristate
rlabel metal2 s 14094 0 14150 480 6 chany_bottom_out[2]
port 83 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[3]
port 84 nsew default tristate
rlabel metal2 s 15014 0 15070 480 6 chany_bottom_out[4]
port 85 nsew default tristate
rlabel metal2 s 15566 0 15622 480 6 chany_bottom_out[5]
port 86 nsew default tristate
rlabel metal2 s 16026 0 16082 480 6 chany_bottom_out[6]
port 87 nsew default tristate
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[7]
port 88 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 chany_bottom_out[8]
port 89 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[9]
port 90 nsew default tristate
rlabel metal2 s 3882 22320 3938 22800 6 chany_top_in[0]
port 91 nsew default input
rlabel metal2 s 8574 22320 8630 22800 6 chany_top_in[10]
port 92 nsew default input
rlabel metal2 s 9034 22320 9090 22800 6 chany_top_in[11]
port 93 nsew default input
rlabel metal2 s 9494 22320 9550 22800 6 chany_top_in[12]
port 94 nsew default input
rlabel metal2 s 9954 22320 10010 22800 6 chany_top_in[13]
port 95 nsew default input
rlabel metal2 s 10414 22320 10470 22800 6 chany_top_in[14]
port 96 nsew default input
rlabel metal2 s 10874 22320 10930 22800 6 chany_top_in[15]
port 97 nsew default input
rlabel metal2 s 11334 22320 11390 22800 6 chany_top_in[16]
port 98 nsew default input
rlabel metal2 s 11794 22320 11850 22800 6 chany_top_in[17]
port 99 nsew default input
rlabel metal2 s 12254 22320 12310 22800 6 chany_top_in[18]
port 100 nsew default input
rlabel metal2 s 12714 22320 12770 22800 6 chany_top_in[19]
port 101 nsew default input
rlabel metal2 s 4342 22320 4398 22800 6 chany_top_in[1]
port 102 nsew default input
rlabel metal2 s 4802 22320 4858 22800 6 chany_top_in[2]
port 103 nsew default input
rlabel metal2 s 5262 22320 5318 22800 6 chany_top_in[3]
port 104 nsew default input
rlabel metal2 s 5722 22320 5778 22800 6 chany_top_in[4]
port 105 nsew default input
rlabel metal2 s 6182 22320 6238 22800 6 chany_top_in[5]
port 106 nsew default input
rlabel metal2 s 6642 22320 6698 22800 6 chany_top_in[6]
port 107 nsew default input
rlabel metal2 s 7102 22320 7158 22800 6 chany_top_in[7]
port 108 nsew default input
rlabel metal2 s 7562 22320 7618 22800 6 chany_top_in[8]
port 109 nsew default input
rlabel metal2 s 8114 22320 8170 22800 6 chany_top_in[9]
port 110 nsew default input
rlabel metal2 s 13174 22320 13230 22800 6 chany_top_out[0]
port 111 nsew default tristate
rlabel metal2 s 17866 22320 17922 22800 6 chany_top_out[10]
port 112 nsew default tristate
rlabel metal2 s 18326 22320 18382 22800 6 chany_top_out[11]
port 113 nsew default tristate
rlabel metal2 s 18786 22320 18842 22800 6 chany_top_out[12]
port 114 nsew default tristate
rlabel metal2 s 19246 22320 19302 22800 6 chany_top_out[13]
port 115 nsew default tristate
rlabel metal2 s 19706 22320 19762 22800 6 chany_top_out[14]
port 116 nsew default tristate
rlabel metal2 s 20166 22320 20222 22800 6 chany_top_out[15]
port 117 nsew default tristate
rlabel metal2 s 20626 22320 20682 22800 6 chany_top_out[16]
port 118 nsew default tristate
rlabel metal2 s 21086 22320 21142 22800 6 chany_top_out[17]
port 119 nsew default tristate
rlabel metal2 s 21546 22320 21602 22800 6 chany_top_out[18]
port 120 nsew default tristate
rlabel metal2 s 22006 22320 22062 22800 6 chany_top_out[19]
port 121 nsew default tristate
rlabel metal2 s 13634 22320 13690 22800 6 chany_top_out[1]
port 122 nsew default tristate
rlabel metal2 s 14094 22320 14150 22800 6 chany_top_out[2]
port 123 nsew default tristate
rlabel metal2 s 14554 22320 14610 22800 6 chany_top_out[3]
port 124 nsew default tristate
rlabel metal2 s 15014 22320 15070 22800 6 chany_top_out[4]
port 125 nsew default tristate
rlabel metal2 s 15566 22320 15622 22800 6 chany_top_out[5]
port 126 nsew default tristate
rlabel metal2 s 16026 22320 16082 22800 6 chany_top_out[6]
port 127 nsew default tristate
rlabel metal2 s 16486 22320 16542 22800 6 chany_top_out[7]
port 128 nsew default tristate
rlabel metal2 s 16946 22320 17002 22800 6 chany_top_out[8]
port 129 nsew default tristate
rlabel metal2 s 17406 22320 17462 22800 6 chany_top_out[9]
port 130 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 131 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_35_
port 132 nsew default input
rlabel metal3 s 0 1096 480 1216 6 left_bottom_grid_pin_36_
port 133 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_37_
port 134 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_38_
port 135 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_39_
port 136 nsew default input
rlabel metal3 s 0 3000 480 3120 6 left_bottom_grid_pin_40_
port 137 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_41_
port 138 nsew default input
rlabel metal3 s 22320 3816 22800 3936 6 prog_clk
port 139 nsew default input
rlabel metal2 s 202 22320 258 22800 6 top_left_grid_pin_42_
port 140 nsew default input
rlabel metal2 s 662 22320 718 22800 6 top_left_grid_pin_43_
port 141 nsew default input
rlabel metal2 s 1122 22320 1178 22800 6 top_left_grid_pin_44_
port 142 nsew default input
rlabel metal2 s 1582 22320 1638 22800 6 top_left_grid_pin_45_
port 143 nsew default input
rlabel metal2 s 2042 22320 2098 22800 6 top_left_grid_pin_46_
port 144 nsew default input
rlabel metal2 s 2502 22320 2558 22800 6 top_left_grid_pin_47_
port 145 nsew default input
rlabel metal2 s 2962 22320 3018 22800 6 top_left_grid_pin_48_
port 146 nsew default input
rlabel metal2 s 3422 22320 3478 22800 6 top_left_grid_pin_49_
port 147 nsew default input
rlabel metal2 s 22466 22320 22522 22800 6 top_right_grid_pin_1_
port 148 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 149 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 150 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
