VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__0_
  CLASS BLOCK ;
  FOREIGN sb_0__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 2.400 ;
    END
  END address[5]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 6.840 140.000 7.440 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 11.600 140.000 12.200 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 17.040 140.000 17.640 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 21.800 140.000 22.400 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 26.560 140.000 27.160 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 32.000 140.000 32.600 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 36.760 140.000 37.360 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 41.520 140.000 42.120 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 46.960 140.000 47.560 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 96.600 140.000 97.200 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 102.040 140.000 102.640 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 106.800 140.000 107.400 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 111.560 140.000 112.160 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 117.000 140.000 117.600 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 121.760 140.000 122.360 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 126.520 140.000 127.120 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 131.960 140.000 132.560 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 136.720 140.000 137.320 ;
    END
  END chanx_right_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 137.600 4.050 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.130 137.600 11.410 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.950 137.600 19.230 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 137.600 27.050 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 137.600 34.870 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.410 137.600 42.690 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 137.600 50.510 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 137.600 58.330 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.870 137.600 66.150 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 137.600 73.970 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 137.600 81.330 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.870 137.600 89.150 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 137.600 96.970 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.510 137.600 104.790 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.330 137.600 112.610 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.150 137.600 120.430 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.970 137.600 128.250 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.790 137.600 136.070 140.000 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 2.400 ;
    END
  END enable
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 81.640 140.000 82.240 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 87.080 140.000 87.680 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 91.840 140.000 92.440 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 56.480 140.000 57.080 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 61.920 140.000 62.520 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 66.680 140.000 67.280 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 72.120 140.000 72.720 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 76.880 140.000 77.480 ;
    END
  END right_bottom_grid_pin_9_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 51.720 140.000 52.320 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END top_left_grid_pin_11_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 2.400 113.520 ;
    END
  END top_left_grid_pin_13_
  PIN top_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 2.400 131.200 ;
    END
  END top_left_grid_pin_15_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.400 8.800 ;
    END
  END top_left_grid_pin_1_
  PIN top_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END top_left_grid_pin_3_
  PIN top_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 2.400 43.480 ;
    END
  END top_left_grid_pin_5_
  PIN top_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 2.400 61.160 ;
    END
  END top_left_grid_pin_7_
  PIN top_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.400 78.840 ;
    END
  END top_left_grid_pin_9_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 2.080 140.000 2.680 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 3.750 0.380 138.390 128.080 ;
      LAYER met2 ;
        RECT 4.330 137.320 10.850 137.770 ;
        RECT 11.690 137.320 18.670 137.770 ;
        RECT 19.510 137.320 26.490 137.770 ;
        RECT 27.330 137.320 34.310 137.770 ;
        RECT 35.150 137.320 42.130 137.770 ;
        RECT 42.970 137.320 49.950 137.770 ;
        RECT 50.790 137.320 57.770 137.770 ;
        RECT 58.610 137.320 65.590 137.770 ;
        RECT 66.430 137.320 73.410 137.770 ;
        RECT 74.250 137.320 80.770 137.770 ;
        RECT 81.610 137.320 88.590 137.770 ;
        RECT 89.430 137.320 96.410 137.770 ;
        RECT 97.250 137.320 104.230 137.770 ;
        RECT 105.070 137.320 112.050 137.770 ;
        RECT 112.890 137.320 119.870 137.770 ;
        RECT 120.710 137.320 127.690 137.770 ;
        RECT 128.530 137.320 135.510 137.770 ;
        RECT 136.350 137.320 138.370 137.770 ;
        RECT 3.780 2.680 138.370 137.320 ;
        RECT 3.780 0.270 8.550 2.680 ;
        RECT 9.390 0.270 26.030 2.680 ;
        RECT 26.870 0.270 43.510 2.680 ;
        RECT 44.350 0.270 60.990 2.680 ;
        RECT 61.830 0.270 78.470 2.680 ;
        RECT 79.310 0.270 95.950 2.680 ;
        RECT 96.790 0.270 113.430 2.680 ;
        RECT 114.270 0.270 130.910 2.680 ;
        RECT 131.750 0.270 138.370 2.680 ;
      LAYER met3 ;
        RECT 0.310 136.320 137.200 136.720 ;
        RECT 0.310 132.960 138.650 136.320 ;
        RECT 0.310 131.600 137.200 132.960 ;
        RECT 2.800 131.560 137.200 131.600 ;
        RECT 2.800 130.200 138.650 131.560 ;
        RECT 0.310 127.520 138.650 130.200 ;
        RECT 0.310 126.120 137.200 127.520 ;
        RECT 0.310 122.760 138.650 126.120 ;
        RECT 0.310 121.360 137.200 122.760 ;
        RECT 0.310 118.000 138.650 121.360 ;
        RECT 0.310 116.600 137.200 118.000 ;
        RECT 0.310 113.920 138.650 116.600 ;
        RECT 2.800 112.560 138.650 113.920 ;
        RECT 2.800 112.520 137.200 112.560 ;
        RECT 0.310 111.160 137.200 112.520 ;
        RECT 0.310 107.800 138.650 111.160 ;
        RECT 0.310 106.400 137.200 107.800 ;
        RECT 0.310 103.040 138.650 106.400 ;
        RECT 0.310 101.640 137.200 103.040 ;
        RECT 0.310 97.600 138.650 101.640 ;
        RECT 0.310 96.240 137.200 97.600 ;
        RECT 2.800 96.200 137.200 96.240 ;
        RECT 2.800 94.840 138.650 96.200 ;
        RECT 0.310 92.840 138.650 94.840 ;
        RECT 0.310 91.440 137.200 92.840 ;
        RECT 0.310 88.080 138.650 91.440 ;
        RECT 0.310 86.680 137.200 88.080 ;
        RECT 0.310 82.640 138.650 86.680 ;
        RECT 0.310 81.240 137.200 82.640 ;
        RECT 0.310 79.240 138.650 81.240 ;
        RECT 2.800 77.880 138.650 79.240 ;
        RECT 2.800 77.840 137.200 77.880 ;
        RECT 0.310 76.480 137.200 77.840 ;
        RECT 0.310 73.120 138.650 76.480 ;
        RECT 0.310 71.720 137.200 73.120 ;
        RECT 0.310 67.680 138.650 71.720 ;
        RECT 0.310 66.280 137.200 67.680 ;
        RECT 0.310 62.920 138.650 66.280 ;
        RECT 0.310 61.560 137.200 62.920 ;
        RECT 2.800 61.520 137.200 61.560 ;
        RECT 2.800 60.160 138.650 61.520 ;
        RECT 0.310 57.480 138.650 60.160 ;
        RECT 0.310 56.080 137.200 57.480 ;
        RECT 0.310 52.720 138.650 56.080 ;
        RECT 0.310 51.320 137.200 52.720 ;
        RECT 0.310 47.960 138.650 51.320 ;
        RECT 0.310 46.560 137.200 47.960 ;
        RECT 0.310 43.880 138.650 46.560 ;
        RECT 2.800 42.520 138.650 43.880 ;
        RECT 2.800 42.480 137.200 42.520 ;
        RECT 0.310 41.120 137.200 42.480 ;
        RECT 0.310 37.760 138.650 41.120 ;
        RECT 0.310 36.360 137.200 37.760 ;
        RECT 0.310 33.000 138.650 36.360 ;
        RECT 0.310 31.600 137.200 33.000 ;
        RECT 0.310 27.560 138.650 31.600 ;
        RECT 0.310 26.200 137.200 27.560 ;
        RECT 2.800 26.160 137.200 26.200 ;
        RECT 2.800 24.800 138.650 26.160 ;
        RECT 0.310 22.800 138.650 24.800 ;
        RECT 0.310 21.400 137.200 22.800 ;
        RECT 0.310 18.040 138.650 21.400 ;
        RECT 0.310 16.640 137.200 18.040 ;
        RECT 0.310 12.600 138.650 16.640 ;
        RECT 0.310 11.200 137.200 12.600 ;
        RECT 0.310 9.200 138.650 11.200 ;
        RECT 2.800 7.840 138.650 9.200 ;
        RECT 2.800 7.800 137.200 7.840 ;
        RECT 0.310 6.440 137.200 7.800 ;
        RECT 0.310 3.080 138.650 6.440 ;
        RECT 0.310 2.680 137.200 3.080 ;
      LAYER met4 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 138.625 128.080 ;
  END
END sb_0__0_
END LIBRARY

